��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ���L����ѳJ���ף�6I	��7�"�D�}ے-��KpV��s�h�n]��[��;,��*��_�H1mTu�<'�M� ����Z�H�H�#����*ծ���p����*�R@�>���Vx�Cl/_G�b)�z)���e5��=")D9d��R�d0�� x��Ġ	\�{���> �Ueڼ{�g�_ˡ����T�x�\mB��޿8x][������v�	1)�X}� E�� �_ð[#�b�$Xt��C�
w��bGe���ʹ����UG٣�ɹ�~V��e"ѦΙo�ɱ���0�-�y�v��CPܼ�Fڀ�2@�E\1l�GN��Ϣ l�iRP'�ϙ����Y������ T�*�g���DO��� f1v�\�w������Z�2���8.�QV,���W��K��� *�,�J�6��jH�;�B�n]��CKxv���R�i-IJK�vC�?K$�Q�Ai�L�����I��L1�Cɂ��[�������x�9ئF��ty/Y��Tdto�	�^�S���/C'iy��^�,��)�:��K,϶>�e4��D��#��#�a��ÉB��� m2���pv �Ah���q�ݩ#��?-����A�1	�)W"�"Q�T�y��]�,�V��~���zZtˑE�qv��C������+	�i�����Kc����|���F���o�|B5Q�L�ν�!������q�"��?����z���AL8����B��<�x4|��<I�*��m�}��E�r{���K�B
�8� ��p�P�ĥ��X���@;;%lcKrʓE���Xȉ+A�|�7q���vI+@���dK�K���.B!xW�����4��P\�T"�8O��y��_�e�dˁ��T$)�<#[�s��6��
�|<�+F�x�� j���bw!=���jT0�����c���r_"�ÞgE$t���!\�b��$��ž��c�)�[�h�_����uK?D��Ĭ��W������B�a�PM���Z�!"c���ñi���5�Q�<�x�'�1e�Km�������F���s��&���0���X�FH-��p(���c����;�ܨjTY��G��y��?����X��&�:�z���)D:��:4-Y�1"ɓ�E�d y-����b����}���N�d���&�&�ܓ(#��k
�\��n�(�Y�Y0����y0��V�]d�\uH����6٢�98\"N�	��4S�4A�n�\TL<����������㟿�£�����8��+���Ħmo��Xm�9G��W��%�lM�<�9�}q5ɋ�)�#u����e�C͂j
n�)4;G$�,I>�
���j��S���qo��['��|
�_1J�ڛ`/|#�|LQ!��p�>s��Swq���j�����KO2-�΅ff�~S�Q$!�<�9!y]���i�AL��֨��|
�8t��1֬�8�s4�W�ǌ9��oM�L!�ǚiy�d�ꎁ�rV�$��dA%��E3�R�� �)3^_ׅXMad����wW.�1&�ªR�]ɣ��Dg �
��j*��hَᣢkW��H�՜��M�a�˯��G픗ZQ�߅��b�g5<��V$Ȭ}��sW��0M�o����H���C������z������Q�����ǭ����0�SX�kLyP�/�o�Ҿ^W�Cy"
S���2��$�Pt��y��l���Q
�k�ӟ�RR�(�J��g�G�o=�,�)nT�b������2_#�nM]�Kv����^`-������"k�᬴_�:��{�����գ�:x�{˽F���_�a>��ūLe�
��:DՇ��[a����k̵JU��9CB���o8���YՙǢ��{ �C�to%b� DHUpH�_j3�[u �*�c�NE!�LP�F&/Lc�S� y/zŪo6MxiM��Y���5�6��Wi��^Oo?����8�{����v��:�>2K�~@�*#(�'�����|E.wg�������Z��A�:��jHKG5nxE ��=�w��!��?Gҋu�x)뵍�<����f�gL d*u�b�<�iD�Ȼ����R����NĘT�8ԑ7�ߜ��
?>'����/���+��kL_�Ү�/�c�W��z���$p߼�t�5��� Ũ3�&���%�u��6E�(��ս����)��8�i�}�z�[���b�f6�c�jR���sa�V_�֣ZX��g��4��ʁ�����ӳ�EMJL�b#�˚"�������m���̱'/V��j��L���c��q`�0/�WL#�&r�2o�F	/� ky�V��,�ʈ�{�Bh����-��B�dv7�'j
">�;>�i�4沤B��_�δ���L`�ѽF�&Ts�]x�g,�q��,C�
�fZ��Ah���A�=�-k(jx����$�'����k^�ِypGv���f�>�*���㧆���t��b�*If��F ���Inq;+�'���Z�M�XeW^%^��c]��Ov�U�/��?"�a��؜��i�i���r7�UT����H��2�7�8��w ��uF�k[��I2��'�9�A#������+��Ѽ۪]꿹j���7S���=s��G�Z��nT��C 	��1	�tU�3K���X{X(=��~�RA��Ƹ����b�q���8�l���zj�}�c)3�(b>�%3��}\og ��;�W\6�,xR�w<׮��K��)�g(/�?�g�O:Z��w��?m�I�`Po��E_��Fv�=Ğ̏�
�w��x�)LS1}�=��S����1Hx�S����m_Xت	������"�uY,���x��9�׋cE���v.�Pk�F�>J��T�-�H���Y�um�_�'�tI8bp.;�	Je���r�p�iؿ��O �zD|�*�H��A�*�撅�L]�?���YX��5򓡹� �afp &w9������+VŰ]WML��A���7�.��@D�ꍈ�/Ҍ2穢�ez�=�P�g�*3[��|�S؆����HɝѦ'�^���K>�7P,z1
"R��S[�P�ZC��8���	��q:��hH��^?��}��M����,"�R%iӚb��z�d	��.s2Kx'� )�ֆ����j��#��"7	\\X��m�t*�n���W���ٷ��D��]�]P�R��d� �K^Pߑ�~�Y��z�G6F��J\�w���t��o��3�t�?Pl�־��*>l["���u�Z}����d=�߻Cr6�p�����g� �h��E������d��T W�A`�������;مȉ+�?�˖v� Jk�f��t�y	���Qz��������A/'���`E [���,���]���P��c��Pn���&�9�(�K�9�����Q|:}��~�LSK�r��^}e
��~$/�i.M�x[���#.�U�g���F���ֺ��9�59��>�mOy�Y�U����S�Q�i��B�L�/����R��QjU��Bj��_���
�X�]%˥^�Xu��{L�|��R�UqJ/�G�l�j7����4V8����QͿkzxͦ�N������KMB5�X)y�"'���˕�{K�S�j*�|WH�H 
����?�K��?�3��N��\q�o�8f%Q���9���n�z�Ѕ�r1�6ނ{�Z\��;�5��}��y�ۜ�C[�L&��ۆ�՞�E��7�!����\w��(�oC�	���[�X�* ��"O��(�*����tw=DE�h�/,��
I�MPm� ����+����,�'�$ ���tⅆ��\b�q'[ݛⲔ?@��'�詨1�?�����Y�O@�9�A9���f|��9���F7k���V��9c�E����a�|�_"��瓋q����������CH�
���"o/�6���v�~9��(|�,���;&���'���A:��X�&���G��r�|J�UL�O>���x�@|����No�>�� �C	�B�����"��BF��z#_$��_?�U���`=�k�d�]��h�����ZM7;��ֺ!�'!k�%N��.b�Hzl�����rc'�Y��¥�H	��A���&�e���Ӂl�"�D�a#'���q=j��V�XW��b�:K41�}�����l|�8c��Z��]�*�$i�(��voE��"(���O��l�=�<�;P�|<�U�&H�ۻ�>seU������t�����Z5i�w���N�łXl�����2߂V�%�JB\��F��1W})'Q=�uxJ$.���@�{�!�Kɤڱ�j��ڡ��۲N&�����y9�YXy��bpʶ�,u�x��+��z�cX ���Cժ�gA��u�f�=��J����f?nFf.ĭ׻$�j�DcJo���a&L�����	]�K��0��ry������l}�A�GEM�2�8�#~�6��ը:}������~=`�a���q����X��Z b ��v��Õ���\�j�MEQ4��5n��~Ίt�Z*��/&�n��ɡ�>���4k ��%����}g�	^놥d�/�ض��՞��h�Ť#7�z���&�(=������h�����k౱(�����ܴdX�/s2#�� Х
g�w5Ǥ�L�o	>߇�����@�-�*��6|� {��J5p��+ҟV4��9K�5	��
�*0���t#=�������S�FcJ�e�(�^�'z﬍η;"�?y�W(�K��a�<&駶t�6������C)=��Za,������A���86��Ay���J�s�ϓ �g;�����#��{��Ĭ���0�y�͇��9��:�)tfH+��J�n�$M����CW���6<h$�Np#����f�ќy��P�E7���)īYЬ�{����c8ƻ�4���.��_:Wќl��p�����c����6B�Y<=NQ�v-�+-�?p���|n	�J��T�PF�_F�M���T�,p0��� �Eo�M���R���~�������m��Q�h6$��	'2Ƨ����z�$F�m��GccTԘe���S�͜7���圎��o�l�
��\���l���.&�|\�A�L�� ��U�\�B�*��O�NE�I�L�X"��/ˠ��T~����}��lg  �L�3?{}N������⢋�L؞P �����]�0�����3�n�v�`b"1�ŭQpQ�F[���,x��T��-�׻�t>:SprǦ`E�x�E�r�%�~C�[�1�nc��u�Șt@L�R�%� �l��;b q?n1��T��8�,��1|�����KjJ��LLZ���\�o(*lc𻇑����ك���aO�G!#�����!��l�D�3�%�u
�64��s�S0e�7<??����+��7)�Y����u��n|/u�N�K�8V���޳���N���9,} H��v��b�{�@���|�4	��\�5Xͷ���y�22�)�T��v��+lX�p�G�͝?_��j�e�s��{{@�N�e��Y�>�z	`G��V���Э�����d�g�,E����9uJN�ѝ��&I�Ϻ@@Qa<�پ:ω#���lll�4`To��ň1��𮡠��2�J 7&�f�yb\�"�k������r��%C�J�֐�塆w�ALPt ݧث6:��ԟ_E���>�W�Z<�ԑA��M����y�p��� ����w��� �Gr���(y=�6l�`W��>��R*x� ��?�%�=[�6���&bI��C���/s�O÷�f�P�Q�οGX�&O��_A��_�tf#�������\<d��At3>�.-?�|Pۀ/���M�cW�������	�>'ɂ�� =��?��G�)k嫬Vl�gp�c��j�B�zND4���d���vI�6�HMV�h��
�==�[�'3�T�xs��M��5���1(ᖪ��w"�m(���B�/�(����=Ģ->P��+���E�&�A8���J�J�sq�ZK�D(4�lhԺ��^��: �Ҍ����N��d�G���B��E�P@�]bh�.)��YՊ��^�2���.���SDS��1}�:x����a��%�7/y�*R7�<:���t�N�Ê���X\d1����M @���8��[��)�ϧ�W�R菏v�HC#�]8�Td�gJ��a�����y;Ǭ�����
ME+׹�1n����Vǻ� ���c&N?�sH��-4��̅F�E'��tZZ:U��X��x	;���'���1�!�	e�.2tt��m�[XުZ[q��N���P����24#٧Y�)r-��\�^� >3�6 k<���۸7�� B��d6���#s�_���
X�Fm�T��
X	��n1��u���IH���>E�iO�2�����C�.W(����ZO��֘���3��:!-%�W�4�H���	�e/V�V��C�$�]�����y^���RBFhR���$eU���7̈́�T�E�Rk_��"'���y �U�VNul�%4.偍�g�����=)�v6�3��l�4���m��B{b������;8�*��S��
t5\�B��zce����k�|[)���{�� ��x�s�i���=>� K��^�^�C%�pu��U�6/G�a�陒���u�O�8�wWb��ʽdc���a���F0�<ptt5�=��j������ڍ�%Y˙:.��{w�!J�&d���F��4_ٳø6t��Ӿ7�v��h��J>��A(<�(��V�&r$劥s�NPe���a�h�A!���@{�!"H�c7���Ğ�)<4'����J��@��[�&-a�V��|�,kp��b�18�T��W
F!�Vڸ����8eMܶ��Ъ��囉�d��9�^*���:�+Fx��/��c��j�;2��~x6��֫��BE���~'*@낝!��
�K�l#�:���uBI�D`�o%}�e��̾5��qZ=�|��P���I��7.�b��"k?�ˎ_b�� A[�k.�@�-��AJ�3��JĜ\�ϯ�@�\�ͩyV���A�cZ� ��'��h/F�����S'���?�������@7��һ(O�H]�}���f�%��?ܹ*M��H �H=9�4��jn8��cd�0׆k�keRoI��-��bJ^��]��X�p��ce5�+�jww�yB�O�!:��n�i�_1f�9�[�
k�?�
�zA�19��5*u��a��$�B��\� aQ���<k�g��`/���TGUS���"Y��.5�df/��L��_�}������i��ч�bRa�o[��r�$��;a��#'����c�� �:�gzOA�k����Of�&H���z$�p�_� [U�8ٹ��9 S��/��-2v�vY���2�\�(k��7hғZ������rK���~-��1^�r$a~6}�)E�^Y�1V���3*����Px����9C�K��YiT��9��g�9|6�J+���M_A��;Tt9f��2��/��g��+�������dB��h��ˬ���	�B��=�J$�z�b >N�!���>��R�'m�w�Q�![�A�j�n?ů�FqIuY+׺&�Vܰ���*G\�M�v������{�@��G��$z�k�+�,+�C���W��u#yFH�� ('��A�xd'�T�2����Q�+�S�ߓ��t���]H����^�pR|�A�&���GM��y:��0 
��v�w��~�/)�7����f�������um
YA��o�]���?ҚQ����T
!���j���QıwE:����*��+�n]2�/;�s�7wsM~
LgZ	]���o�i9Ə��PȳZ��L^ Gpe�j�7�hm���x���+(��=���7u4�'��&��LI~|�L8?/Ŕ�p��0��ϖ|�t��T�n��d�:�az��;PКb�c�� �{Nخd��)b��c�~j�\��o]O&i�[������EJg~�w���w�X�J�6�4��*z��>�݇�i�=_6n9��gi�.�>�g�*�{�6�����@�c����Η9p��No�{C��d�]��ߢ7kh:w7u�-E�QN��Ri3����,�ΡŎ��Ǡ�)�Y]m ��5�@��Ҝ�� Μ�����t�8Q�����dY���T�[�k�`�l������ܡ�b?^-���s�'���_+�����{
r
j��(�E��-����O�?f����NV�TVX����fr��+����-ٛ���)�\&H	)ɰ6���M\�,��՝H�!��Oe���}�٢���S��G�����5��K�룎%g
Z�s�T�|����=bo����/�$h���РH����t���6���Y�L�X)_��T]#�Ǐ�1���0y��@������̩H�	�g+իH���@Δ�����<Cu��֓�-K���Uu�N8,̺��%S厇'�Pv���;~H��A��y�6��.��0�h)O�e>R�<H)���8=��@�����S��*�|�J�H0j��.b�zTyV��K����횧��h�OP2>D����N�l�j0����n��^�A.0�j�X*B��o���cS&�B��p��+)"g���S�)�Mz��	;J	xPX�8�<x�h����X����@����w�9
dF�,��t���Y��鋕څ[� �`���&�����:�j	�^܇f`%�pſ9�箝��|b�%,�Yy�P�=ɼ�}U�pB0�[�3�J+h��r�e\����8�-x�!^�ie5�.�-VQ�H����g��9�O�c�Y��h}{/ݷ���>�$=N��u�qg��������yk�l�������1��m]�dx�Da���c:��'Z}Y�����b��K�e���\�0�0$=���g���B�p�^!�V3+}�����~2c@�wM&������4�r�i^+y����m��F|���T@Ǎ>�Qz�V��,jo&�j�zW"O�v�������#3NO]'k )}��r����`��yY��"o0[�F��}o�#iӮM-s}Tj��p���ЏB]��"�+� ������ds���K[T�i��,��H�.Έ�X#�˿��Oasթ���^Y�}��(}��ߢ�J[�a�+g����}IYQ��T�n�|5�r�a����^���Z�G$c�"����Z�����À����"$���!�� U.ʻ.�~Z��-7�gr�
d�t����]���	.�(�\�Wd�b�ԆNÉ�|�C���[z$!�#����׊���?8���m���[��*��ɛaxLGg��6��+"l�.h���Ƽm�YT�V��u`/�_z��|�O���p���(Di���6�g�����k+�� )e���yy��|�[�6��.��S�V���l��9�=J^w��hp3(�C#j���Ix�PJ<� �xm�0g e�,q�2�����t�O��0����.�Ez�F�nE�'Bڱ�Fj<�@�e�3�u:�a/!�����
�`�H��P�wY��.q��X9�}/��v�� ��?����(�
��]|��t��e"���-�/��ڪ��"�y�{�,�V��$�9��x+C���v������@Q��~;Ck�����$ᙪ����.`� ��`4�EK�7ή���C͂<K�}b���X�)p�Y7�X"�?�S��b$tp�Ʋ:�;�g|�HF�lz�)�C�:Oy�G���-�kx�.h�7K�|��$!�.�ґ�}8�<�:H�^���r��lx��ȃ�톤$[�A��()��d�&k�γ�)*m�Ĺ:Z<��](��~?�F�+5sGNG��8��|�j��F>0fA=��H�w]0��$ԉ��$����'�JO��4��j���̥?�>�~��0U;�_�v�QǢ?��r&�
B>Z �����0�)$�t ��������{���Q���M�Bb6��K3��h���1�v:	��Ȅ���wj�ʰ�7�c�fׄ��<����P�z5�V�PZa5��x3zD>Z�f��O��+�mW���2����n[Q����nj�չ��D��h�̇	hrz�QA�����y���� �Dv�`��8�.�a%�S�A�����4��E��+P�}q�C���o��w�J���x1�A�f�z&���uɀ!�Wy�4�(gj�§P��160�5����m\ecg���`ľ��J7b��Qd=d���^z�۟�Y�Ѽf�`��RLS4�Ɂ��

PM�홪��>�S��Y͹�pШEChs��2�+'/�rLF ,qK�'��C�u�o�R�ǖ�+A&sÚ��r$L����Z�R��<A��+P���/����\�b=6������ҺT6��Ղ�����=�W$o;��P���!2^G�T�ֶ��7�~8��e���~�lQ�<HO��3�-7�g��)0�Za�������fn#��C��T��S�V��q��d��k�J�
J���z�U�S�7!���N5:���16�"��q �K�kE��A|^�����D)�
u�'�PD��4�:�������F��oՒ��p�ː�`~ɭڬBV~��KZ`D����\��^	�����r���v��Qr���:�9�{M>������[�*�� #�r�ɶ�-���ؑ;�ͷ����?'[s�	�|���N6�*��޺<|����U'ׂQIA�J,�!"����q
��U<�n�5�eU���������+�B�P-�)�ݣvR��;�fh���[�2�;#�-$C���ۼtx�A��=��\n�'�K{T��Ir��w���9��-�N]�Q�Z�'�����G�,7������5�&D=V��'��o���i�X�F+
ǚH[¸<{KJ �H�zbݾ�sE�h�m��y��#>2s<�,�����i�6��=��z��f�%t��e�U9B)N�3��\omR���j����Du�d<٥#uZ��fm���Z�5Ҁl��@[���ڥ����>��Y)���~���/���h��^���k��$��@���:�����,pR������6���I�L�-�h�"bS���08����vKU���_ħ��aq�����G��v�MLv��}�|��}ϔ����M���ۚ3̴11�g=��hq��j\��I�9'��@x.���gS�/��i'�J��D�}}Ի`��O,t_�S2N~��&lla�}��q�j�6���
i`ධ�Z怣��%�[4�ފ��h��u���y�\��b��SD�-%a֜X�$�m��D�R�v0]�
|M�-����	��j��צU�Y��aR�� ��@a r�f���Ͱ���-����2��<��l�B��bt�*G>��G<�|��~����ܫt{k�,�N�V9��v0+<v��aC�LR Y�B] +B���O���]���TD�K�t���m!~/���Q7Nn�we�<�#^`bEZ�T�5�]�Ef
�m�~�N����0ҲJ��a6�9KZˌ{"QtP�#�k�j ��FH�Y�FD>�B��6�q٘�V�Y�_�Ɋ�3sG�'|�3ݬ���t,"q�����ZN��yF� ���I�IVWwf�1�UyJ��9��5��A,��K�ft(9�h�;��-���V�x��>,nܞ9*���r�� ǆ+�'�^nka
m{:�m��EŖ޻v�e�ʓPum��/�͈S%ғZr��reĄ
��C[; J��u�¬С��mg�~a�wM���N�``��N�:J2��*�.r�@�=Z�K(�K�)� �P���QX7�����!�9`r��k���>t�GR�[���'�_�($�O����ǔ��L�PE�Z�D�\���u��.�\����
,���#�S²�Ъ�TlC�G��O+�+H]*4����jT{�皇}�D#���x�7�м��?-��.L �v�0ZS����?���[ao��g�"CW�y3�Z�������z&��{�,���V�\O6I��m:�b����s�UZ��C�����Cj�.�jC���_q��0١C"'�Dj�a2��#��lP�֎È�A6��_K}��QÇ�Γ��ޠ�q��v�}P�nʥ��X�qǠ{!�YȢ�k�_��/ %?+%�;�}e#���/���5C>��Q7Z��6	�'Kt�_g��a ��ꊗ�Z�����8�L���QD�����e��UT�V(^ ]�����uP����j��D�5O��p�No&�	�q��G��ĸ�0�ۈH�o�n�]l�y?� ���ـ�Bdz�A9���q��c\eT����	�fn�)L4�˰�?'�f�k�_Q�F �@S}���%[��ֲ���3�[��u�>�B�ʞH|�����mJC��ڕ�o!u���W��4�n�����T���9��AS8l\6-�k���}A�Ϣa�T��}[���;i�Ɂq��<��hfE}6��yLend5�2���`��NaL�%������@m��\��{q�G�`���e\U�Z��J9���p"0���Y�jf�E�|&5[;� '��;ep*��o��J�L4�F��>?�`�����<��� �)3M�0qXQ�� w~�і�ݭ���H
ۦ"
y����>ߏ6y�a���醐pľӘ��䌼C̸U�;�s`fOmj*�2e?�eoD��B���_=�{?�Ȍ)XS�%���UC�m�,�x�}�_Z� �ZA���c��PZ�Qn��	:ZrոT��q�J�(?�־ŧȁ0K���J���dj����h��k�yw�����9Kk���|�)a�Ygv�?
$�����jꐢ�H7#L�?7 �թ��
!�ڪ�'�7��a��������0LS6�H����H�H�������bfG=�E�CT���$c ��;���ǰ� qv�S�`���Wm����L�9����?D.[��D�G�Ӟ��Մm�bQ�N��[j�t^+�E��D�eCAvV8�u�|�x�y(V�GL��`~�1�Oq:�Ðo���D�.:4qG�!c�5F�t�nô���bv/yIO���W��V��`�MQ�<��1l�u��sa�"�\Pj��#�2{A������i�X'n���Ɣ�Y��>�+>�W��}��B�w�T b�ă*A�e�b�Q�j�&?�RE�}��
�t�#�L�w�H�耓aS�'�=~������$��q>^9�`�����mR�����ɟ�f�(T�,�K$�  �!�d�i�#����۠�L�Y�49*�"��7� 8؝���X�������Sj�|�F�B�.�����U"w�$Չ��7k�1|��%V+$�M���*�Q+&�e����+!~iT@?�ʮ��KOv�٫Kq���F%��2�ƹ"o{Z���"��0���iP͓��_S%\�g��E@������m�n��J;2P�1�����	YA���Yf^����"U�;��7���`�n�E&tR~�Bd��+e��d\)|�sf��k���b�C�,C-�������4c=�1SŤ{D 	m�3P�b1|�P浯�����"� 7�71�a�;Y0��L
�+��}w�R7�����%����>&&6��s�ί�T����8e!d���D=3g��j��`��(ɪ]�	�^Bt����rG�f>�ğk���#mARD{C���B���sR�Pp�љ\@�u��+���.�3MT��i�[K�pu�jgG���#��l�3zªZ�N��'t*��Q�.H��Z}2�k�� ��Gr�`�)����8B����쥅^
�h8�F*fT�+i�j���9��1&D� ��0ÑX�h����ӖO�P��2
�7�4˘n�8��o�4c/��h�4��mM6 ��\�ω��ǫ��4����^K/��n�9�5��ž4�Dű��I���dTf�D~-Rb�2��N��K&RӱNǾ�J;{S駭�[&���ˆ���R��c�ζ.��t�K=3�o
�Y��Z�z`/K��
����OD�n�H������S�4���Mu��[[�ƪ/���q���
Ҩ���I��7
����_��@Z5ӹ��㣑�9�yʄ_h������?X��dq����qF��]:u�̹MY�� �cq��-�R�i��qW�Y��#��_�*�s�M�	T�yu�s�hf}'�|�߻��}56��`9�T��x�x��W
V�ܤ�cbudkjF�bUܻK�>e��D�����
�u�T�-�<��SB1��k���r�?u#���.!ы(uų�6�V1�FGJ�� �ua�{
n$[�g�J�Q�';�2|��	4��!*;�_yV���D�S
�v"�}�����k_������G���L�_��$BA��|����=��]y�Ӻ�U$�CX BT��k���gY[��=�w��ǆC�ӴO�k�Ə�|���)#��]�o����͞ф����ʉ��QnZ�M�Y��z�	��FJ�J�D�[	���Z=�D�rx3fFT��4�Tt19�i�)�����ŐX-I��YYʂ��{�q��2熁��+�BE%��lu���'S0$c=�� l��b	��]X;$�لк�]��4��b )E��2�_Ѭ�Ew��,p�K�`��<QF8��޸�_����@\� �h�����E�_*\����#���0-c��b�>D��O-ysa�-ef/x��l��) �����r�p�g>Ӹ��/$��*LVl�iR;\���b��i��=uF��ZF+G�����'	���Gi�jo��xXݲ?��v��";ٝ�\[&���N�B���'FZpu����2�ԥ��]��)f�r'�)<�	�b��
'�!�opw����$f�],�bhB;��Ч�i��4���۰_��^i`)�CxأWf�J��R&:N2���dOg�f�F�[� �x���>|��M����z�]�4l��;�*�<�i?4�ֲ����#Ƕ���Sv�����B1���fV(�cK��_���4A�~.U��cQ��<���F���抦B{��Žuͼ�[°���,�i@x"K=��m.����f��[=|�:�9��	g��5e��$�'��>�f*�ѝ����'3j?�"g<���)������Fx��S����[U��p���*wFkgX�YZ��uk�:�5a%z(%��4�������+���nE�����_(7��tM,�%�FV����� �������Q~I�գg�ԈY�+�6Ƶ����S�-���osL�k��jq���Ѷ$4�]��B��חSN��f��з3(�~%%�ZT��
4a�.�K\+�4�ׅ�?�h��� �hU*�$]~�U� }�� �!�Zi�@�O/(9'��Gt���	����}�ƞ�̌h�I��H�mU��K���<�M/�ޣ6�B�~3s��$״����ƍ�C^
�N�ǟT�&�B?�ю�dC0ʃFi���U��H�c�FyX�r8��\�����G���Sq��#7�-�'q#Q�5h��cv�B�4�z&ˮX&�����=�j�|i%�0�Yf�k��S��$DK�j��*-;����" {���aF�ST�Y?rkm1���lP�U�@�lV�-9S?Y��g̋Zo���Bj�����d��i����6v�
.�DZ,w�خ���ٸʕ�`�[y��1*Ou}���Q������]t�����V�]0랡��u*�FQA&���y�y��+ͭ}{��.�r��Ny�o#�]$er�#�!�5�������	rg�Rz)T�h� �9��p;����n��[�?2��#��HqF/ګ,�����.�ZՆ? �ew���2�(�z�L��qlx�J���K7u�i� ޹�y��V�����E�!m �|w�iq�_�W�� ���~���=�hڪE�]�(=wD�b��x�G�Ա�Iibӹ��
���UW��i�/5����f8 )�>W;Dȯ[Ձ��|l��@e�Mh���k��m|�!7�QXːQ���dX�5Q0�l@2�1�� C�SH���:n/z�y�|���@5{ �Bcr�#Y��Γ�_��=�O�����@ ����=Q �t�-|�͆!�e���;H`ܲ�=E�<YI��uI`�9���8��ހ���(�ad���y�	�р��{�M���(�A�Pf�OB�ڑ���\ȿ������ ײ�Y8 ��m�p�yR7����}�G�W����~1ɒ���1�d���[�T*ƫ(zrh�2䭣~��MkMC݅~���(=;%t��)�qg�MpȆjQ� ����6#����V��hy5�@7�O/%� s0]XE=^;zӬ�Д���ͦ�w�;d�vt��\�o�<�|���^j�Y��R��xd;���GBt����ٓ�4����T7����'��G�~z��>�2lR ��$���V�mGߙ"N5����L��(9D�1f_�ؑ�%�<Kv>o�v���v�P�_�F��7����N�JFPa�v;6$��d��|�N[���*�
>�����,�ނg�8��/ܷ8ó(��vR|�.u�lh Q+�u �q��eP#�<0z8�ꟶ��:B4�b�\m�^v���TM~�ik�����=�ge���ڭ�U��l��R�T�s�bu gE��4��=�E,��ԏ�p��XN��G���x�h��,��ض
{6zm�����X;:$��|����Pv+l�X�d��=D���k�C��HS�,&���R�8:�/N��:���$�Gr��g��#�c�O�Q�=�a�r�6�i-_v:t�wB��-�v���$�-ݭ?��,�/��P��m�OO��Q�7�
���,��A��Q�@/��?�-Xu)�܂iѢΦo�;y�H=�B���j�������LՎ��R;�2�!iS�*�T������'���e��U���n�jI>���E�lL�L8w��Wf��	}�\������i,	�r&})$�k^��:.�5�P|&_7;����Ӗ�����JX)Q���Qm��d*���D��}?�Y�zs���_ZcB��"�z�XO��5���<$Q�뗍ek!��p{�o�m�S��Z��j'�����:�H�)��s7�d�H7#Ҧ�f�����k�� �&����RJA	~_��S5E�[�z�n�K�#�J� /�B�s��(��Y�+=�o�f�-7����5�(N�mGd'�̞��ea~R�+:���QCR:�gp5�M���!�C�Gc���kFBI[�e�a�{E�� �	�9vŘ,'�,�*l捝�DJ�]T�T<���i�8�ʋUܘ����Lg��8�c�Z��
��+F�_N&�X�����?�x!]�
��O�6�`�7p��A�m~���U�[��r�_�=��]���H��Ʉ�"�+�_�z/%���ˀ��l���_�A}]��!�*
ժf��X�F�Wx���R��K(��΍x�'=K��A���w:�BAvNZ��>�1�o�r������I�����Fa�����[��%�U�N���xJZ8Rdn�GOn�.�f�ε¨�L�r8}�ŵ��-��(2������]��B�-j����T{1�,����
Zk�Goz����!�ɤT~��7M64�;M��y�n��O8��(�\L`�8(�Uɸ0�3賊7cA�>�1���Ş�n��ީ��Ԥ�̽8���'�U����;qs�}c�������M_�E�9o֪2%X�A�a��_4X{!�$T��H�P��	|�К���'y�a�X��Ŝ��x�):��R���r�#�j!�6���qv3�v�Z�5�\�
�
J�>B�Z���ָ"�!�cV��u�a蓫~��RM��
_G����-(��H\�@����Y0�F.a\?MJ٣�s���R�K �3Ȗe�dg�n��dPD�.�DB�-hN�����#�ȟjh2��IM����I%�˹�U4ۚ�(��)����qH�0���R�I�)�'Z*�c�(����Q��c��A���7��qQ04���d��$��ca�K�m*Q�Y�����Σ��qr�E��Z�~a����A�I�OiW:]��Ce�|�M6��v����!�^�]��@W
ț�0�K��N{|g�t"�Y�����8훾���b'��E�'Q,�_#��lT¥c��F�^�dm��d8��㽎j�R����YBۑ����Nu��=y��ɢP��eyB@z(>|P����q?�=�qE�Ggl����4`�Ƿ`Pf(�Q��H�'��?TF�98��/_�9χ�p-i������у��tX���M �<53������O@m"oZ����J�x�i�=�յK�*��7U	��}\r�q��M}�B���S��9T��;eh4u�7ڦ �Ǟ���qʓ�N��i��@C@�N�Ɩ�+v�G�^��ʵ����W� 	'k�j���D�Yy`'�b��L��/�
����ڗ���*���2���%%�7�u��d�zv�����֬#��ࢅ��e��O;�L��ѓ�z�[()��+���1^��ĺGY+�k*���Ѕ�n�&)�b����>Z2T��=2�۞6������Z��b�Ͽ�d4OE	tlg��*���N�m�4⏽�O�L�ՙ��ԫ.Z�n�c<�v��VNE�娛Dݏ;&��@�ad�(n@R��NI"���bH�K8��*��2Y�f�s�c<���U��g{%�8�H���Ȋg���è����@���/��.���iF[p�|��~DRڷg�c���ߔ���8M�UjA6|���N��ǮZ������� ���0Fn���Sn:�W�r��o9��-���i�[��V����<wz_�1���������>+\��ְA����Cˉ�Ni��bR�Ǿ!5�����1}VMٲ�9�E��̠d��Xv�J��4o�z6������80*���&oS�Aa���%�DX�b�5������m��
,� ��|l����,�/���k�S�$�K�0�F��}���Y���<��4W��{���u�p�������IT�+�k��/��./Eҧ�=*2Q[����h9;��ԝ��|њdQ|��;�!JJW s7�I'���c�y���DF{�02����9]@����G���o<쟳�y�.oh뾞� ���l�V*�t��m�dd�?M
�F)Mf!�l�o�V�&�����fo+%��߶%y����]־ �k�� FP���~a}R�L��ST��_��.��M�&�Ͼ�Tk`h{q�� ����ס6N��?�u�
H�������X�(ϋ=O2�=Xl��",hz��҆�d'�r.JR��)!ND_
y2.�z�Р	FëOH���C��JR����84�)<`�; �U��	x��3n�i�Q���=,o:;%KV����fm�^��X��(�sgU���W
�б3)���:�|�N:3�^���6H[g�<}��������F��$|lD��
���bTu�c���<��"�p��d�{alu�����H'�Ml���!�����Ur޹[F���u�wy_f��B�*�x�l2��lV䄆"3l�'�H��R�wc7ɧ56��;c���
�
��,�v�q�JK�PM����.�>��P���[:+��m��DZap����a�Y��|�h�����,4|�r�r��&���^�鍪�:�t��q5��&j)��-��R�$�94�A�Dt��r��0�}`��W���fޙ`��>�r��v��o�szݗ��ksE��_K���𻆘�W��S��_�6zm�s���u#֎�2����?���H�s����Y1���<j�!�ID��\i3N�P���>�w�d�`���<��iSiخZ+���>�fap�>�o�yr�؅c��c3Y�ţqG�6��2�;�r��l�2H~8���1%�5�c׽����kW%�zv2��1�o�g`�I�������>�]#r�:��i���(⢴=t	>d��&�%��o�iFQ	b�Y1d@�x�ƵH��A�Є��Y�*E)�8rh`Y}Qb*��t�
p)=�NZ�@�ob�s�YE�@�yR�3*�=9ð߫�L�K*�mnn�رu[W���IJ��X6�wTh�Y�^���Ŕ���&fM�0�}ρU�9�[0Das��`�(�67R������ߥ���:��j9��D�:�L�2��Vw��}��@�n]F�6��}D6�������{���v���2�>��W�g���v�r3�H�}�HN]�1Q�m�-�^Ji��_���=
�#7�r��=��D�3r1ǆ�������,�[/�;��q	�|�|Y�*�.5�p= �[�3Z��Z$��u�(,^a�d��e!+� �28%������#�n�tk%h��;2r��q
�1����-�]�(MirWzB|)��ci.4�xm�"7F��~��[܇Ll�en���F�U�#~^aQ޶��B�B�Ĉ�_ڧkQ�\
/��&s}�w8m�đEZ�Y�X<w�3�i���H{���U��$���0���tH�b:���)"��Ոj9��U\�Xb���1V ǽXd$ ��nd�[�F8�߈7\h���o�kȘac��u�Ŗ?:_i��>[�����6��TMI�@�0
��o��0��$�2�������b����4P�m.�v�:����2��)�k�ct�z�cZ��l�6�*?<�p���3���E?��2�.[rn;?���f��4vJp�2So���s��B;8����1�3�_mh 9<Hit1o��!t���3Y�o��(��Oi����s�o�X"*ׄk�7(7�������U�b~�zg���R�=P��}��C�4�:���S*�g;�:��2m���J����^�f(9Y�weelub/5���M��3�,G��h�V&�KB\�J�)Qqt�#� �@ٽ��9�-��j���d�O�����Y)B�~̗��{F+x�I*�����P��������K}���R�RX��ٌ2�'�	��j��Gv�NB�&�H��l)��*��~"�\���_��t���qC��سٮ݃KBv�2���<c�J����L1��g��_�-U"(��qok��2"��5{���W�Fu�M�8{
�O+3uW���й4���x���H1 ��Ӭ'�������.h�ԭ1M��
�	u�8N�]����f]��E{Ǩ���'(`,�f�P@M���@��"7�Z.ѕ+�B?԰wU2�q�9Z�ޤ{�8�w�]�����S�@.Z_�b!��YU?�Уƈ�%x��F
6p싒^�(|̠^$��`��]��+ރ��kN��\͆fێR3�3t���9��ϝv ��l! R��x�:L��њ�6���'i��Ar-����Hn��Y���b��F)[�ߠX�����$��.��N�fdŹ{�#�쐮���+�a�j�c�������V�y����L+�D�;������ps�C����o�8s�����m��=�������-���{�6^iʦиT9���{�'��ؐ��N�����͒�-4��2l�z��I����Q�J��I���M�h(�q�i��l�R�b^t^:��FH̡��m��	+d�A��Y�e���iL>-����l�!P�4н,�\nF���=&��N��j�<�k�rQ~��	03l�iPS���&�Ů6,��d��w��U}�1��f�	�%Us'�2�x���,�����yj����`Q�0ρ���[����(�'�ݹ�ü)���=-�Hc����Aj��X1���՝�HC޷kZ�͡�(�Y�02s+Y�9��ɩY���[���6y��Ѯ=�殡~��N_��\�0B��*z�K���T!c���#5�td��S�:*I�=�+YAW'�!��>�g�A*�T����~}��ф+�~6���=�&�P3�%��9&*�Y��}I�E�@�ꗩ�dQLǪ����ŎI�o��xڢ%W `VY������o�(,d�����칳�1�R�IfW}izA��b���̟ɉ���_��W*��;�����y��g�^� ���d�y�wHM�-P�������V�����4����Ns��\���t��,(���6�<>�k�R���}Y��M��ĕ�Q�{����|u�:do�X��w���~Gb��z�rn�:J��`z²�R��aNj� �I��˄$g��σsCm���b<"'�B�j��L�R<-�	)�H��w�5Q��0���?�Xk�#�]gҺ�W���i��oT-�pנ�RQ�7EZ�I�u0L:�6�{%Wz/�: �q�b�of%���R�~k'�h�H�Xo!�J�Z!�%�xw9�J$;|�cùl)g�ªi�q7K6i�rOȍ��?	t�����c(eӋ��`��>�.�(̪f`�����4R�����ǋ�T�j�~�ܕ�OF^$`��gOd\~�S�P���"�A(�?u#˽�#��ˮ�M#�]<���� ���F?Z��!�T�Z(�Hu�?ӈ�1�n�!�q�ٲ<$P�4(%��������s"	X!����7n�[2���1C�?O���۔�̘�O�aQ8m�wh�u�� �y9�"c�VV����<�A�_5��JJ��Bv1��K�#�5a<�&���r1�Y(ДI?vmRDO�ַF��^?�P�4���4����%�w��)�{��u��WR����h�5x�D�͢��:K	QT�*]+�����HC6%b��e�C�B#�&8�W����_%���!���b^��AC���e&�	kH���>�f���7�2��oO�.t��^V�����G���k ^ag,���Z�+�K���]xO��(S$tէU(��m�]uv�2�\4�2��x�p7Zxi,E�U�O7��x���0H���v����S���a�ږ��シBH��n��s��[G=��2x,G��ά�����%��z�|�	��#����`xlSHX���O.1��P��5ۧn�{ԨQ�u�s��v l˶���|���n :�|]��蹴�0Nm��*h��h��(o&������� �\z��i|�ǈh�b��ab�P`���_N��y�v	 hT�㲛�l�;���� :��,��T��-�=���h��_���(����*j,|�HK*s�s�C�j��D$�5����0��Zp?S�W6��d�%U� �ѡ�)����U��EA���FGy�3ɵF��^�D�*�t�A��ʜ9��D���
w����ш�U,��T�JIF��8ɍ��rt|
y�ʵ�b::���{�݈��^n`�"2�hA�@/E�0�!����띩^��IRC�篴�&� P��K<]ѮLл����*��Bn�s�}��!U�_W�`5 �p=v�5I�R8#��G�`�-?�ȼ�h�K�!>?�|;&�`JО�]t��V>\�8ᯱǤ!���ame�X*���+�H�6�%qɛ�E]<���c��c�I��h�ns�*	V3ｔrڳ�]?r"^gg�T���e��Vg��^����W�$�����������%&�޲I*��>��U	
��ߛ�ZI�(�F9�H+Ćc�P� �JR�dEg�*���;nYǝ*>��kGT X(D�Iv\q��T����b��v��l�Oՠ�`
�rB�4׫x���_`U���A
I���\,y����K��s(`��K�{v�71E�s�w��������閄�P�� �6g ���^��xX��7!�J���CT�-h!Uk�O��cx��F9�)%���=�$�L}ۋ�-xm�=�>��9� ��w�Xζ5����Xe<�b��v�ZBH�<?��Xll!���}炆:W����������~�iD��%P���d�_�pM����أ6��A�ځ���bUR��76#}>N���Jn+-^�hI�N�C���;P�$^����C ٮH��8c�3y����K�N��r��*�~U�Ѵ�	�����	���oTgM��m��!܅��O�)�R:W���-����J��怆}q.*}�������m��Qβ�p?>Y�8���v�p���6����Jbo6�R�����H�� ��Bf�G���^���Z#���~ҽ�N~�@ٜJ�O~����1�m�"�q����<� 葄Ȍ��X��,�Q�?���a�к�r][�R��Kҟ���������3f67��嵲yf�f)��'�� ���0w��uG�ؼ�hW��W"wg8ءQ�aV�(����zI�U|�K>�˵��(l���?oś?E��<�]�`B�_z�t���?^��P2ow`RV�4̥D�m*V$�i6���TJ&�e�p�	�
H��ׁۭl)=!A��X�8\��Bl���ٵ	���#U�P&�ŕ�����k��0�e�S!Ǚx�/�h�!%��TĲ��a�.(pM3��˓�T{q�"xH�ҙ� ?�/ǲ�匓J�[h�l���-�hx/*]�K��%�rc�{q��A8�q�J�^���?PS/l�7Et�B��Q̯d����c�~#�»l����L������0�dIoG,���N��AM��W���m��o͎�B�L�~�������R�r�\������+Ya�=Ƚ����o�p�
�k���WͶ߉�g��Q��H�Á���w��d=ň,&��c�Ǩ�9��ƪ���p��7<�S��*e�$�a�D@B��E٦e�3I�z��9G$F��*7^�?�_|���M��ռ�Z	���q���3�I�P��Ř8Cj��ŧ��L�gD���m�?X}���Y����%�~I�C%6�D�;�{��\��靓X��1�VD�r�~,���,��aF�n�	���[Q��a'���`gB^8�bu�]�O��CV��"�+t���W�$���E��{RTŎ��M���#5�k���$"
�����\_!���^{�I�M91 g�I�����}�ǲe?B�U�_w&�@-��T=nD��L� -���o�"��#@����z\��B{i��8Զ<�C ��w�,mn�3����%+ 	�L�G(P	�3!D!�$y���\�j1Qv��LZ�fX��D���-��Ø�F`��c�GlŖu�Z<7*�*l_�IH�0�����ްqs��eF\�V�8���o����w
�Yĭ�R{�8E�AR��kZ1W�S�Գ�������?��|\h�*~ET���R syi�U_���r+�ZJ����X?b�A��yQ]7��e>^�˚>���ħCP!J[�6��21�s�2b�"�q+��s��XV0d�m� ����:��;8�hvx�,h�7P�;���'�VL��K	�� n";�J�+fy@���*˓�鼽eIX04Y�D
�3+`��2ir�� Ł�fW����f.>?�0��؄(��C��B�}R��h�m�fY$�Ƿ�SӔ������|���_C��/˳}������o�j�O�F���6`�4��ٞYׄ���7e�y�2�@�N������_�O� U>�UC:4��M��&��APe��*ߒ3��$�Y�!8�����0��y����Z��8O/8�G��^��/�ZJ�_ ! s���ɋG~,�@4GɆ��v����D[�cmO�8'�%ڼB�'B��H�f�͎����ܣ,���u|!g��c�9��|3Π?R8�X9'=��g4>̐l�,�e{a�>�`��r�_c��Z&jW��&�""ցd�<���[Ң�?_h��,�]�PJ<y��czϲ<ou��0g�c�)���:�"�<�lc�z�JZA[M�3h|�?ĉJ�r��hQR�������'V̝o�ȤE�,ISレy%���;�p^�^��A�"�,���X�� ���s* iAv�T�I�1H ����#��
̬�A!]r�Ͽ�^(��v�F��&#f� ��(fh4!<��F������<��ʍ� �W��ih0J =���V�jG�o=������ OXFȫ�Tj�Զ<Y�z�l���c=�YR;�8���;�=uP� ��d��Q\����R��@�E���v?![�h0��-��n��������vr�)���eu�hO��Fv��yn�V �`�t�x�T�/�X��F�Ąf��i�`O8"��j�MV�L x��3o͛�n�K�[$�F��W�H��V\�w��h����*��X�'�q?Z�`=��2��"�o����08�B��U`�ݰem$�E�	/����W+i��i*{i�3{���< ,��R���\M����z�F��U��
���ǄU ����:s4M�g�km}]`�<7�u�h2���|����t�{�pwސ�U3}���OJ��;6�?����_ ���uj�*:�ssPv���c�wC�s�}��EV�ma�h]s�	�ME[R}�`B�f����P0?��IG������?��5��1�"3���!�Z��-!f�5�;k+LC�!�֔�1g�&Ðh�}�OP1^�|�\�yiP�&��Yд����X!24g�*6���a���)?ɼ�g{��0bb�e��Xyg�J���a<�����zB?��8�%>&Rn9¦�Z�"�͐���@Wh(��B_�ڬ���
��ڹs�]'����c�����/��(���nؤ�SWY�ywn��EU��9���k�C�`�@K�gAy�}�l�!@���
�~#�vZ�ѡ����#�ДZ}��:Rs�W�����1o�uMĖ_�2N�K�5?[�^��_r��՞�w��x�!T�=���Mc�d����hsg"2��ã�)���u���?�OA�d��)��pOwʐj^�£,��)��j-�F�m8�W���?Wm�V�Z���*5L����[�U���.��FXAp%�ٳ�7���˅LS��b:Ux��r�#�B�F��|���:&�����؇����C)�0/�ʼ���7d��J��HcK"5M��^Q�A��7b#H��~'��f�r��������P��'��:�Ƈ�]��Sޤ��!D\���(I�f�1�J����r3�t��o���z�y�({[E��#�PK��;U�ӣ˫��M��A��T�5�ҽ-$N쮌���7�k9�|X9#OB���6�Er� ^9K�Pg�iIH��t���7wj����x��](���,pk)�6�K1EO9fs
z��B�M\��(/|bT8qu�슣�-2����Gx���Sj�2��Y��",
u��I)O|$⺿g��=@���ΰ���y��B7��.m����*[��\t���{�#\-,ղimu.�@��q�B�p��D�ö�d�X���9<#���lm��|0c]*P~ޢ�3<i�@%�ij�����̑dp�h����H�V��v=Ϸ+u7n����[�,ܲ)t�C��.�!�t,88bI�氺����	'䒣�?�~O3�OS,��_؈t��e'��TA-��$PW�����Y�5�YlFߤ,��2�'�g�ˤ��2�At�.�mi=�#�z����ϱ%D�� v��;	%�Wu�kY�b#��g���T¬�D�ה���yO�X��X(����q�f�v7��n����VZ�m�����q�60���t�˻8�u�����$:���d��q�B���.�fI9�	���d����|u�%]�4"I�<�%�R��r��z|Ƌ'��p�7ZU$y����+�+�3���2@>{)�_���Wx�7��mm��=B�:m"���Q�>2�4����P1,їI��v&����L�H��JM|ۗ&g5N$9�j�K�[���ĝ?"�B[�q!�J��8�:��.ݸ��o�� �W;��x�� E��2v�=ߙ�Rp%7���%e�iI�����^�y��$o���#)�7Ŝ�)�ab��iK>��豤s�{��Y�1?]�{�B'
pb�=жM	p�s�}�<�_ڼ��G�7�e�}��l_?��؛={yBi�1�Y������FQp7]ucEv$�)f�	Kja��6-.�U4]�!��R�o�y�(�91��*lG�bDn�M�^��I�X�E��5�V���7`�0�ݼe��?��\c$�l Ԡ�0�
�1�d����kB���H��$����n��LG��{�6n���ə7�S>vz#@u' �.hG}_Ɵ�9�x=v��9�H����%Z�*��J"���!��,k����֠�f�H��#�q �}f~t����3��j�;0�KO�&D �e��Z|3n:��_���`xK_[]�cr�t��Ř�p��-�e4;o]��8����T�b�mQq+7q/]�k��@�#�����tG+RL0�\�_N�̣� ᖿ�.F���K��Ǘ��Ep�V�"��1�d�R� `Zy�M�9R�������@J8>tG.5jA)%/��9SR<�A�3҆7�@�����:��L�`��+��7��΃������T0��x��Դmz�p딹Н��_���01��4�PQE���dQ�d���R�ݫv:4
O�^��#I��O�k9	�lm>�Pt,����(��Ӷ>�b�"���M&�n�b�E��xE�\���H�İ�&��֛v��!I�Xq�|�HKF��3����,�_=.Ƅ�Z���K��tq��gg����(���^>Ⱥ���b
����S�h"ĨbĚ�U"�1
�/7�2�K���y�E��b��wW��N.�8S<�������oY�v�8�db��c�W:߮�񅐢�nAW�ދ�t�Rv dC�W�H� Drl��^I�<D{���gH��K�!��$���V��	��LF����a�ӽ�&.t�Z=]pZm����@�:dhT(� v�8�nE9�b��`�\��� �	�f�]�G��]hp j}��{PMw�������p��_I�!s~E��D���`<m5��R(̙��kr�N��8$�b�/������X*A���U��jIeU���!�Rv�o`�4��X����U�Gݑ�N���;o��AZ��� s��SAȭy�s>��F\�7�cSEF��h�.���	N;�x��%R���R5yL�i-ڧ�Y�ij�~p��ݚ��YС!��N#郛}E�Y��Rխ�D#=n4�+�M�-j�x�E��ş���r�z�>JfǨ���>lw'�M�n��V,��0{��%�C1dM�n�k�/�b��u�N����(_5;�A�D�L
���E!Mx�m��}B���M1���L�yL���x�pE���\���Դ_��e��z2a����`K���龴�,t����:"N���3���ښf�����KRK�ܚ�;�E�����9]�.�ź��g��1�$'��_`ޞ��ۄ|��{�@G��M7<'>7-+R��9IKȤV����O�d��ң��E��orA����P~�Dy�+� {�c��"0qm�ƤD��j�Б�� �&�>���AپT��ײ�K8;M�Y/�[�ׯ��AZ�J3�
�7�q�2��lc��͋�[2�W����xϜ��12�` ��]Wv?<��:�P��+c��ǐ�N�D�;�nK�nU����P�l�t� >8`��7�&����1�Jނɸ+¢��ݯd���lBh�
K�V��o�B�<]���	
�QK�7��P��WD��S�� �Me���_d��涋����J���
���K�p�/İZ_CB��:k���Q%��`�*�L��a�c�0�7X�'��|����b-
z�ٴ�d:Yt	t��D>6�%���_��"�-Q�11%�L�^���o�Jɤ�~@��`M����"0F��|a0s-*�!�j�Cȩ6��nX�5��7 C%���>��_��;e������q�Q�`��QF'��u+��ʂ�Q#9e�۔�x�m��(\D�qA�������;iI?X�T�H��BE�P��rfb�����a��Y��30��Ӎ	��=莰�t[�4��N^j+b�[��'zut��EՇ	�C�k�U�nc����ʀ�_.���{���~��[h4S:�*ؽ�� T�����rv>�MuC�%z�Y4#X���\��J��=�h:a+�R��,��Gq<�la�
�c��	EC&��9�E��K��4���)rk��Շ�w��R	!��9��w6����y�83�W��~[^�N������	�eIm��p�;���`�Grc�Gs/�L&��||U�5�9���q������F6p`l�`S�	�Ӭ7y��%�y%�wIL=o��u�p���������R�G9��~�����;}��^h_���9K�a�R#�G�w0e'����C&r���D7=�&͍!"wG�V�O��B�>) �i�����Y���d�q�"p�>#��ʥF46���ZӞW���;@uV���F�-|ڎ}J��eomp�}1���5��Yrܠ=Є=E�f ��� q��C�ϒ~/��l���k����|d�(Q�3ýz+'64(��Q�N���}u X3%��,M�Z�4�����.j��>�A��\��a�7�Z}��D1�<��|M�����B�"��K�0 ����z�����*�/h��;U	c>�e:����z�����Ɣ����'C�H-�m��a���V���l����tR"Ѣ�1��r��"�?"fg��?�LsM&T��ݘ��ʑ��`h�c�H�ߴ�~�����}*Fx�5]9vy�{3.�d/�Ғ)i�Kz
D�Dp�X���\��ڰ��Ƥ�寬9����$�����J��!�Y$��ZF�a�/�0���t"!���@i�|�9��>�X����a	e:�VSmD�5Q)�d��H�������Q�>�x�/1%Tn�AY����xc���E���+;���gB��O@�o��M$L�@Hc��Ps{"�-mݩ�2wBԪZo��.}���1E���e��Xqhc���qTo�x��~/"������z_nH?�����ڃ��cC,�-s�L*��~<�9��B��r�����P���E���'�<�]���GB��ŶS8��3���9�J���󺫉�\o�;R�R%_�K�/o����Yk�������.+���zM��6���<�}����C��(7��Tqź|^�.���ߴ̂�Q@GmR��pƃ�%&CFT�:e	�$�A�N�x����͗0�!mh&(�-#M�? '����)�˪��<���	�;�Z���A}�:����Ñ*�{�f������&�[8�w�i��5��]XH5<!�/���Gi���%
>7=��$���^��t�۶�d~���z�9��qj��;�CDY�o�(l.^�@2��� r�8��+����z�z(ƣ��D�����T���v������A�<������"rGV��N�9@=��'\&h�r*� ��]�.��n����Q���t��t}����Xkg�%�P���ݍ�$�1U`��g���+�3wdY`X䞘�%#7��''��/Ôq���hF)Q�ūγzQ�Â9�xt�'Y�A���W�wD�Q4LU�,Jy�:�Ɠ��s�H�+{|x��M��Yۓ��J�/*O��U��j��&$S~p��J�լL(�GՌ�0f�TVl2�aumj�J���4@�V���5���s�����{�n�\�M�>m%�U_x
m7?)v��{�	�r��羥F?d9�,��w�r�J`����Y�g6s&�/2�a |�ssϷ��8sK9�ѽbs�7uҗ���XPm�IFU�2ׂ\��C�l���z���A��	7�V��)U��1�=���i���v��g��Y��J��̄O��9=J�B�<>��V���>2,udf(��"ś�����:��o���7!;�٨��!=�qѤƵ������ۧ\<A�|%��i�颟�!�k�.���h���m��Ҡ����v�#[<1p�ֳ�iki�
�A�C���V�>��5=q%�T������jaCʲ�6p�L�U���&)���m&=�{�b�'��d��qv"����,��?pρ����8g��Q5p���",�}n���\~t�\A�)̗�v""�,��4��D��C�Q�\���
zKfd��[�_k����F��L��R�Ԩc3��Ϣ�Nz�nD��:6ޚ�̅���53Ss��%t�)(��r�lĒQ秽	�s�}���W�)�x��Tx|���� �(�4)?������X��e_���ൠx����A
*�>BAmŰ�4P�����*-�B�,��ky��:=�,(���w���w	t�h�r!Y�\���P#ԙ\�wL�a1��pI�
D�#�{<�2X�?��.ڋ�9e�=U&����,��!�\�$�'J+���,���*5D(��;�i���'Բ��t�����=�JU�a�<����f%N�O���g|GI@�9�GW���=/��~�6�ܮ_���M�<���ՎS���7��z�@�����ZH���2q���Ml�?�H�V�/��O��;
kP6��Pj|�|n�zp��J�r�|7Y@A{W��M����6Ɉ��k������h8]8C�Ɠ��{�j��]�������u>�j�>������,�%����j��G_�q��7�lE�&>�D����mQz���k۝Y���$��:���;/��!ʭu�0ϝy�\�>T���|���Opi0E�������ɒ��f��Q~��>:��0��7��W�o�֘*���y��;��s���o��b}�%�m��@i��`$�~u����N~l|����9}�7.%��$��u�byx(�X�� ���J�����<B*s�ԛO:aX�h����4��]��X�3��,�]9QUI57�9�sN;ʯ���B��ˉ<��]r''���|YG��F�6t���=��f\C��B"çZGvSq�r�+����vs���{� }�p�/�˝{�07_������i#l���F����� ���D���"�ms<Gn�Gp{3�!�ŵ/
;���bCSy�j���w�r3MF��P���)ZPY��3�-�0��4[06�]�@���F�F��S�M]U�V��W��iOVz����Jl�����p�$�}�ͯ�<�E�8]�[f���9N3H&���<h��&�s2a'�+Ǔ�b�G���QtR�-E˩��FH�o��%LZu�L�p�AE=���)=�%�d��!O�r�H��a�J�	�3��
	�B�yn}����Z�i�@"	�D�Rp�gT7h��GE0��buY#;}�wv��F����� �@�]#�%�?�%�7m�����E�q�.����k�A��Sr��L�ʩ��Zם��b��xoT8,O���TM_B�)�9�&w~�ԎǷg\>��r����k	ȶpù��G�x0u�	1���_fx�H����)s=+��6���j'�Gq�-���M��H� �d6�@I{ ���2r��$�"Z������mz\�f\V[����K��;,H4�?�p�Q}��e��Z��$� ��]�!�}ul�e0z~P�A��A4�n]ñ�S4���{� H)	�?(7�V����1�,��]�+�hv��ոN���&�<�x���6�Kck��0�=�����b���8G�j��L�p_�GEY�3�{���U�ij��$K����?> ���N"|��bnO�)�����r�=����G�|����"!��%^*Q��ɻI�q0&c���/e]2	�S5q)��i�E5n��s-��ں���fM�:�nc�\��9�o��냔U�'p�h��)�8���C����R@&T��((�2�@9��!�N���.�D�j��4R�Z/�/�-Y���^,���N�MOi����ޞ�Ibef����j$��_��k�A ��+��_�?m+4��}Zڴ]��Ki����Xi%
�zo�G�N+�34X#�Aqܷ�iM(��i{}a���et\�YCf����T��$3�D�Φ�ӫ�?����:jEl�A*2�$|�aeu]�T'�1�M���=5�t��T���t����.3UR�S�P6[���9�Ll��� ����Ř�3�ꍰ������أ�#_r���M�o���+J:���S����Uh<�?S��j�pG%l�[j`�At��( ��^z�;�����*��N-�O���(oi��f�ǈ��\om	sT]�2KO�7z��E����0K�s��5���m�Jvf��E�|�YO�]��@V)6����l�����ݦh���n5�݅-�-�z��Y��ƨF����Cc>HV��3�t}\[B�	�L����������fY=�l�&�)J�����Rp�c,ԟf6��b�)`)c\��L���)n�(Hx1 �.
�yQ�l��屦��m�B�R-=R��U)�h_�龔�:$L4�0bA��� 7�-	�j�
�A:�6���~�g_�48�7��˞{]�ޖ��t�zY����U|	���l�V�J%�l'�N�[�c@��T �?Z%�ҫ �.�3��CH��=��'����M#d�|��:|������6��Z_\��=����>�"'����0Ϟ��[��%a�x���@��:�
B������Č�´V���r^�2Nsk��b��� ��Ws�'�z+�$�3<a	�C�w�G�(�O��уw�Q���&!��M�@�a���\�3w_GO�v�I��������z�){m�F�K�oz�_�����{ ��O�O}�v5��(�2`v@����O�H��Ձe��r�tr&�|T�$�bs'�~�pWr٥r����f�=R��D��	��w��d':�����n�L����KUۖ�:��G׿�k!Σ���L�I?��*�8v�A W�s���ϥ��8	G����펯��K��6�}k%�4V� 6*
8��tY��VGB��h�|��*K���+���~��)����ɩ�i�"� ��g��X����g��9���?ig�A3R��/g0xh�&a��5��Jy�-	�)iƽދ�?#@�<�1�T�1���@��rm���0�j�/����X;�P��y��Uw'��e� �^�W�Ov���Q�T�&��0H
&XQ��]�< 0nN�Q��vx��������T]o���!��zƏ�M�<h�e��Q�wf�ID��*�ؙ ��Şs��jl�^�,�A��M�?ʀ �8x KKd��ۼ����6vl0���/�\��
	�hs�Xn�k�T���(����b��w��L=⺭��NH�
A�42g���b,�<�Lˣ�V����y�(�"	(:�l&��Ά��>���<߼��B�
vq$�o�������l9��, e��9�Q47bD���7�ZF�x4{Ur�c��TMmGz'��L��^�%&�U*�Xc���Bޡ:��8���=Zr�(^g{��t��+5�r��s�Ns��V�#wZT�6��u�*^��s�K����1�
�t�U�(�5/4O�mDW��A��]g%�*f�J�rzo�\�*4��4��j���E��:���������]WM��,ێ�m�F]�k�P�����	�Yf8fv�ւ՘��j�n[-� )`g-������Q�"�8�&�-���Z��?�ʅ���<)�����Wl5��&j3XѼ��ឈ|[Ϫ���>�Y�VKn&(e�]{H�ŖK���k�gF׋H?Y?�[�_�Iܵ�}B��d��\���	X���J?������Wc�D��vy��sݺ��B��~Fq��>4�Ώ[]d?}�P�`�9�h7C*z�R��:d.�O@��rA�\̯y#S��ʋ���$�NmR�
)��tazUxKA�s�����k`/�~aGt�ᣏQ��z�'��w>1�����j!i8�"���1_�9��D��r�Y�sI�<���BW�W�?��]$V���S������(}�h�}2_r�"7�]f���3j�3b����`}7�n��l�G��3��+E��S���\�e�~�L��Kq4�P�*���'as�U�H�A^�n`z�e����[�#"�*𛿼�$���:��Nő���A,{�ۨ�J9�rFY�$�Z��E �� w�I�y3U�4���_=:���c���X����-!���d`L|a�A��6�@��65'+)IN�0 r��A$�����7�z~����8�9���Gl�QMk�H�n�Y���Q�^���KsdäK!���窓|���T#���{h��QC���!M��<m�惂e�t��HU����>q��&��LiH�39W��k��p���A�Ґė�8���R|$�din���?^�҈ό�(]�;[p���ر�X�k��۬��%[��`Z$|�\���'�%a��=�ɓB��W��	BL�����ʰ��ڙl��b�H���Sȥ-�$Dw�de�Q
�����&p��j1=�\�g*޲G� _���5�ﬗ���9����B����B����ej�����,>u�]%vKlbZf�Ҥ�x�Hλ�&�Ǝ=��x]�5j����:��T	��T����ΙE�|(���C��F|\z���Nm�u�z-�����~~�/j��.>���i�o[��#�F9�msi�y_�9�G�X��	y�8����淖G�'h8f����T�� ��V�5ŵ�e�(C3�[��ĪN#м#���f�= ���]NV!��[�cTc�ȯ���d�-��!�ڗ�G ����UFzh�t�����j�ϵ"���3 �Ɣ
�{	��p�M7;�<N"<����S��U�j>oF��+R�Bv�����3TR*��DA�ސv��_��2x�d4K�/z ��rb�JTozO��v<Y�)����q��x�o�UǞ|:�� ��_ �I&VC
���+nyG�ib����򥁑U�\,���>n;��sl���w6�7��\�g/�B�74z��bJ�z�+�Ra����_Q��
r��_3��#rΞ�.8��ut����nL&�j�5B�r��]�$���yM[���0:$�R2�f�`0^��S����LZ�2i�����yBM���%>�gTaT"3$_�8.n���#K��4;��}>�vݵ�q��1HY��� s�&��|�&��5�,W��[��U�%WAG���u@�e� ߫��~Q����z�Q����R�19�ہIH�D���s�� 7��8}	���x���Y,���*ٜͨ?7d��l_���X�
�U�7x
���LۢGܗ�&6�T�&��Xdnr���ƚ��v��r�A�#<k�<=ݘ��?�ZH���&m;su�s���#����1��!"=��&�9�4XY�%�{,��b*uG���X�T\}J�Σ��W`;�)�7���>��#,��Z�8ڵ��%JR���uh[��5��V��}���%d���1��53�����Z��h�|����28��Mw<x��;D~RjXg�`������0�m�jţ_@a��W�K������s�������O�0�R������J"����oĢƾX��9��V��/�.*�;c�����ZQ�l�Ƅ��m'�^)66��N���콅��)D��"o��Jz;Cz�������K�s�:�?tt�R�/qJ�J����K����'�Ģ��"}]��ꚬ�v�����|��8�pQ�z̧��m�$:�0:��[�yQb]�2�KE���՜A&����Qk �B��l��]�fB�-�V"�� Fd����BGbj6���u��C�~�]���������z`�W"�>	�&����E�$=������R��; '5�h�m̕u��~_�%��ƿ&C�-ESz�����I\̞���S�W ��fa�&\�`ve�Bl�#�37���Us���R�"�g����ނt�������@I��Rg��51`�ˡbxR�A�'u i��������Ha��H�T�fJz���;\�����$FN:��0��r�O���9�1=^c3�)ʕ~�	��c4��9�qT$�Cr�$�����@���Z�4�aRD���N<|�(���c�I}> �ϋa���GS�3���y����H�F��\� �Z�LJG�	���ˬ��
*	��9d�$l��Z/��
�]�L�Z���4��u>m�}�/������?�VYt���O��;�r�7�Ĵ�S�hO�e'�I�K��a�h�9�)�(l�e�A�}��z
��K�޻�J�[=��t"�F�G�z$?���*n����G���\�ͯ�A���Mu1���fryn��:�������U�!Ee�YI�J#*E�r�p�����E3e�
���iB	�k�b�7!�:a�����L��8�{�vX�p�S�Z]���qh�WTB��um�8��]���|	�5�p�O���V+�\��] ݋�W�~�����+�m���ߎ�1B�W�O���&P�o�=mu��* ]����U���]��L��}���9�o��g��6���֩Nx��y��J��� Y;,��o�H��<V�=GlE5?�H��Ȥ�ؓ���94)|�ѡZ-ʱ�H�7�(����^)�~NPi�ڔ�di��;���#.�b0�O�Ώ���]	מ�u�qѾ�z�ٜXu�2���z�1f�ˎ�,��W��2<�Y@S�`Px���H�]#��h�g�t�$F$�/����U3\N�'�����؄���#A8n <mKX=KEK��ѹ��Em�Q_��9���!�Z*ښ�ّ��`�CM,4	/�Rr�nR�UU���,?���ϓ���ݗi��=-�K��NdƬ����?UI�[d�e皠�2AZ�)NI��3�c��V���E7�'X�q�ܶI�:�_�4�����ӭ��,�s��J��#_d������כ�I����Rwٿ�@�PBK�FN~a)ǭ~	0�?F������`
0��n��,zˎ�w�:�Y�4
w��0aEZH�;���Jy.���5_*ņY�4x�"J��_0�.������d�-��:-Z×�@g�le.:�7[�JL�{��Fh�t ��7�8ɻ~R��*�d1�����}��d@e�aV�\�w�NBF��[�#Z���%яHoY���Y��އx�#����_�F�F�Wq�̵�+L�"��Qͦ��9�$�޵��Hn0�`~_��U�b��sH ���W[)D+��>5
��3�ދʒ��Tk3��+sY�۟_E'����ʄ#l��Z�W�rs�
�� ��U�d�*Z�;��H�����Ȭ��.� B�-I8m/{����8JG� ����Yz�H?z�8
�ZL̟�W���u&�9;����Z�M���#���<n|��K�L�\���-D�!��16D�{y��=@l���=+c�W$��{�t.�A�O^��;da��
�����bR#��e� �8�b��0���DHkK�X��+K����t)
�+��&�Im<
u\������w��".�������t���rNMf��LB�Y]!���cDE\��_2�5J ��� r���]a�H[��������m�6	A4���b��yP&�N���u^Fq��u�ҏ�iS����U���+^/:yR�J��=�c�Q�j]LP�� �w����蹱���v?���.��)<O1�$ټ�Aݒ��mT^��6�����ѾL|��a?`�T+?)�3C6� d����ꞩ�x<vOD��d�Hm)�.��Ym�Z/����'��X�L��X�$ovT(Svn�_�w#�As���?��7��~B���6g!WqU4�������Rk�u�{�ڲ�	��r;����;I�{5���� �~�qͯP��b{��5�������s~�([f���ڇk��ɜB�k@>���� ?S്���z(�	�ݩܸ���	�����c���HM�����y��G��B�C�Ć)����c��bO�l��7�VT#�US+�g^0���R��{���"�w2�%cf� ��!�|>��{XUD=��z��45web�y���b��,��&�;�m�Ӝ�<���%���:i -�!�n=*F�BB�ד���7����`�\�k}���2ܫ�z�]C���bwqj�b��t����^�)��0��8��7җ0��������	6.U�|:L�U����'�Oi-,?Ol	\[L)��lX�
��u���U�D�)<�z�� �h���1S*�$[�	8����lv!�JF�j�����B�5�o�Ƞ�]9N��߄.k���s���Y��� :#�i�����&k�^�A}Пd~-���c���N:�^��P���Ir����Wf��	m4��
v�R��W:��t�(�Hȋ"1�(Z�_rH�2��+)����?i��\U܌?ttR�� !�;ϮU�Z$�4��+��*���-��Ɔ�2�T���W0S��(�K��GJ�kI�'y�锼u���ҙ��9��� "�ߢ�!y�Ld� o��, @Ы���f�~d�n�n}�ݝQH2�WY]��&���k�Q~$��Q�/�i�R��j�C9��/V�����|��
b�}�Z�Aȅ�ZR~�J�
8�Hν|�^�[�`"��z�`{�B�@Ui^����_2��C�WF��P �����%�|1�I�/�J�:����O2rL��~3�����7�����s`���ub�E�)����e��t��D��u�Â��1��w`�.��:�V�1L�|+�|�ב���L�@e{iJ�{3> 8�e�yYߣSq�^���靖]Į�6�K;�F����?3������BJ�qUW�'��@G�F?���J�7&;[�#��	�U�[��6'��,w�`P`riƼ1FHy[7�� Yr��]!���8�X5�x�}I�X�]AMA�Ym�G6�}h���Y�t�!�D]V��i )�C&��&+�Z�tNW߆l����B���� M���ѹ�w��R�*ԫ>���H^�a����������N��{a���s�怑�~�4Z=�&�}EǗ	42��ވ�DN�Oi����4gO;:}�&�xQ��Em=듳�0�i��d��r���	��oO*��e���Qp��˱'���G������.T�h���B�I�KeL���Wm���ow����h�E�)��p�ů��q��R�Z*�ܚY�:q6D_8��=e4[��l���I��<q&)�v�<k��t�F�~�0;�õ=zG����NĨ�J2Ք�WI��[I���ږ(�0짥�Zxۅ�a|r�B�I��*D��o��a�{��G����O�� n��[�*��, �X30ƣʽ!�6M�P��,�;���=��Wƭ&]��zZf�'_r��&F�"��-�����r�o{-rPQM�1����,N���> `�K,|�|���!�[=3Y`,"j��Ν[糼��9�|/8�C_~'�M[���J�s�&ӁKr��u�U�	\����&�;q�q �B����� �? -��F�F���>M��w8�!�k�l���%WN&������(ӎ��<(6�,��S���=%���:~���]A�VB��征���A�r�o�v�S��$Yw��Y�㡅�:]��ā�u�>���Xz�@s>���|K��򣥟��-��,�}�zLZ���~����U� ���m@�y����"�Ղ���S�^����^��}��cn�: v�_���n��灣&�A�8���Z�:���&�MշD�.\^g
�����N��@<1����� �9�qZ��buw~���`�/���<�E���맱z]�S �V՟�, l���ou+�r�3}ZR.��a�!��b�`���Wh�����(5(*o|�~'�,���|��J��<mn�O��/~�'\&��OcN%PU5�zI(fV��}ʣ�������2T3҈�i囉�L��$�ZT��x��&-@�s�ه���q��dɫ�񫐃5�S����yZCr1)��������=R ұi�
0ڽ��4���~?��;R�r�b�J�E�cg�;�E���(;3/��ږxC%�9_�&3�u��.��)4 �*�Ϙ�x�����n�az4sr��wl���,�&���7��Z��nF�k�ݓ(/U\��ҽI����hA�҇�p�/�~�h� ��[�(xjĨ$1��_Խ=�E0���w�	un��u.F�7���j#��=Hk�h���i�t�V��b�Ht;����1����(�NB	3'���ڸ��tc�8�Ow����w��ې�_)������	��������Px�**��r���(m�l!���q�)���~5����@��  &����Y��W�`/W�9��r���.K�cbV#Z�M/nii�2�&����(�J\2�"����,�J����Mb���zGV��U���?�ԼBHb��p�i�/m�
])�K�3��]4�Bo�w��<��Lx�.8Nc@r�Zı��JcB(]wK+���4�yk.��,�,BN
S�U~�w��A\�Ѡ�f���N��!�A��!�U��r)�p@�8P�mvu�x��]4��¿��/ʜy5�tnZ��6!O���!�yD����Q���Bz�i�{��=�����P�𨂊'�Ql˃�q�gn]��:1��Z� *�	?�:�K9n��ZC�/,Z;1v��|.�O0�9`�<�!�;������i�nS������N��Oٴq�<߬���&t���h��a}P��l��!�1N'ٰq�e�
lΓ�����R1�CeyY*3-�{��ڸV���Sbe����}ϱ��G\rW})G�5$i�5)�&�$������,������ S��P���}���[��f���a"c����9t��$l�N�m,֬���[K�C����u~���C~j0�:��� F}�#�.�2�82hibOx�k��T�ob�QDv=9^{{�RP�-M�L����T�A����֬�łx��5'v-�c��|�ե[41���{��8��gT�~�Ne3�4���7�����4y"ڕ��Rk̿����	wv���-�ng�@����c
�������^	A�n��1D�Ӵ��T�E�s0L�LO�� 4,<� A�*F�#�� ���HN��ޜ�ٕ�/�ሧb�'T_�ߎ
c�e�������-&��V����b�{����r�KЀ�e��3�e�Dk2r@��>���`��R;Hc�F�b���w��Xe��J���f0��	��"�w<�L?�f�3����5�ruj���g��Jl>#�� �o�������5��S`U	>�}��:x'��mv��{0c0����Z_��A�N�p�Y�x9�6�U8�f���^��:w]x�˂�����4����pd$Ҋ&�������p!,�
	qFj����QHt����f�'��RDϹ���c�WW�E�[�չxjr�XRF�� ���
�!� ����HD����Db�;�������B5����#��{���fy�%3�z��=��W�U�t�-:����]�~w���pniq� \q!��5�k��JL�d��A�[��B*��~�b.���PULX��e�5��s�&���J M�C��<5z����[�h
G%��"uTWf��d�	�u�3��y�2A.	ј���z'$ꀣ�]5'*��̠,��k1m#F��dhJ���$+y9�껫��	�˳Q~���K?h��E���s�'�f�{A\�@eW�������f�Ib����A��>�O��P��E{�p^LMm*c�˷��"�_T�ax�ߐ�O7&���k�+��!�tnX��!�! � ���أmz�P<��&�@P�����#����KWެC�(�D����q�9�x�+� =� lXJA~�o]`z6T~�5ud�,�=cG'S� �7-���[wѷG�Z��cE��\0�/c���熦=�H�j��0"�Z������ys���p4F�%j3��ڢ!�o^`GP�鋝�)&��p��v����ia�v�ԉ5��(»�=���VF��볣Ѭ~���(-��SS��E�� ��߫��J:�$8a�7���KqA�LB��@F�{�FOr ���]�0����W��Hf5��6������\j���Ŷ��~�
���O|8풦��IM���,�c��Է��~�W�<����ZfZ�XB�š�כ�.x��;g�g�/E�hE�k�j���Go���LÃw�l&˧io��t��B�ms�mP3��,��/^R�ЬN��/4KM��t�m�/1��b H\��𜨛|'�5���m%X�o�0��R�5	��u��wu��Z���n�Ug��	F�k���w=y�<���K�̛rT�Hc���-����M��;�0?pb ��(��r�����3�;d!3�1o��nT.�Gn֘] ����F,G��X�_o��Ӎ v�����iFt�6*]O�N�����	�>��B�3����O�r�f�R��`���j��XVV[)tͭR͂2>��G�2>T߽�����/��ČV�������� ����}YB�n�p'�(:s�����lљ
���fxV<J�������G$%e_�e��"���Ԛ��b��A�Nte`�a�s�?|el��Ѳ�)��yzf9��?y��q��l �ئ��7)'���8�n�ٞK�
!���T��(��v�Rȭ�JN�,%ך��R���@��%:E5^sG�ҩ�Y"c*�@�ׅ�����U�������l����)B=/A0�m��EODӸ���XO*�	&Sl�����4p/_ٻ���D�V�keCh�Aٓ��a�t�RC�_�/G�;�Uƚ��T��Fn�� �S�|��X����4fo��_r�r�+3�Cɤg�0�Tw������bx)��/q|��(VS[��Q��1���ߊ��:}���^���:�e�@$ 𩕦��L��I�� ᔎ�<�%=�]�0��^��"肌���T��af��+��$� =U�3�K�	4����gmJXw��|�`3(WX�k�o�D�U^�oM/|��i�Y��BN^����x�#cxȅ�)�?慥��P��,4.�&@Cl��K� }�7b�x�
 Cg�]{�n�?��X��B�Nɹ�ߨm�ɿ&�c]��vf��07<U���c��QؾرI�:��a�GU'�T�B�����Tdן<ouV�����|�㫋H��J���{�RKK��|�h�:���/F��Ciu����z��?����ҝ��c��`l�;�m���Z�h/���=�J�ʪ,N;wVU�9�����)�U�WˑU����i�Jh5YOj�Wz|P�)����y�����������?f�i����y$�}���*�2����X���[��\��J����F�C���w��꟢��(�!x�'� �]�:���
����)!5OBhA����d&�ZrL�lm"/�S�����ü�?b���k�d'_�lX"f#�����
��b����}"�񙿅7	y��� ӭT�ֻ�cu�x�g��B���Jտ<�x.��!ךFs�	-wS�I<G�+���N��ǽa,a�6��2>��7�B�%*7��z[�ށS�R\S��t.�P�;�H&�02S�6�ky������� �퓐�� ���3v��U7~��څ����QXM5��jx���� hCXy�Ɉyu+e����Q(���Q���
�
*��G��hH����#�* �Q�M9��/$��'�����t�aC[�=�U@?7G?��p�vaZ�%a��Tq�)�v�����rX�O2�L���N\1Fv(��&��2lB5���k��C��D�Y�kbX�A7�|�{!���ͧ�ʽ/uK��ʳn[c3���P4�0r�8k�t����:V�~��j퍡� �38z�%PD��6�5�Y�%:(�B����l3"{^?����A���Mz�$թ���k����#�loԏ��v�l�����V���r�|ؑi0���۶[,�"�A�|\%yrn�����jh����n�����{[�v�H>� ?/���5��GP��?ޕ�7�C�K�]��lo�2�@������8-��e�?�[A�KL�����k� ~���������)o�g�de`�t�?d�����E�&�{e�K*ǒm�u�!���ѝ
�uxq��:�k�
t�V�,�R_3Q����Θ�5`�����N��� �Ӣ)�o�pܪ��%}u�{7�|���o<��S.�.�XT�q�֘��H��O�����<k������@d�d%
1�f�h65�խ�Oe���1�Z]x����#��]��g�=�m�����r#�Al�8Q��Ir?����pZ�Q���TbF/�T�݋��,�bJ��v�R:������@�h~��],RX��
	�Vj���	�H6��șҰ�M���Z>��_Z�8���OZ�gNa�t���8�n���n<O�&B�96US� ����(�m���{�tA�p�E����I� �_x��ݗ3N`��-;0�ʃ���OǷ56S��*��'�t���Xk��i�	s
Iً��m(�j��j �89PA$1 �A��[�b�rRM	��3@�p\]o�5�ߗqd?H�:n��rFm�Ol�~���_��n��yXFbuŗ9��D�F֋Y��U�����L�p��&BF{�J7v�a|��W�AA���� �#��p�a`�WU���Ut2�-��5	2=�ʹY�	cMŃ��v���ɼ����Ԉ����X�z�%��
����p�T���HG�y�E���S���$�b�L�p1�"l��'3���'�0ӂ�5�F��~�%��,��dX�p2S]���y�k�*��s)ĽI�.����7�4����"M,I�W��u�U�4�ZVdk�-�hf�T/H�WA�NK|�����ƛ�~��+��[��6&9�G�A��ɬ�8v=�����l+^��׎��3&6��`�`�*�� �U��fx
{��O���g!Ġx����4�#�^�����0��e`[��Z�.\�6�M*[�.0	���נ2s --~ܲ���˭̛ɢ�'�D����G�2����Օ�N%-�憒�����Nlpb��b�c"� �b+��,���'����6������6�Sq�ѐ��Z��z�秊]گ	,�s)@�]�q74W�4&���e��)���'?iqr��S_��[1NEZ�Z�`�`(�Og��NX�|�=����I�Ud��L�}�[4�U�X�����������$rb�y�U������T��0����$�4XH%fsZ5%nCVY#�� W�/I3ҩ<�|z}��?X�q-��`�.=�%�2����#�,C���^�+}��KL����՝��1�
=6v=�R�d|���ת��碘gu��B�E���.0<.ƻ����������m�9�{#�A��HI16�����z昝���[���&�����<��dE��̵���g&s�0�OE[ ����: L�5��~o�WW���A?˦�>��g0CSp���<!�Ǔ�6����z��p駩Ƒ��n�A��=���b:b�Y�����#����o���0Gfiܐ��d�	�P�G�n�R.@A�~11�]��D�pڬ�h��� ��<����>.�#��c�>t���U���_L*F�^�k�	������6�,�~bOp;�D�l]^n��e�
ĺ&�"P�{p�i���I+CE,%�.��|$���7A_9�W�J���1� ��֊��!TrC���e�m��5��(��8O�j����ร�2[���"�{�Z��r���)��k�D_������������R&ڈsU> #�}|
�fc��p�G��#+ii#���9�:}uh�m�b�κz��YSn���۱�����_|�h��Q�	g��W��҈�ӔC�� �?OY�������w��㖅�����%9�}����mL�*���IzC�ˮ����dX�$�N�	�����E�O}@{X�x$j������h���uuSjO2�-[����DDY�I�:/�Ļ�Ղ�т/U�@7��n �%k�S��x�t|�!qM�u�t�R�[��������gp���"�WO@Q-��$_��x�G�t1y"}jUO�i�����V*�Bu��(s?ymƄN���Wg�'��|[]�FQ�RQ{>]
�Ƃ�M���u�og��[��4/h
���XK��A�(���qց$�@֚�A���?(Q�.�׈/�}i4I)Ǳ顦x�wk�ڒ9:�`�]À�FLs��yzG��6�Z嫑�|M�G�@���"��nT���?�;=�Wҝ7�B��Cni`�l�Ђ$r���׋sƶ�4�bY��:���$�ޞ̡�U��eB`�WU��v�S$<�cW��;g{7�(>�,'�ڠ^ &�cR	3<u�75���R����lug��h_		b×m,�����||����;�<U{����0�,��
�`�n�1#�o�xLP֑j56���Y���Z� �2��t̐�a�3�G��&�U�~{$(^x2s��W]g�������#��9%}���D>�z;OS�f� rq�T�k헤�0�t����򯂎�K�ԥ[P.){��Z����4"CO�"����|��%�BX|���[Ɣu�y�9t��ߴ�"'V���+�G��Z����rx�k`E�Z�љ��.�2���H�h`�����[�f���8@(���툒Gi}����(� 4N��M�!��ק�DJ`�H3i�C�܊d%H�o	G���Wp�8
v��c�9e�lD؟��K�۽�6�d@~�4�	dW�� ���Ѿ��*����Y�D�����sE�&���jY+�A�)������OQ.b�8����[���f?#z��W(-b|��S��IP2�@�?���W�H�:Q{)�7�X����i���R�{���sG��W5t��)|w���p�:ݍ�T�~���'"��&���u�iA<��O<�a;�c��oD5p�;�S�4\�Y~T�fPC#�;l"�j.%,�q�DR������@��Z]�@�m:hX�^�}�� ک���v_��������xO�k'��  �i<l��J����*���
{(��Jm�!@�Z����v��H�݂2�k����N����]��$�����X��*z]�'��fr��4���:�qxǢ��;�R,�U��+���J�X'�B0����":^A�.a 7t\��}�H|���(Ÿ ���L۬�%Kb�PQ9a��M������ú��#��=�i����*vm�.���z���杄��q���vB4�P���o-�D3�I���p�#j�2�H|ͯK?u��͖L��	��
���M�+"��j��{N�����җ�,og�s� [i����琔��x<y��ؖ4���v�Ξ/M�/�Nk?����0=P0]8]���)L0?q�^��>H�iʲ�|X�L�PÉC,^�2��*Ey`]#:6�	P���e7�RԷ�hC�����-�B9u�
V�`�~��<*���]E�ɜb�$hG"f�����ϲ`��@�ϳl�w�Ə�lHXSol�y��qT��M����MF��WsLvS�ik]����5C�T�e�^�_�n�n$��<��j?���x�K�{�w��Û-(��.��"�Z��p޵��ͯ�/_0+����N���,1IoPl����&S6��~t�1�s�|@!��wSj��@�ފ�� O�/҈?\z.=��^M�Jg�nr��	��F��k����@��J�٩m�p��[f��~OFH�����޹�B��7�oe0��V����?�Y��P"�2�&}��h�"A_O��>�I���)9��X+�kl����W���׌K"<��1j����������꛱����{K$��x'���|Z�����a��m[x��q+��OZ3����|>,b�%{)A�n����#�yN������J�4#�}LE�PK}�HLb�1<��a[�q~��[#��<�A�U��%M�a��h|�@C=��POL��\[)���G��
A����aPh���C�L�4�/:?Oi���;44�A��R �����wXQ���FJ�L���p��M;]S�ыXmf� �K�*�� ��,~&��5�̫�4�e�s)PjlEt`A��'W9' .�ĭI�9�[|6c�����{��_Bg�wm����O�U+t�8[=�m�UG���(����ޱP>L��J���>]C`/�i��]�诎�Mi���lq�<n/
|���&D���%��}I+^��Nf@����� �����ԉ�3N)/������	�o�?��V
��oN[�Ӽ��|�5�;��I���aP
U/� M;l��S6���Ϭ���>XBB��L[	����ehz  ���F���j���S��*3�l4p"����)�4���2����QaE�:�|fn�g����`��_������
�;�����t�\D���S�7:�)�:=<?W�Xb<ɧ��ߗǷ �3eoF�l`ޥ� /?ku��À�x��'�o��$^��7�q�ݫ�`]�z����aaD�C���۪���^}Z��l���t�o-dĶK���C��tc�L7�U�o'�9���g|��}�'�?���eQF'Gt�Jn4�@n�����}�A����˸㟌�~R�L���G�s�E�� ^��HC��y�Q�8�$/4���By�#�Fc,K�mm0���M#S���1f�
o�b/��/�|�V?��uO�m_!ۈ�����|@g��=%i��/�+�'!��u>���L���3W�����(�Jwcxj� o�w�x�jR�oΣAqGF�M�&�f�#��1�)�T3_�<+r�k'���Z��������f�E�n8D+�-Z��n��%���-BZ�'�7"kհ�?�UB;�.�F}�.��,�U7�����p�ıf�� }��r����Otx���n�!r2�V]>j;A~�[�N������)���]ԎT~�%�|�p���.e}O^@��"z�����o�Ki
)��,k[d�E�%\e���8�	{����.�~r�}a��5��aG�~��d��0�΂ fh�Xԉ_�vH,6�@^Й��$�r/V����I"@��jz{ʐ�4��ɓ%�۶`y�d"�<��0�',{���J�Rj�^�m�6�2�U���|�gc��� t	���>Ӌ+�R���V�ܶ�Yp��!����t&�п����o"(�jg����VP�0R�~��,�U���I`*�;R��Eӷ��;/�pݒ$,-I��XCW-���CQiP���ˋ��X?�����݅�B!��)<p�HT,:�����ՙ��NE�/n��f*�F��ͽ����M�p\m�я���DÝ`�(�U$@�c]�/��b^QߥYV�6k�t4DŁR�M�(>�����Z\b6"R_���ޱ�~~ب�V@K�Wz�lq�6ϰ-���޻Z5��W���4dg�|<��TnZ�=9��J5s��g!^#׋�
����=���{4�
�|��R�Y��g�rJp~U+��
\:�O��/���v�w7	Z�?��X�k��_/x��0ż,-�fk/BՉ�	*X<���4z��c$w#8Ot�9�d J�}��11���iR�Y�&�"j��b�C��+J���6Bi;lt�����[��ϩw��2���"lƧ{���miw���aݧ0�B!q(,�B7!�?0�3����b羌�/�å��F��X���HC�n�pa���B��y��0�B�=�Uֹ�z	�,��<��RM��j�ѻf��vv*`�~��kQ�oT��<�a[mV�LnB#������30�Ћ�-�"�wo��^w(��ddp� �V����9���?)r�=�7��������I�<�;s*K��]�_B�uzA����BP��Έ��<BYv�ήV-�f���ҊY��	xF!��R�(Q�n;�;�%�q!{x:G��'�(8Y�m��h��*�L)�%���}#/����CԬy���
���U�$��@�@_��J�;��F�P��ؒ?w���(Q1���f F�^%�K�b3�^?4E����o䰫[�����ғ���P�{��?�5��=�j��ݦ�N5i&�\E�%��!	g�]ި��đ�MW<�U
�x��$ѕy�׾j]t��쀀�\����-xD��v�#e��<Ea���1��$e��А��� :5r�-6����{N4��&]��(W�~]����e �･��@[	X:}fϪI�����5��ì@��.�qJO-�Ka"s�&()}�h񌀺���y�ߝ���*y�l�=��<ޔ�ѥםC���>�%ce_-a_ޓ�7���͙4���_��p���}�j�W�8��6�5 `��xxB�U�\��J4S��D�\���2��?{|���i_���_��\F�>�}�n�O����q40������<G���PuQ4�AD3Ы�*`�\�؀�m4!md��{2M`���j�⛠�Qj�0/�;�>��@r�F娺կG����>�R.��S	��b������B�I0n4�0�赣�#��@�)~�r���X�?��b�g
�Q�b����¼�E�����ekS���+`h��I0���J�)��jD�L��-�n"N_ח�l����%Cq�,o¿e �Qr":G9�}�\�[*�o�2���{W������7!�ݳ�D�o��
%	29����>�����E q��)7�`�i�q~�Et�K~9���6߇���ۯ��b���m�iШީp��a�!�rq̊>Yβy3���W�����q��I�b� �&�����0���1-/��D�i���h/(�A��_4�R�Ւ��iBе2��|��.M�,"c?�0�RV6[�+j�0�D��2����藉��������L�n1甊׿[%ăE&�O���U��n�l����' ?�+t�$Cy��]Ȭ�3D���Ү���@[��:UQ���P�R>��#��8%uF0'P�p�H�˪{�D�i��E��Ǐ@��1��ӥ1��|��=��w�P�\"�B��lH^}���L�A=�}K�k�/���%	��'J��}M�!�ׯk�Td��g*����ߖC���bx�������M	;���+�R�+-�G ����U&?��[����j�D�o3�Yn�11/ ��z��.�ؒ�6��'Z	���Un'=^��>ç��T��21$�,�� ��ە�:!n���)k5d֞Y�G^�5�NN�xa�mK:�G!&��n�y��1H�\?}�N�!���X�iy�h���
�cQ�6�bB�ҋ�rki�3:�)1���n�H�x+�ȕ�\Z���ի�]AB`�M���/���^o<������m�=���u�cN�Y�r2+u���)ep[�$���-L�yj����d�a�&a;����S��//�!F|���䊮#.�p[���6��U:	D�*�(�w��ige�L�n�H�q���Z�֭?0��|�	M|��l9����v��v�fB����cz>�W������������Z�[��� ��10*�p�(3X=pX�~d������K���)t�ko����q����"W�25�إtA:ѣWՊu�v�kӕ\��+6��f7 ���T䵬%zl�v֢�e���#��^F��Tj��n���&dv��[�D�<̃�К=��1���n�D��H��I�^�K�⡥����&��v½�,ywXiM�2�+w/�F�6�Q��l���J+J��w`ز5ﴥ�+c���G��Q:e���M�F]����a���Yk�9y@(��'�19!�#M5$D�~6n�;H�<�ǜ��yx� �a����� 1-J6�ld�3ւk�m;|y����D����un�=�%�.�RX=�����Ɣn����.�R�!T$i<�i���t0Yp�ޤ��"�;kg%6�c�kd�����1>c.��]��͏��w��3��]����=�@�X=�4�X߭�:���.�寬��V������ˬ��:���m��[��10���_�ùR��������~`�&x�#��b��1��=���W�Qs[���f �هL�r�z
w���D<���_��d��kV�~R�	�Z���rIKd���p�L�-��jJ�G&M���L�YWx��Y�ᩈ�e����$m\�<�+�x�6OB�lE��<�e�,,�<�ʈ!���S9>@EImQIb��mp�4Gt
9�g�% �`��J�9U�h���>�l���j)�&ڀ�f��R����E��`q1�4�40��Z��&n'�IϷ���p����LC�|Cs)kA�cb�d�Q�/�Wk��&�j���=�=�ս�n�����$�x�m���BX�P�A�1���Z�?�m���Odf���P�εF���}#�A�:]�+�T�IX��լ�č�"�eR �����kX*L�	��Mn޳�� �PmP�%��&,.=�f���L������C�+�JeY.���0�q�u��L^�}ԫ+���9)?�n������6�`��6��lz c�d#W	GF��YCI�nF����\f�:rMĬ��W���7�������PRƨ7�	D�Z������ߞ�R��f�<�0@��OH����j���H�;*$�1�>^���L���dQrރ i�4m�o�7���SLz�۽���h߈�ֆ~�>�V8 ?F��3[b��8)������e�����4�}/��08�m��� }q��%� � �HxU�+��h>�Y�k HR�޼8���ht��X���~S'�c���b.7�s.�3�Е,V��v=���(�R�Y�;`ɴ����̓���MR����ɢ%��韛�����c��X0��g�~�Nd %X"�
�~+R���_�{%C,�>�-1nprǦY`і�tp��h��d����A2�C^9��$g�֮��H�C>�
A�T$z����n��\�F�~���8*�F����a�8�X��"����Ǿ9�,F���M���O��6vP��K`�q޽�Y����Ғ��̮���tv#���[
5:�<����khJ������zy�-��7�e������-��g�α�5�/� ��Y>��ۀ��Y;6SYe���[T��8M�1�ƾ70�"0q*�����(M�Y9n�T���&����V����]�	J���c)qg&�^��K�[��n�����p`�$KZ
�s��p�A7��/qf��ڲ0nE}�<�zI|pM�.ȱ����Nj>V�sME���Đ���殭���=m���#X���1.₎��4|�A�쌧�1Ķ�5+�)�NE����������9/��WQ>��P+>�=����:Ia:﷫��d璣c�.v�Y,ћ�[@��T��q�!I9:���)����8���՝�����|���m��gB�`R'�[�#z�ߟn��s��#�7j��_�j	�ءa�٤���A�Q�[M��:����o	: %�c��%���ʔM����_PE�[����ȁ�IVڶ��8l�`PS�9��&��ͳNX*��hN�kT+�] �z{zf���2�s�cg��A�`�bP��-t������}p7.�}�8��pLo�� wW`��6}�ն�3��"�Hi��� ��������.���,���S��0f�F�۹4�R♎��]�Rn
�u�Xu��vXH�A��=�ƣ�h^f�$�	���/��i�y=P��}S_��h��W���Tv�({��0Ҫ9�e&4�R�j�}�*�w���|(��]�Ag���h��*i�b��G$�"�ٳ뺰}�{6�W�nى�^	M�rw� E��g.eU7T��y�h��ӻ���Q�K^��=�B��)�v��\�Zʹ^]��+n��/�=�bQ
���9����P��kI=�]N�����}@�و�ci솪$8�R3��R�5*g�'����5�XB��Q��hTB��SQ��Wq4��]�f��x_؄0m�ݡv7C0[��gUn�r�<��~_�lL<������1��N
���g�@����1�Xƽ	C=��R:�s�"�Ҹ��P���1)��Y�}k�l!�a��<��sT-12�t.f��S+����ju63��#/U!�����ఊy9�co��LT��!��q����$�(e%K��;)@u�RۥM}�Gqž7��+�$�-�O�Q�HgHkvQ��������]���x���9z
�CsFVg��D+k£=y^��F��־୾$;x����E��?��^��e=��)'����8w�mː!�T?���xc�/�A�I��ߪ%��
IqՇ���k�ڄ�����)�Q+Lx�����2�����ħ,�&��ݔ9�K3s�ʝ~�t���l	�Ms���.�<��}P꼼�6�zX# l���n9��B-y-��v��Ѷl-$�(�g�f�ξ�n���8�9D�JG�Iޮp��[���[�����@~�Rô�l�f8�j�vB}�x�)���0d[�1��Ñ��g�F�I�>�_�m�����Y�pW��a��'���T���E=W�����l��,�R���=�}A��fz��K�"~,���;����xݎ:_���5�|�_�L7]�ʹ����tS��-��JU�?��n_���2g���Y)�tӓY���|���;�9�� :��(�n�5���u?k}�w�"^Ͽ�L����"�� #U�<�b� g���1@����O.P���MZ�����T�!nm;��^�ot*РV�*���,��z� ��
|W	M��0�.˅Gf�eF��Ȓ1��\�������-<g�\�����[ZE�-2�@�u�fvv᭤��L�z}��Ҹ�1�Q2j��D }�����{�-<�m}�g���������909Q�j�P�2����d|��[o������+k1��q�H��ԇ����zq��E*��>=�V���t�n�9�T��T�<��Rt�f���pxhg�tv��.�Ko2�Ƣt�$�9�2*�a�F��!��gB8 B�h�C�ؕ+��ӿz�v�`7bxA��L9,9q�������oU	^��<2?���^cd�Y�ßFfKe�|1��U�.�PI���
�d!��x��.�%$��~�-��C���X[\��~�q*g7]�q����Y��5������4v��`H^b�E�x�ދH��o�Y�/�=��?)����[��R]X'�W�b$;�$w���l�;J�!�_�lj���i�[���������L�D�Odt��9���:Z�������!���������4�����g&����Y�|��1��ӈi��$�F"f��g���v��"��)��7r�7:�rS܈�
]HV��)p�S� �f;�{I;Q��^r����E���8@�,�)Jx�R|�� <@�!��k�pu<a�$ҡ���0R~��@	��𮥒3�
)k/�-�]�$�T\����'Ġ���u?A��W��5d�R�|�/��Eg���+K��B�����&�����^���Q�Ea�"���T�jN~�ٵX�a�ݐ$w&���΋�PL��l�-���"]Z�p�[`��Pmg��)�9�k֩��Bb�~���L`|��j2�g�鸓�6�MK�Hk��gl��տSƄCy�	`�fl�^d.�z)�}V�][_;	�k�˫�2�'���5�n��h�imUCY�|��Rs��د?�0�HJ�L�TAJ��c�7���D�/�h��T���t�VK+ �d�j
��^�$��Ued+F�X�|�yם��̀C�0\^�I?L&;��ND=c��6�ws�Q}hxV�F ڷI�Q�&	�)�:&���1�[4
�'�T�����r[�PF�~7'��$�VE6wk�e�x��|�~-B��n�f�ѷ���}F����K1z����{���چ��JzNZ�b�AX@�R��j��=�U!mWp�Ml�����N�ۑbꩌ���|Āt��-����\]ɭ|~Q�%�E"�%���08sy�*U�.�lvT�����.�Qq������!ښ}PW.ȼ@��x���/�W�6k�gY��Ӌ�y2J:R��?�o��c��"�)ߵ�}�qQ�m���`�_���%U���V�B��n*#�JS�gO�b��7J�/��
��nȶh�)��-�M��RTe.j����?����3��G��4;���D��a��z77��a�����4���r�`��%�՘8� �0��M/�Hۿ�K�5�[��u��*�4�)�o��A �}�����3�}ؤ]�b�
."4Ogh"B�6��$���D�z�1{�3��Y��;D���\(�w���z�/�ڦ�H8���Ĝ	����t�����6�sa,R�IT)�@ʦX��G�����p(FLB��4� *��p���� �#��:]��\;=W)ў�gH����溰���r>����pa�2����X�#=�����I�,v"ک���m#�<��B�����g�>DY �"��k�}ZM�|��u��OQ]�L �)$ �x ���Y����1��E)���;�}U��d��nIxn��~B�
](��u~4����Ө�cp��֚'��j�SE��c���)��r�*��R�:�<ϝ��)Som�E�Х��_�g����Ћ���5�q�����+�oB�`S�o�:^���W뽔�����V��X|����JD��uM|�����Əq?�����b�I��r1�N�3u~�D!4(���� #�ȸi�@���
�Ĵ+3K�Z��3�0�XS8�h��+&]�c\��N�B�55&�P���L���Sf�*7��&��^qL,u���d#���V�w�ë�;j��������`N����*�ʩ۪O�P8˙n��w�b*z���{��(�������[U�P)�-m� Eh�E��䥋Y�
�A��*�z�ss	|�s�n�k� ��:z����*���H�����h���T
6��LH���R�9�'&n�fH�!�����S|������u�We��V����c���SKe�XQ�TOc�=]+^�r0I�WR�
�މhŀ�B0mc����m�'��Y\�نsO�����2����s�0��Ҋ���;��O�>���X��F�-�4I�zd�lA��N�ZJ���/.�Zۦ��x�6�Xݬ�c��}�c�@)�픘��9��c=�2�DtG�la[��΄�\F>~�S�|�q& �����.4���`v�_z"Fsj%���J�ן�z��q�Oj~�C>?�C>��I_�Ez2�k#u<<L�߫�az8�a7S�;��w��GG_L��V���|By�ۆW���} "�4��:%�F�����M���+���^��kefp7B��T3H���T����^��X�dņޥ�6	���FaA.�����a�.���p��cG���o{_&�G{�(%\���N��_=�r�"*G4�S�m~y0B�p��B�6�7n�7~��ݲ����%d+�J�Q3��,�>�e_��:�ÔX�Ek������ѷ�QF�)0Kq˛e�.�! ���1�y���hH���E�*;i���m�ǏF���`�e�Ȼ���bB+������7�����;/��(Q��82	��+h�pFQS���=�U�
�Ǫh���34+k�f��C�X96�K%gyp���ދ{�ז&�;�	P��ԳhŻ�#����>�
:Y/U	2?K��Qzr�N]s�t{�R��͙GK��<;M�i�����=P���gF�d��륆)��R�3����6I��US�v��q�3����>�}{tz¢&,AtF.���?:���9yȏ����1o��)meW�����𞹰��qF�l�>��gO�˻���h� �C �l�lG�e�;`Ǯ^�t�mU��@��Gl�q��P0�+�����/s帮Pޕ���MI�"a��]B�`�3F�n��J�����!0g��&�N����x�A���U�Liïp�ģe�69ëC�G�F��5��fg'$����,���O̊=�� -tsbp�
-�!��}Cl5�n����0�m����]�Xbe6/�4`�uP�N
D���1K+������r93��DƔ�����T��V�k�Tl���l�U~��@Br�k��1�+���:�Ć��j��Ց����z�Y; ��.�MѢ=R]t!?�۰�x3��=�p�$Q:7;���2Jr)��Lj���lvw��g���L4����$�Tr��o�^Gm����W<� �#�L�;k��K�!hP'�����5*q������7�:x�&�y)�|�_�s�V��S��PԷ��A���Cgue��] ۛ�g���0����v�*9|߄�|�b������,�B�;�����0������,�+��e��=�V�� �lR��h"�y�>�uݮ�ߩ�!̃\�_�:���PO��H���(����r>f{e��}� �K���r[v�g�#�o�+�:v���b��c0M���S��e��2H@�;Z��g�lSXY�A�<��|2�5�`��Ap:9���D��ng��+yaw�>P��8cv�+����Prȋicw�>��
��z��Ɩҳ&+P��]h�7܀iJ0&7�|�b����[N�����4ȉ�Q<��C����~��)t{dyq�/2�[#n[z�ro;"����Xņ��K�*���x�o?�^�5�HU|�f������Y%lKok�r�Y>ڄ�>P�)"�FN���b�_�*2E ?��2ba��ʼa�WÜ�o��M����-�?�Z2��31ﵽ�Ib<WpHCƪS���k~�����LA!$��M*C�����������y�'����ݜ��Z	J�"��O���P�m����r�$����O2
O�H�
��M8����,�	����=�p6�iS���80&�Č���>��G9}��y�fuz%����J�����7^��`i����̭;Д]G�6��s�N�>He��5�)fF7�fq��Ր���V�!��O�AY�d�&Z�����#��C�
��1G̪�	
��2|Wg�#X���qa��|�|'�]k�b�vN7�� �7�l�~@�_��C��rM��8�s.<�V�>Bum���q?�?���?�2��м~��!�X*�la�@����hTn4z጗����u���~���5�{[se�>���ܨ�Ћc��Z�d�
�!������jp�0��j�������g�^e��WD�#E䡨�b}�[��Sq9	����p��h���1k�	�B���L�3S*��o�~u/˘�G&R�v�eL���!2�t���*��pS�c��	�j~�{=���ۏ|x�ײc�C��-��E��.�/�A�L M�&o����#���:j�2�zب���(�K촹�n�/f��fќ)�tn�W�#5���V�`ƒ�$ʒ"�y�8.h�*� ���Ѭ@!oO��4�� �(����t�WA���w�Y���$Q��!��PK����=a;����Ȑ�O!��YA�*�I���F��E�x����Cb����Q!y��}nP�[ �뺦y/ �ze�$� n�r���(
7�wF*|X�e�ͷ��n�#2\�C����sc������.GM�8-�
���#mR�(@�T����B��?9�KɌ���u��' � dM�g�$._�����e�Q�b޺)ΫO'"a��@���0�ա L�j������c_�`�z.CK��엚��v��i�@��o��-�*W�x����(�%j�gjz��۽�$( "ڴ�����rFݪ�4i�<=B�>��R�� ��[��[Ëj��b���������8v@�<?(wm�6���r�jg
,Szc(r�Pb1���� ��ȴj�4�2��jcbʡ\��i�*�qs�>��؊��0�4٠+C��%ٖ�-��hY��S�S���&�4]}�y��`HD�����e2(��ߝ��HY[;���Dr��G�fiâ
y��;2��)����Oa1b|A-O�y,�C���"y�M�KF�W5�=8��P[�kn��(�.e�Hc���V�9�1L^="Z>����̝jRj�j�ewچ���ܑ�ʪ�Az�'�2z~ipr��:�}�Go�*�j�e++G�B�3$G�Ů����&2Zp�D^�whX���3�"3�X���^)�&/q���_o���ܒ�
,��(�O�`�J�y�:�(E��Dq!(��^Χ��)E	X�m����fϧ/�@�y���z��	���V~��{~�\Q�;An)�0������y����m�*t���l�#	��REN˘�%Wk܇�{v?����?Ȭ��#��c�U�+��"�@&,O��P,DhlB�_�w�9S.c\���� ��9S��>CȎ����Fc���ߦ�wiY@���J��o��㬯:��Z!Bp��咈�I͂k_����9��oP:��%�.�>%E;��#$+8�0���a���2�)���h�ގ��' �uj ��@F�i�_����(R��1�+�R�9ğ�U�E�.(��t=�A��:�3�R~�o�c��c+]Q���M�P�ԛ�S�!8�q�!����nȭ ������������G�875gL�7��(�	��.e����{s`�S'F.i��|o��+�l����A���kГ*�A��F����°��7��=�Qz�^�$La����J\гz�Qc �r����tF��P����H���V�qM����A�+�lD�9��b;�ԏ԰�����1F��5�|I�*8��ɗ�<]�^�[��J\b��B�Aj��)��L"e�x�0�bd����#9������oCx���b;�3r��[I����eH�*�"�]$&�G�i���4�,�&d��Q8��K��P�e���S��-�'fZ&��H�0�0 �=�S��ݤɆ�������GA�u���6�G���v���S�T#��	/88vB����ρ�TD��,�E>��!ִސ�9(�O[��.�(+����z&b���w�}2��Ȑ�Yz�8A'@��&��W�L����.m�p?ٙ���(k��7c�+��e�Y��ު���Kg��ӮY���@'GD
�~����:,'�)%l�{H��& ����=���k�K`���7�#�U�������.n�^�Z3��G�R:�Z�oBU,:����"+8A�_Qp95�,=T<���,Pn� ���j��5
���F�"��a��:0ea�#�	�_��nmu��L|N��T�E�ߦa�q�.�E�)�K��E����R�9w��H>%��2=ƣ�E�%���d�m	��ؿ-�A��K���p����GOPa�2tٌ���Y��ˠ�a%��Sy���0��lg�/W�����7	݃�;�ܵN���;�@�I������i�x�,D.YI�޹ �P	1Y�Gi���s��E��M�^���!u��W����T�.�4��hB������雉�D?`�*7:��F��sd����nzAڶ5&T���~";.o<!�2x�g��>����@�|/�u�����������w����(A�E\T�k�DЏø�!�@N)}�e��W��?��PP_�;�U�hcR��C=[�f��U)�X�I�k�_7 Hryn��E�C_�82�k�B�I�~c���zm�&_�Ժ�Q�n"+V�[\�V�!�V��b�~�i��iz�ǋr��k%؛&:ҭ{��^BeA-���9_jX��[4?�1��X).R1�vX*X�(3&�v���h�c[;�5��S�⽆���&�(xOV�t���,��R�?n|��%�_j�T�N��Xa���$+`K�a��������ƍp4heH��'�Ô���F�i�l�&۴|b&4IU�}GD���B=c�Z�"�!V2/��}�]��M ��C�5��֔�·9&7����}쥕���,�	GU�	RR��aA���dnd��v47�^TH��E{-a��>P��B��q�]gL%�Յ�)�����
f]^�AT�����4g�}�9�� ���1[�"~AHK�:�d2���A����I�`Z#4�4,~������)u�k�q\4}��(+K?�;�Cc/w	�$k����2���3��X�Ѵf�G�~����C�-�ҷ�]�v�,ܝ�A���%��� ����8H�}�ˉ
�%3�$"��w�����!�p�Kub0�lP��0ښ�l+w�D=��L�m-jT�M�wM)u]��X���+;{԰�#�����P'�%��N溰>��8������^p��kQXd�$p�K٩e�:�ޱ􀿋q-����h��[�n&����_�N�
,�ޒ�Qx�ij�i�!��S�Df`�s��1*��S1H�Ԯ����j�b_w<�Y�9��E���9(	�/��րĂI�<�?��.q�Ň��kV�Q���s�oɴhܘ<_u|@$�:1қ��UZ*��;���q�W�~��8ɨU��b��w�K-�{�\ ���"��&0�ߕD���[�n�g~I��oh���,`����q�#���g��޼p���C)�F��UF񯨦������>��"�.5цU,YXx��d���!<[3Va1��	���m�����	
����H	�%� ld�~�iW��@��������o��)1o,!�&s�P�7�/�@3ۀr��R�b�bL�����u��ywk)'��B��9��m��&�"��L����ѫ��<�ҵ�L-�.7 ��2�F\�9��`��V�\���eW.���rS|���ӟW�#��|�Q�����S�gI+S��T�����a���#y��]IK��u����=�p�ݥq����o8 I�{�^'Y I��º$����r��,O�PoԾ%z��c���y *��l����ۢu��ҽvɓ��r�h:�UV�ec���`�� 2C���=�D�-�Վ��2w�j��/,'�ɈQ/��`?���@�K��Ҍ`��a�(5��ў�Z��7��v�J���6I�ƥM��U� ^̾l�I!�QS�Ƀʣ����qHb�ؔ�O�>閳"P����b~��0W,i��G��]~��@Sar�5�֓�{��Y������1�(q����s��#;=qU.p�6�BfB�0qU��K�w3|�\9�,'�t<��Z�}���j��,���*�&�s����I bU�ks'�S���� ���cFo�E�}jY�� �re���K���u$d�ͼ����;D^���:e�c1-�:ܺ��픉9���A3u�̍�C��w�hAI<��47�y#0Xѹ-wxًB�����"���x��c̞�&�^z�C*/�Pl
�	1X�4�h�?�SȽ��bQ�!��m�h�PBm��/�3DS�}�z2�n�l8�Uy����@����q	'#����sG��(S�mU�3��S6��`5�di�p�?�hB2� �D�Y9DrVޣ}N��4^nœ��Pⲏ��Ȯ'�Z�G�����p�Td��S꯮�Hq��/��1�[)j���;�abe�s���	P+����j^L�����xK�c춇`w�I�H��M�$y¤� �f��D@s捀9 �c��n���:�0ă·L��:���St�P$�|�Ú<��{����f�mT<���h�m�IUgP�����*�3:�����d�������D���q����o�ڔ������y�����	����{IH�{�/d�R3B<^���`D��p�S�_��fX+5f��g�q��_4����~-����z��h!�É�&�S�r��G�����c�t��g}��Mz���n�������M�M�g��imH�C>������U�n
Ԟ�On:j)Պы��(��?,^@ �="����1C��O1��������g��9�4iִ��T�J"����H��%�z5y,��o}��J}e��)Ӓ��1Y����h�z)�o��/Dg�H�uS�+xsׯ��s
��&=��������_�`6��p�<�6( I���qK�B{��M�ֿM�i0A�#����������F��i��v�#�����Z���F���#���o4�,
/n���8��&���ډD��f��{Tjv��?�[,#��q���CQ=�|A6��{W��]cL�|�`���-�����Z�^��P`Jpy�-�V���ët���f�u�����WQJ�2]迿k������}�����^1�}�R`G�8t�
���]P�lY��K�P��f�����6���}��P��*���z��a;o��7�p δ�~J�]��_6|��*�����w*��ː	I��II�ʾ����b��/_�}N��?U5��;��(@�*=܂�<c@N1xp@�ƣ�шQ:�_V
 ���5ҜPǯdv_: @\X��T�0m=��� ��Q�9Z�c��$1��Y<��.�{F����s��O�yM����B���m�C��1�j�=�U���]���u6�wT;ꮜ��h�s��a|y}{�ss�>	���í��n`ڝ��&��zA��
�����j/\��m�>�ì��?X���U�?�A�]���k�+yԗW�����T;i�'D6>�<���i�/���x�rH|7w���*Ȼ.E��vY�̝��	]f�~��7<���` ��-�+�C���Ԍ�_ʔ�`)%A�6>6�D �K\V��#;`=�^�Q�b��F�z�SK�wm"���֡O�s`�P�K�W�8,_vsv(d,M4��<_��KO�t�]I5*.�U0�$.�M�+
�yx{���ʜ�XI�x�/5g�E_ϟl��b>���0k7����u�f��i�=�E��f��ݦ�W�$s[U���sG��W�DT��{x�n�����g	��8�����ރX�x��,K�SN�v����	�iձ��`[.}�G��n��ETr�6����d�
%�FT�ח�Ԣu��0��?9%��mz"N���y��1�k�F\64(FE?����C�s��@�T^jͮS7���Ej���.�+�{8�����¸,Њr�u����;p��.N^��Γ �i����P����a��Ϫ��V�+���Z?�8��]�
sG�����?ٓc .h^��|�&ߝC�%�+��٩Ϝ�9f�	�^;������vX3Ɖ�P�,ūy�rl�X֮gy��JGH��X`����"(��ͪ�^/����E�;SI���F�d5�KBq~���QRw\���`X��~�ψO������_1�A���yy�y�qG��V��)]��I��H�2��(L��خ�S� �xv�a�0���B�h��w�ћ�}d]-�ji���)�Pa�����٢�Ĥ��������i�es���0��ʺZ�./���.0��{!c�����rQ�G����=)[]�S$ZUy���{U'���N�j�wR[4�?�������?,������[\UcI�� �y�`A��֍(����N?���Uݎp���=�YH0V���ol�kZ�K��v	B�"�v�[\�2����6��s[���]l���N�#}d^8@��"��J)���~h!��ݎQ��J�������̀&M) �s��fR���CѦeN�|e�]����R���2��|ްB��E��	��x��|��}� �D먭&1�Z���7G�D���s��h�P��o����¶�ų� x�; �E-ANY�Nv����0(��>�$v�Vb���Х���a�������(^�_��ݓn����������F���g��5�D%ᜲ��Qu���.�g�B����}7E
�ԇ=�ˬ.[6��9�]���S�	�a�e�����Sm��[P� ĬAN�W�=�ha���$�70���k|��_O4��}|�b�y������7*�U��54id<�;�����h�LIϟ^��M�솈0�S�?����z��uPj+/U�hO󵎲X��3����M�ņ?4����� Q6���}_C�B�5A�<�_�`�ڴH �S��N��	���B�NCCpL��;����:O񑍷b~�=.���Q��2�a�[d��3��!��QN��)����40��7�Z؍q��й�\FlY�ZS��є��9�!q�G�w �]o���%^��v��ϻq����h������}�tҢ�l�U_�L�×�,E61N� QØMֿSW<� S���X���=I��.-���[��bH�y���N,�AM�Z�L6M�p�2�%��:�g$u؝�E��~�1�I��g*��-u����/.�!]r�����ނ���Х����ڷZ'~$,�y+�����.'���G(R��^���������b�x%��Q!p+e��[�m�j�� n.Z�sS�z��@F��C�0���i�uw�&��'�ħ���=�}�
L����f�)��4N	С���n�[��|(��Y�&'��Ңq��[�g�=�۳���'r�g~�SU���9=Ym<�J��=p�f�b�M/f��My��[��|C�-�`�0����u����[.� \�i��I�z�,a��p��d�F��2�0�*4V8g#{���5t�|�Z{z�P/r�̕w�	@��f<O�@fc<������
�Q��mqϪ|)�H�8��uN�#�$�wt�:���é���6�|�b�#c{1����kU �i�����)��Z��>��q��l@��&����w8>�۽�I�H>\$w=&fE�`��v�p զ~�DB�1#���Kk"�䢔�;JK���O�A�2��XE�+�&��>,d}Ɋ��<;��z�f5�ƛ�1�+�^��S�M��}A�?C�B kЛ�J�[a�4X��;��Bm�mC�T.�]f���H�H��o���c�3�& �&�a�'LQ��-��/@���GŊd��&�	��Ez��/_��*?�{\d���=����Ԏ�Gu��=F��tԼ��('�`�hz������B�+���AS�O���k�hwg���ӵ"2�����*j�B$;��H�QNǳճ�P<ڒ/�����+*4-;�I�����js�m���ݠ�̓�2 �V�^fޑѪ*Z��ѹ_-m�<�@��K�(d�C�E���k���-���W�d���H}�y�vñXf�f$�U��W� ��-@@�/�W�-m
<���i�/��H�������bG3�24�l%d�"�����*�W:-J�4F�˶�Ǉb�����V�e/( &0����;ڥCI2���X���ٛ��,!�I�a-�F�Jj�~�D�l����]%{�i����jv����߸> cv����!�IL7�ƾ�"�Q��1�8	�ٗj&F��Ŵ�
ct���.����%kڛ��jw�T� �O�.;��W:�;6p��وz����ko����DP9�'�ގD�t�J�{�:���QҶ��F��kO�>�Czu���ՖK�S�ô��b���M���,ʫ�i�N�N�0��-,���(������q����;���q;۔�3瓽��8��7�YyZ
B�y�Y�H�8�+�^�;wec���m�,�����~��4#�d�s���|�W�p���t���˓!X���䝟�lsp���[}�;�Df�hiB��� B�_��a O�j���༔�&���c.�d�ڞLA"�������z�r|XB^�L9�%���Bbq4���=��J�c��aE����;�_��H�R/e02|���7{�38��L^�*:݄6z*V��~��a��Q��%��ѰK���P��/@"���i����5�վ^������9���hW������06���BYx�q�@�`S*�3Ш`���,���86,&�}�-9�4(D�4B0M/CC�fQ�ܸ�ϗz��P���܄z���{8\�N�)��a��M|��l��F'�������>v]��y��&��A�⑯�8�@�МT"�g3���
	L:\ޏg�Q�Q��j(�|���<�`Q��A|xboa�A�n����.�豳#M�]-���1�gmc`���B�H�FeC�@2E�T~e�]	�W�p�����Z �ef把	��Z�; I�r���,���:=��q[��Y_~:�NB�D�pU^.۳lua��{�9�_N8`�Hލ��'��v�4)m�g��e���M���b���@���Jz9�}�N?'���+)4Wl�[Jy�hq�:4n���Dy�I��)Qm�v��"JTxء�;��5d6�*Pb/i�{Za�C�J"� {�����ϻ�ܿj1����){	'�:�o =�C���ShG�b��Q$��Z�_q諕Qdx{;z �mȓ�ڱs���7�ϰr�,a���Nj����%+��!*ـb�� �`���p���>�� K�,+��.�}�MQ�ӑ�I[�f@�����_������$�Þ;��Y�,tK04��I�|�/���Cpou�`	�+H�!	��ޡ41�ئp��ֆ���,�h��$i`c㜯�s]l�$ґ���M̖�/�>���l��������U�X��WT�o�
�.^��'��8S��U�S�k��[T�� �
'�j����⫬ml�sjI':���f1ϋ�����i��8%�5�`r:��˓�;$$g��94�=�6��;�{��vԘ8��C�N��ˉ��@�[.$�����	}#�'�dܒ+�bAaYc��V4�ǳl�MEKΕ蝪�"�A#ڜ�o5��c�Rꑀ�$���$��O�Z=8Z[L�h;�r;K] 4���ܘFeՈ�+����� .G3]�3=�-dݤ�{��L��s���|��NӾH��L�/D�N��Έ.fZ5t4�
#�|���Lh��W���3�h2]�$���@.UNcZ���>�1��vU��x���`�'DZ�s-��s��x��6��N�ޏ�l�D��E#fW+�*>��"��zMo�9�;���'��90��������2��Y1�p��:7S\y"\U���\!p7j����-q[��~���[��x�G�z{@���>Z�K�oU�ާ����!��1Ź��ݚ���DL��N��z��T�b��+��*U��*1C�� | �=�����SW�^���%.��nr���P�� /����
l�#�"���_�C�q1�k���ƪy�8l�%;y*�g/���TC�rM}�5m�N��%Ps��������y��U��� �E7%�$ ��2c��bV@d���'p�*6���0��]͋��P��.4�_nXN7T���c�:�æ��nsb������1���ĸ�80Ţ��]XO�`�*Ǳ�"���7�j���5�9��	$�������'7�6��,*\<�-���c0���7o?�E�8{̍�1:ʘeN �]��q\N�Si��:��nk�"��g��	�`�mdx�cvrs5Q}f�������4�l!��QJ��tq�J��$�Ր��Y��c^��1���P�8���h�
N5UH�.�!���^C�<~���pe�ႂ�o��7��c2֥��� y��[�S;j��w���$�"���� ��8�sj&�'l�~;�jN����;�P�hkG���4	ʶ�t�ڨmk��x�9�[���s�(�9�
ڌp�@�{��IA@_�.�Y��4��˟\܃�C��A#���mj���.����1!h�v����D�׊�wn���%���t�k���U�0��#�W��{�W����@#Ko��N����w�Ċv�[]�}���o�f /)�E�g4��r0P�T�y*�Y���0�RX����y�6t���^ʏ����q���RE���"�kWz��Hn���ϋLj��� J⑪=�J��0RJU�1D���֎��w9~��6c���r~��M畏j��o
e��('y�W�7��MgWz�wYΨn�#����̓�3�}���[*�\0J�G|6��b4C<P�"t4R�����je��y�Z/�2pc������5U����U�>��Qr�:;���r�<6$|s�y���g�"0�7���?�˟�}D�?x<m0|�a�����y���$+_$����H��lQ�Za�������H�`�E��A���1	'^��2P����>Ρ���	�4D��|mڂ$D�
vz0i�]��4<a�"ݍ���l6	�*u�d:�t�Na�Rmj�x�Py�����qe�M�� G|A�� X�B��#BK�.��o��ʬ��� L�_,R���A�3����.H�S�d�ɠ^��^���-�{��r��ll<��+㚐�J�S|��������B�,�2�6�m/22��*��e����.,�e%&���c��{��f�k+�T���\[زW�����IQcz�T��׬Ǡ��=�W!^���5^��$�}<���������%B5g������ri�~'\ߧ�h��q�H��D�sж%z�нQ������O�3 ��I�b>R;����	'�T=L%�������w��>�K����l�c0!al�u,-�\�WgI�>��@�c�5i����~�>	zBK>U~ʛ@NK�\�Rw*R��E��l��4*2�B�Of��un[�bPR�í�F~�}<���� Qr?����S�C]偎�[(�� D�ț��v�U�ET�����d��7�E��UK�v���YS�UW�d�G��������{��gY�^��&/H?��!n���ҭ�0N���z����|�ʯ�҄BV5�W�V�HHFl�P�=D� ���Κ�ǻɵai���R*����*�2�QK���U{z�����|��y#�#��a"&�� �h����,͋�<<���5z�w���u:fϳ��8���k3=�����2�c��Rd���~�E���})!����{��vd�'Xv��N�5R:���+F�{����j
��/�B,�OZU@AG9�b��/&(�X���Ү"�	@�>,N^��l��o��뢷����?��d^�K������*��X�cظ�D�ߚD�#���m����B�����j̬6�)�p�9lZ�Kdw���5s���3�B�� ��2�0˒����7�JK��)��L��n�o�A$Gy�{��r4M����Ng���Q�dY�@b�u�yS��2gh+�(4- &Öɨ�:�;%�L4T��:b�lh��@�N�I�L�t,L�����#̮�A��E&|Q�[����"��OSA1��E�&Q����3t�����sm���e�k��־ɬUv���>|aG���jͳ�oA�e��З
FR�7F�母\9����`1�x/MS�����+�Ò��3FJg;b��J/�H�Nl��}���v�Ewv&�}J;5f�}VT�E��b�4���ח�����v�jOÅ�ˠ���F����n�V,)@��u�� IK[�����s�MA�	��9��=�1?ӻD8���#iR��x4�	`���|b>�ۘ��:܁iۗ��j���P��-\�a��^�yE��Ţ��L6�}��jd�Qh�
�;�4�T%'S���5�]cʨV^���IKu���0���m�v��Vp�sm��Y�����>�+��N-�I%)fsDbN�aP~zC�ͅ�~��������sA�@pN�u�9FW0�C̉�@Z�j{��.��2�b!�{��l��N�U}(���"��G%������	���7LH���a9\��<�E�ă�?�*�~�P_��G�G��\7�<mN��2Q]�)o;�ۅG�����D�a��n-�/�%�ήʣ	�����E�hEp�]�c�HC��ub���S�K��,n��B�Ze0r��P���#��-E�U:���K�4u;��S�P 2يX�B�Lh�Ln��_��� F7I295w�T"�Z�^��0�u�/	��0�͑V4T��9g�����c#��	��F ��>�:v��A���C[g�J�i)Mg�HRz߯�\I�1*n��T��#~��R6�~��t:�E�M�A�#$4�]+Mɕ5��������p����"r�1�����pt/��ZF���e�-Ĝ�+���J�Vm�����j�kLh`&��nB�r~���
N���Z�'y֤oxa}�3�%�Y�a��f/�=>��[�	���-L���M��	Ty�y=1�����X ��h:0^jf����s)#p'�lG�����XH@�cCBI\Y���2�d Pa��g[��HHm����ǯ_%2֛a��.�^�a'��\nȪ��pV^� ��걚	_��ϝ�-���a<�.���|��Z�@"�����v��S���.�
b�$Z>ȶ)���?��s�L�PwM��ĥ����&�ܹ��`��Z��S���;�1+�\%�++���&�����u4GS���Ԡ������v��:�>�~!}Lɂ*���z�O�k��k�\�[�j:��y����(h{��ޙTr����~@�п��;\\��ïPh�p�"���]���fΣU�t!"��x���i�iC?홻K��6ZlJ�]��p:#��P ��hT�"n��������~��;�*�^������N1��֙�Ŷ��)��b%����a�/�(�"n#:�u��aK"۝�F��b�����{�.�7A!ܒd.�������I���8O�O
)F��U��!ǂ��ߓ�a��$P�p�JJ�(��ާ�f�Aiq�a}�ޱTޗ%�@%E�v7<p�F�J�OC֮+�^�T�{B�o�q�4���|���7A��t���=�V�pߦU�L��i�ҽK�;.8�P���X��R�ø���ס*ѯ8�`GA��r�ۗ�����f-��Y��vv�J�ڐ���;���� t�#Q�vwI6�G�_�)������p
Wh0��=G%�a�^��W>%P�T�z�,�0e~ T32��.��R�N������8�2p�������{��+i���A�p٨�2g��΂�^g��a�Y8?�*_��T�o�SK,J|4?�q
�G}����W�?$�Js��ѭ�$��}�0�� �G�Y�����0�ɄPY#,�˭�$�y�/��=N���8Y�1@�g O:��3���A�i���ZE/��iۚ�
���ސ{�ӧ=s���3B�����c֬lcv�0\�7���j xQ��=;g�K���<���12���;��gz�C'��˜���q8��~@���nl�	��ŧ�Q멬����Dj�?�^AP�����i3�U�hx�,��u�SW��c��#0��w���9�lQ� `�y�G�99x�9��^?ۛ��mznS�q�-a���h_��AgW�K0�bYX߿�"=��?���;�/�x	��d����P���b贒Q��z+f�1d�5�3����L�´-6 ��o��>k�"�8F����S�nZ���Օ���{c�	��Ţ�,?���I�E�h|�}�]������8��/C˰ހ���쓤���ҽ*r�?ϙ�v�$
�����Y}	�� _%}aFA���<�l�¶u�vX�%�m��%�yao�:5��J�������*��5�񥠫��p>�`���4��e���'�Fy`�>��s9#��gp�2�d�'?�/@t45ss&����@�e�]W�Z`2e8y��$�A&�3��8�VUGx�*9���P��а�S�A�Q�u=���$mf�"w�n�V��x"\ȈR�o�y�m}Nal�����s"���S�����n����>*�c͗��u��ލ�)?'��t
�2�rѦPX�u��$��տ/O@��S۾j9��ɋ_��&;dMw4N�����i֡?��蟘X�B���!)�����|���-4�5�pĭ�Vfurͷ�@�����]KR�TL�2[�C���~&.63eP?Df�r�|� �ef��!k����\="�
K^���+:�i�>�����BEeH��/�{+AD�)N�o��0~��sU.Py�+�2a�s687��Ǝ�*ǿ�]�� ��}״��]l݅�o�{`��}�o]��#�m%Wѧ��U�M�K��Wa߿����Sm� Y�Ɋ����^y��S���N�ۚ�#T�pt���� ����� �!75*��	�W ��Z�ѧh��T�*�9�u��w.�w�S<6�N�0�̟	��"D��?���v��)�~�7�^]S��^����&&V���Z11���[Q8�#�����)�R,�����gI=p���#����EQ;R{�v��p�M�2x��N����ma�e,?�)@.��F�r���o+bP@��B����y�_Jc:��YG0l%�M�V���0��@��򒆠>9�����_��f�iX���kUHC&��Ѳ���sa�H�N���{N+��>\�j�������i�f�J��ԧ�%o�<���l�dJ��|T��<;I���S)�ot�9�D6�@dg�a�eJ�<U%�\YrdT�^��h1�"�6���Ln7�
��B��(�d鵭-6O�⏞�����ֱ������7�D��(����Dpm��ĂN��[��b��c�ñ��mG�(Z-��@<*�{!��z9+�%^��I5t��z�b_`�<¥�Q�J�Ԋ�������00���:�8Tr��>�J%�VЉ�����UrS�K�����ɕD�4}�v!�b7/+�Z�	4����6�'jvw��!vW�>�PC��ա���kɣ����y��3$�)h�|��	��\�(��1���M��~w(6\�'WY0-�[�΅]���4�)|¿�7���ڒa��X]<��ȯ�!6Ͷ2���
��L������ �u;���rQ�~�f�bm��,|m�u�f���dx���P7?]���ki�-�J�>3�S�	A���~�SV�-h{��1��A�B�k`�����l��!���Q��rP�jC>,3��LA�&�31�(g�7�C�VvR��g�(���dY����'H��0�M�8�!}��:#