��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܫk�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A��#��Hb�а~�g����o�+5FL�cu�ȗ$��ƃdY=�7,�����	G7P!�P#�l,���1:6���=(�Kza��@�F�U[Alb�6����M�����nU��ݔO�t����M�Ȍ'%ͪ�����qrLx���|n�`�c3�A���;�l�Ol(93��f�w&bA�x�`�T k���e�*5�����{׎%p.�$6$����ݡV�>���\�Z���:�?����� ���֒w�T	J-�<}�NI.	��^Ǆ�f^� ]xkWd�7��Ԇ�J2�C��ܧ{v:��|�rM@�eD����p�W��f�*j;�����L���~�T���"V@��x��<"c5@)����W��C�ۀ!H6�5@��,̂u�`����D=k�����J#�w�"�6�?����g��� O#�H++�S2y�-��i6��y�{���S6
jAR�4K��4>�h��ʓi�����\�iY^i�}7�=�Q`��ֳ���|¡��7xب/.��	��cl4a�D�y9kn��{GZ�F���wX����	=@͡0�ui�Orػ�*�^��D�S��dgm�	H9�r��U1붻��JtqI,z���녙���x���m����ɹy+�� yRl[�u���"��2���2�"⒩&�Tn_RKv߇6� �� "�e^�͵�w���DJ�M%0PQ���\AL��K�aEM�TTp���l!�9b�A�k�p`6�i%�*��3���8J��o���&�.�P�J���gGE��q9�&��
��V6_����(��̷I#�o�-�H��;��4����C��\W9��4�*m�x+$!�y��3\[�`�-��� X&���:ڬ��٘)��O�I{"�#��;uM�� ��B�Q���Ǝ�u z����=�0B� ���~��R�9:frIs��/z
�{�o�Sr���`~=~�L16w�.�o����i�$�p�eH����^�KF᪾%<�KC?�N��.a/�&f�����ʭ\��d��`����{�]��R�l:��+�P�>%$�?�g��RMa��Q6�����U�a�̫{{c�zj��)��Qq�=�N����13�9.7�SЪ�R�c����"$�:Zذ��PtZ�b>�!j���ܺ$S'�֘4�[��>&6��1-pd�1ġB"YlE�
AO&�Pݰؿ|�7T�������4<�=7W^��Op(�w�]�ǊeJY_����m�Q����������/?I�	v�s`�|'Ң�A�+�D��^�u��bU�Zb����6Ҡ��n\Uy��&v2�5�n�X����PFD�:�f"�1�bE���w�T�� ���2�{��q��/�����FT2���pf�0T�������+�T�o��6����n�����m�kҡ�"��T��sn׹E=/^�8X�&���x���Ց�1��A[�kV�2�.c���w�k��x�$8!E���Ⱥ'�t�����b�'l~�l��mC@��Á\��z���L�՜ͪ���*��ﮯl��]���\�0�F�$ᓢ��:�N�];'��Eq��h���4�4+���|�X9�d�⼐��𱗴���K�Kֺs6*��dJ����(��a�gT&��#��N&<{6ۀ��o�lE����w�>{p�\מ�j�X�[dvxtX��!�⨋C�SѭOИ�3��}��k9�6��H�]���'�F�%V� �����R��1��c�f*]��c8+��Y+����vYL9���C�y2�w�����Y�a-�e�y�B�>�"�L�f#x5���Ve8�}�X�h�RN�j�%�8��Ek���UB���Is}+9p"�a��Ĝ`���T�&��ȠMH_�L�2�6I��ŵ��,Iz��N�X5�*l�kY"�!�JͤÁ���7�����`:�����>�����*�3�]����2���#�-LAPJɂ2��n���%�*K���mǥ_��t[H��i�|����$��ȥ��1:���1{T���FP��z��GɔuO^:@9���� 돉����7�$��J]�^פP'�N���</��Q�m��")��~���/{���1[ }M�=7���l=����u52r�B��o��I�ڀ[\�gN4�톙������>�_��o�{���o�W<�n��-��Q������6|j��O����5U $1�j�F��5ܭD��3�H���+q�������p:�XR��g�7U���F���<��Q�����H�}�f�{cZ�؀4R��ו2.j3�+N�]&�P�\v$"3��8f�u�Y�<O���[�cP˰�����O�q:ZǞ�C�q��m�&ܶ�P�9�N! ��`?�/��4Op�-��� �yG{�K�"� $����/�����@g��l"��-Ƥ�_��}�`�C9��F�p����g#L�tփ�c�K�R�"Z�g�>B�5�W(���%���2t��=A�_$"L��'Y��+򎨑�����d�� �w�d�1:f�39u�V���PQ8��ݺ~�~C��J�Le����eԎ��Bl�n����@���l�3=�j�⸕���Ժ�1b��=�D�7ϙ��s��qj�AQ�61��:X�#����v}ؖ"
��C���=�;�~Ζ_(sl�bf3���?4����]�p�~�o�z��Z)3�.t����Z΍��O��WO!�� J��b�~�� rm�cAH�:J��]��p&������ `�4��(�m �>�5a�'�|s�9"���qL<dF_�2�/ر��wc}#�2��C0�Ũ�R�����z����w�X~N�o�4�ץ�k)��Hk坼�0T�g!p)ʚ#�E���֑��Q���0,�Q��a�*�W����o�tW)���}���)����撓����m��E#4]�)@U�sEn�]ף�#���Fb제"Ο�r�_�<Ñ���v�d�i@9��atj������ֲq
�y�V&�B��O�$��Y/��B��n���WN:AU{�P7
{��Z�e�n�־�
�K �%�ڴ�O�Ƞ�!�cc@���������UB��T܍�lY\�^Ma=2YE&�۱/`hNs��#ՠ�X4R�g�+.-Ȫ��b��#��s��o�KL�.�dT�B����W�������q�6WbBU*=���%�{nAAZ�H��(Y[0��Nu�$$�	���╡L�K����x"�_ ��]q��/��Z;ܕ$��֦���~�i�nɽ=B��_�2��-5i1�"L�w6���I=�r(n$�|� ����`�X仼��w0dA�2�`Ž�}�f|���M�x`�qz�q��,�����r�
����Ge��|�~V������u�h ,���:rҸ��E櫿
YKj�=3��Z9��Lōo�iĨ ����f�^��v:4��E=%��C�^�"���k������������bYj{���-��2T�2��h(�L��5�Z݅)\k��������f��]x`堮zL����ҁ�5����k~�kzlޚ#�J�Խ��۬t�
w�K���qo�)�P�'�>�;bVчE�\R�)��L6h^O��Z͓a�5ͮ�n\3v�9V���a%��w�1-g꒘tID;��G��f���ԝ��/>��� d��#��Q2�'$ý��1{W�L*��fn�MʣoJ��;��-��:�	�9yt�F60�᪈���&�rİ1�x�Z�"���)K	n�b�qY>�T�;�)�\<�Q}02� j���O?nQ��tH4��&(���U�0Ҟ��P���ٱ h\K/�܅����{�����g�,�Ԭ�a�2��?u�����}�%!:+L�{L���ԯ�  �$�7!�|En���%Ơ���Ncf���|.����p��<�?2e��0uv^�}��9NF�B��;I;]UzʄG�f�Cm1��h�m=(�@�G�;�Y#ڕ��z�sZsW������M���\;�zQ4��UtD?���w�$�����^�<��n� S���`�X��F�O#f&���e�_�C��Q�P�
 �
'�u@����|T��E�����7K�2���63��ْ���̥��K��dr��NIQml�q�)�itpn�8�#��cw���%i�S��fs�X��A u��+�MRY�o����Ŭ<��wǠ�ZJ!�+,QO�%I���_�4zvQ��eQ��װ���q�����?i��j!��4�,��jO-��՚�_���|d�u�*��y�b�{|D��I�׏�����y#&����V.�ϧ%�^�X����Vr^�!:����U�ۯI�>+o�boǜ����⍖T����T]��3^	"�a��%�������X�,��8_l�Ro��>��`�Сf��V�u����)��3��e �`�F�t5;^�Ԑ-=�K���O%h�j�%f)B���Ȏ�]���|,�XJ���ұ��?c��!�����+oĊ�Zbb��V�X}��r�[�맸��p���i�ϼ��?����9Ws�ʋl��ƻ��DW�SxF����!��DP�gD^���V�wՖN����=U��Z��hZ�MÉ��\��Z�7^[���ٺ�(��"��h,̲� ߨ��=h��'!�d;�ꍿB�Q�