��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�ϯq׆������s@���'����j����դ�P:�Cb�{�'�t�ɟ�>��(Hw-�u�� !i�^lZ��C�{��И���i�-|�|�I�Dd#����i��	�4�@$,d�������v=�3�A�pO�w�tE���M�ȼ{;��?4P:ٮ�7���F�ڦ� w0=L+=~�&P0q[��^�-\ߛw�T��e�z�"�[S��B=q��È��A7�D��]�!Tl�f�+K������<d��\�毙�����gpȷX[���;ފ@n�%%�WNr5��X�hqҶ�=PY�0��WΈ>��uX�+4 ʿ =�������5�i	��,�Hɴ���d��h�(P�pFtk_���'E.ݷ�T�q����l!�&˃S*��, �FȽ�'(�k���=J�?�>:̃�7�\���9����Px%[�C��a�d�%�}�qyh�!�ۍG��x�58��Θ�|l�zFSg�\j=)霃��f��L�U��!�@C(����U>�RRrT� ���X(�A�G���I?�/�I��"�?�Z��E�T�w>�3p�>����G�FJ`Eޑ^��&z9P4��,�N���*�
;�˰d~4�� ��'�L�͛�e��ث
|%��QLZ��s����9[S��ʝ��:W�7��������gG�^:�6���3=x;-��;
�
��_a���-�V�,+Z���N�69"|����a��tZ>�G�.�/�2�7]�Mg�S@~_m����7�ZҫӁ(�,�	2?���G\�^�����c,Sʴ� ���F�g�\OA6��-+���L�����**l�K��:H�\��B��r�A8��ѵ��1M jp��x���?S��p�k��ʷ8ώsr>!w�2�O���q'y,�g{"�b���ipD�L���#2d��!��K��VFha��_�
]{P���(���*8����N}��^�g���\j'|�
����S��D����ͭ��\|ȹ�s>��@�d.`�t3L���E�+�*?ҩ{*)�D݌����E;��Iy�bm�`����8^s�S�+Ϡj6e�A���T0h�p��v7�`��9�ʡ9N�E�Rh�\�s����$/F�ި�� kJ��M��?�,�&�+� r}M|��J���%��������$su{�C
Ŷ��vƲ�����g�"Zut�P�I
Þ5��������O����PMI�7��RL�c&G<Ɗ Ny��Q�H����X�Cxq��Ԕ %.��Q8�ӹ�c���z}���A�_�����=Ǆ��$k�'7N���3�K�^�yw�Y�?}�S�:Z[Q��&��������T��͇��*�䖈n���Ϊ����6=�P��r��>����,��a����BQ΢'�@zA����$h���ʔ�WJ+BƦ��c����)���t=�I�`1�O�=��t�]��������9��l	<�S�Ό��ڮ"t�͟[�ψ�5��n�nl뗤S,�H�o�ʼ�vxv���n���;���i�^Doae���-TK���6e����D
�:zN�[����2:/e�Vo8#FZѹ�	2����Z��Z��%����ޔD���{:"��F.��<L�L��)Lߢo��t_�F����g
�S�:}��!Z(N�/�C~��3g�������Y%�����9(� �D+��N�%9�a�1��'w:�gSI�޴��Ek���%[W��l�K�x���e���\kh����{1�~t�V�Y4�P�j3����$���C?	ʤ�� ި�a$�Y��I>�,���˷�6���;��R`�A�\�D�R����f�@�<eV�������|�&�t#�O�i���k�8�K�G!��)'�8��oT^\�m���=b�9�����i=�����7)�ڛ	v�z�魨f��6�B_B#K�3�σ�����62TZPS���������9
��l��; �H�a�܎ix���{��a�-7�6�J�H 艹�OX��ّ<1N6�6cJJ(�{ҭ5r<������)J�^�*lJ|�Ug�o�4�4�F}�� �G�`<e�L1	�V�N�����s�@�����Z��>�Ɋ^ɥ���1�s���[	r0,�Ihk���p�(w� �V��C>.^x���U ��*�H�S���Q>,��x
z]\�Z�%��=�{!9C���؏JD�t�-���gd^)�
C�ԇW⌆�Hgי�"-���<��5"I'���PQ�@�@~��NkJ�|�}=&�#�
���:�Y��;�g�xe%��k��g�c,o����|~M�x�]xi�w:5�!S��rW�S�\�:��^Շ�xf}�ϸXy�L�VV~|��[����lԝ,�\}UW�ĹR��N\��s?�T��sM0��`> ������0�ϒ�Qc�ps�� ^.����*��\���N����`��;*w2�*I��M���,!���l,�Y K�����y>��V·y&%���ȁ���#0���i�M'D&�V�N]5l��};��Ua�n��ǀҬ L�ao2������0�U�4�W1��J�jS廗;���v@���#W^���'���N�5�-�gS�;���6���r9�������\�g��wѮ�=,��4|��i�c=� ���Hů��PK
��`�ٕ=�]I��x"gr�#�U�%��I�o���:���&�E����k؞ޕ5��#@�������%�JU�!7��F�*"E�^�%�@@or�.w��94���&��x��ivQ����o+n��Zj�01m�P8d���h�2�7c��=ܸ�YL\��S�6��)�I�D���y?_�˘�(b��b='�d������4��8�?���[[؊�ֿ��cI�yp����Z�$�Y�@��K59�ҩ�
ճ~�N��_��' A�x���iP��p�?�#9@
��Ӧe
)���{0[T�)H��ՠ�����L�����j[:HKx��N�:<�(܌ՠo��*cR�t���$�
а>m����ŕ	x�:���7����@�Q�=S��ǂ W?>�9P�Y��a��4ʕU���~���nM�����@n�Dw�jS���zpJ��w��
\�����u���tC�Ŀ�@��΅�H��-[#@��_#�u�Ǟͮ�?�����u����o�/ՓZ�z�H�]E�ȅ��i�6����O9y!��1���;����j_��!1���t�}��/2��?nL�NC(SP& ���S��]�-�]k+z���})aX���C�!4��Υ�S	�*]٩v�T��F9��Ј��0�L��@��I�3���C\ޚ�<�v��zۭu����w�<�B��3�%u�5%φ���%�L�p�cAu�x��:��˖�ϝ��ylo8���ȵ"*���^��:������;��j�%���k�j���1��L'�C�x`���m�m���{�:��o3�a��a�Ic��W��Ɓz�u�ma�#�+��2}&e�k'\�یg=�'lۡ݉)o���K.�����R�Nn6e�Jf�J�3��-�S%
̬�)XL,����1���η���=�&��0������J�b��(�iP�B�-�f�T���Ț�[�A��9�_�˷ +����6|R%Ԋ$��>s�m�+�F�hMR�ޱS��C�9r�H̡B��+;G���:��׃.w�IlX��NN�� f~����2�k@�WT�nF(NN<J���^с�5�j��m�m�	��N��I� O�聕H���Q�U��(�Z�=T�ߠ�1I�v&�=�ؼ5� [n�q}(?�)	�{Թӌ�-�"Y�x1�ׂ�R{��t�������Z�?"�tp��w�%��ƛ���MbA?�w�n�&s����'�>��f���_	���6XA*���E�ӎ�l����g��G��d�M�}b��p�_�)���Fpt�	��1�24�H��d`Ԯ���P���H���&	�#�=�+���e#��6+H��]R�=���9Y�˚G#xs�Y+>�Fl��Վ��^�R�ߊ�s�w8��*�s���قv@�Xt-�������m� Ȧ/d�(�sy���q��IH��+0fYXE�)�?� E��Yo-�S���(��mjv�6����q�0�m/�;Qnb��n��'�0���l������}�D�./G��ъ*���._NQN�]y���R�絵sq����y����%p�����U�uD9��[N������In���$*�R͉3��?�`ɍ+��(���K��U7�1d��.�y�+���2�3��0��i7m*(E��[*+ŗ�7�����#�н���j/H�!'D��l1���������_R�Xݫ�$��o.+�_���Ĕ���0%+V����4�$4@���Z��ƅ�t=����3C[���mbGM�)���K�9S`����Buԑ����Q�Ǟ]���@A����6G���0�{���i�Iˈv+s���#����+����Qm����@�P��Ԅ�B��?��?�N������P�P����Jb����m���.� �#�����,����F+�r��y���H�T��%XYx9E����#)���6?9�9^i�g]�[��~�I�4ۖx&*)��s�~�5U�fT��κ��G�P���k��zڌV4�0�NOE���,C'��e�i��$��%T���=�Ƌ�_]U���:�})�2%�'�����6Nu����mq�fڶO໥}e}�i��\��
��֋q��B�7nǅ	��;�ԨB\��1�F��|�B�v7#AQM!�V�g
�I���n,�4*�U�a�9��E��:uw�B/�2�cϪ�?ɚ2Ո�/��wI���y<���r�Z��莶�#���ا!a����?!�B$��Ŗ���@�����5=,��b�Q-���s� p���*��N�1q�9��gFs�M��L�x��p�O)�gN���Iz[I����g��ޙs�X.�ܪch�!OH�>��b
����r��XBȖN����?V�)[�[�8�Ļ�YR��M��A[)�NoN�j
*���	/��5�&悺�+����'6j���ӌ0��Rľ�B��
�~Mk���k�9�s��ԟ����rHʟN�Z��/,HO.�X�Ԫ�	.��6;��$|��1���	/�ј �J�KU-B�eY�Y�"��ts�ך��7��<Ç�K����['W����֣��+���U|�+����S�kl{������!��g!IBp�	DSpM&K��y�q=zy�Ԁi������˚/l����(�c������.�m;�Ȗ���u
�7qLB�y�q����;J|P�{�GCY�N�3Y���\�1�߈o
�DV0��^]kdC�n�6~�Sela�7+�
�ڵ��}/bQB�l��C+�=;l���.G���v}��0ǋ�D��������.'�i����.:s$V�im]C1��%����~}�M)@j��p��ro�I�m��9�e&�@M�ū�]� )!������w�?��0�gh��Ư�x�:�}�[�5Q'dmi�m�rj�zP��i�t>}!ܹP�be�BY/�s?x��ٵ�{l��Vw�Cن�wC3��HG�z׃��$��5����qhP�c��5Z�Z'<D�Q8 Z�)�fe_�=��^���E����,9
a�<L�����'+.R1S(��?��RP�E4(	f\��&Oy	��h޺�B�Y���L)��e/wx�!Z��k��J������zD|M�{@�2;�ǃ�:7��"��j��Q�M�y
^��=����2�F$ �.���-4�y^�!�"NT���>丛����!�9 ds��{�%��7w3�4�#}ǈM@�%�Q�G��#��/��ǜ��8a5�2�[��#�o��#����T,����	`c�.�F�Q��RJ���\�����?˃��x	���'8�1o߈���ī!���v+�P&A�`@}q؜�q�F��2�EB�l6>�h���<(2ȱ�0}p�2��"+��.�+e+l������o�QN硙͒�d
)�zI �z�K�C����P��T��(�-N0��� z�� ���Xc�و��7�R��Y>;�I�P�6N�<=(�ӝ����_�_�z3��d�ݿC|M?y>&���T���?f�Z!F.����������3�zCK�,�܃	j��z�^��q��$�!��2�4��ț�>ԾY0��Y xXv�!C�Y��|o���'��Z&z��:2Z�3���/L�ਫ਼��UM$+31�N]T�=$���e���(�|l�.h�5���e�*~?Oj0�i`;[�z{�x9s��`�Td�.x[����S9�ƌ��3.rXҧ�2�����j�������H�k>�������H�?�E^͓H���
��d���A�wSd׾Fh�o��"��枸�,����w*q�h|�a���Q�Yl��PC��ز�[��I�Y���L�9�{�E�)Tu�\�󰒇?��E�l�<=l��tu�5�`X����oE�t��H�����㒗7{�Y=�#�S}�޸?u��+Z�����W{���ͼm��\�{�����? һ�S�X��U���Aܣab-�`2���=���Z� �(�P��ͲPV�-S�s�0�!�
���`nPT>Ly8:ʣ0��<r�N���h��}M>%�P<�q�Q��TVюss<l��B�<�ά���/�Be�� �Δf�h\+�6�T���A��2�s����g$>�Ye��Ϸ�3˱�"Gݧ��א�޶��g���K��7�į9�]��Zf��x���#��)^��'etS�k�=�ס9���+�����~p�d��vsw?+�I�)��jDc$���D�{��W1߆�M=�5�{��M ��Y�
�9��
�9�r$�:���QB��Z4�!�:��]0KLqf�*���m뭽�lZ�w��e�;��Ϭ��:�h<L>sSԵ0S��P��G*�s[((�����R�M�
�Fe�n�C'T����lC��90tqu)�|؎��B4&E��Ϲ��)�Y"��uZ��L�J�0�������!.~�1����ṎVS
@�e�O��\�ЖAm�H��'#�ՐIx��ю5ϡx�ĺ�nS�~f���Q +h��q\:�6l��Х<ޮ����!~%���p2X����.YՇ<w_��OÛM��|�x������.�K[��/j�%�(��ߒV�۬t����!���(��q#(J"��[�U��Ì_|l��k���?,���������A�/ɟ#���'�|>�|�k,��fG�Cms��c��^����z�8�yXf#�5�ԡ�>Z��5U:�T"�t8Z���߫(�;���]��)����Cm
���o����~>�}���{�ܧX��
��Ѧ�|�d+��l�����۔�Ԭj�.�Rܴ��F]s�'������d�cwqEb'���j� �yӥJD2�L���3Y��%g�d�/��/���<���ub�x��]󲴝h��+�L��f.c�>P]����b7��ט�c�U�]��ޑ;��Sd8Y���N�U�Zl����n)e����aO�-N�Ǭc4�W�L��
�p��G!ʑ��1��2�m,[�� �pb-_�hF�h/�]˥���6����;�Ik��Sa��)<�0��!�)k4�m��(^G�t�����(�RD͋wGV>��JD?`_� M��=A�燲�y*�vss�k�A�/v�-43��M[sz���g��}�@u�F�Ѿ��ZdH�ٜ~�w��{ۆ��"߉3���eMѥ�m�E���>�y>JX(S�G_��v����mhΑњ/�$�W$%PM-z�R03	��;�0��C�",��Q%���C��9�^^�b�k�7&�[�P�L�fK%�����P�[:�v�k1 ���OE�� ]�j�,��{�_��xs��Ek�,�oD8���fn�7�%�U�����~-T׽>^5p����^�ǂ���������b�k,5�mZ�����k�R��Mܷ����� �#�*I86�F��%5����͊MzW�.8�O��㍧�������kVX䪦���/�?X_����|OX3jP3`88؋gjC�%�N��g�dS�̔�EJ�!v�ʞ%�0�N�6��j?(�+���x�}%ќ. �<��h[�[�/X��՚EnR�7ev[�����G����\��"U�Ͼ��g	�I���ў7������oU*^�+�Gli������#|q���g�_�@�(9���I\j�f-�Nw�ȋ<m�NM���M
~�8��h?d�����-����%� �L� (
�W_;�-��8���<(w0��S겴��ms~Yj���ӳ"NTr\���!�j��E�����*��(�iJ�Vgj{i��:��%q���]��e�"tt~��<�t��y�]�{�����S�����F�R�g�JH�L�t��W�=�1?Yg���J�=#��l�٬HXe�G!!Y�I�?���9_�؀���x��Hww>,g�؈�).�	-�8\m@o����q3(k6giT�S�wl��Q���-B_��\D�t�+	�ҽb��j��c��eD�W@.g��g�Ȳ1�����$+�h\CW:�x�K�5x�kA�������r1��0����U���Fd��w{q{͎��_���i��k@��:5��h�88����=m��̭�"9g ���C��\^k�ߩU��ݕ=��G��T�N��C��?����f�ͬ놋��z u�����y������C+}x�8�-�i�3�����Yc%�E�.�昀%ՔLa��������}%����U��=9v�c�9;�z[DH[���yD�SN� �2q������x�ݯX���洁���H4Ũ���t9�g�L�����L����"/�(�O�Z�&��h��ӽ���L�9�����`6
��lRI"n���o��A��N��Bv���+4�>c0�:�o�C�^,��=I��I�n����������	�JK�(S��4(��P����#2��g��7��1 8 `:���ߋ-~^|��6��J�3a��\��x����@�S��d��d��Q�"!텊:/��q�h{�4݉�p.�}Hs��#GZ����x�p�O8�I�I/n��?Y�z�*J�^lT?�OomU�*��߷�K�C�}��՚�^Vq��S�g��H����:z��:�(h�۔�CF�z�w��?ٜݣ�U�@�� �/���FΙi" ko�b�I��h��B�u ��g�S,53a���r�*憸���x���BGV��7��y��PZ�R#`W������x�r�P^��($9ۢ�jD�K�Q�VVY4W��W�����Yp�G������&Ϧ��Z��b'-��$�g%��񼗩���=D��y����a�1��-���8�ύM��:A4g$5�ʡ�D��,�Bq��_�DN�����1~�?.*�m�����kZQ���vv�G7�b�4U���n�"��0^s�n���$ﶉ�����A�H?R4�S!���ʨc�vV��^]�ՔV�/zD�����}����:������v%��lӋmp�H��6ߠ���:�ۓq�TM���A�s"�[�٦��'*�rSXr���4e�Ă�[�`&E	3�x�4����8˸/��[<߿��C�Y�����f�����.�����c��4�yb���7#��~��+'W�N ��76,I1�nx��:4Fn�5_��)�Py�i� �	� ��z;8��ۈ��f�T$&l,��̼^��#��Wg������F�@����.�b��秧� �ՐL���5`�_�\B�AN\ϊ�ّ��8����ѵj0��G�	�d���L����bдӉ�D]V�y��	tL2@Bh09��P��HUe�ܡ*zay��c�
��{�-}��h�r�LZQ��X���HL��a��s�Z�����2F:	 1x"^'�z�R�~�"��vE,��'n{m9S��&Z�=cL/:��Q�&p��F�p���̃�	.����G͔m����!�?d*�j���JOK6�u�F��
1��R����w':��	7�S��Ӣʼ�(n-�w7Gn��^�Vg����lZ�'�	�_� �{����Q"�s�Aj����\N���b13Xj���[���45򐎓%