��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|e����M`p��E'VTEB��A)���7W�9_�ľA�}�����+A�iȘ+6�[���u��y�����9g���hə��:��e��oKBm�Q|��P��2�5\�xf��($�z�Y��L8&*
������ЦU��C���n����td�t]�Fc�����K]�\���M���jx��7^�V�\�)��5*��`�k��<N�&�Y��mJ��O�m?8����ÝA��������a��!`����?�0BYJ�I�_n�f��ǫG���%L�����j���rk�ѐ�Gݴ��������O�Ȃx
UV���;=
�8/�gX}�a/��dVP�̹wȭ�$�Xe�>��"�>�3��Pik]�������Ye��ö&�T�[������P0I{�X�2\� �����	��J�V�C��v�~^1yn��z�u�W_�
j���/͍������"�?7�p"�,�I��}��z�l^�a�g�N� �?(5�ۧҔ���WY�T[!�!��Wj»1��^mYȁ�������w,.ȓ���w��	�z[ף}��J��7�Z4efR��0�k����f��6^�4�O5���=@�I�$I�H��aD��Nin�)cZM�����<9_$��y&��QF�6��Id\[�'�q��&#�-\��f!r?�Q�A�$z�-M���z�m��]@]kc��k�ҽ=/��ccQ��D�Ŧb8MſP��r��+]���5NEZa�Lb[�R�H+'�9&%t3��0�z֚��&|Q�[N�U�����A��M��Ф����:�㾣	�S�v»b���F��N$��'Kj�?b��Đ��J��%閾��d��n
�9{��SW~)���$�`�cr-/�q	�a��7wf�̲J`t����i��}����jȯ��9�F��1�u�J5��q��Է���>���'�̢2�܉��=T����_n�f(d|�T���U��qi���z���b=�ó)���5�H��[-�h1Ir'�=a�_�z��p�B��"�_z����Ue�s�2��`����a�t9h���C\m^����Ā��9��4R��91��������ڣ��k�aPCЅ/���_WF�ń,����P�F����x���tNA�3�?rɋ�^ ��ך&4\�ŀ��q�'���1{k�qr����>qܢO�n_�	�Q��i�Nm�I��'����bg���g	�
O"�̗�j�����dr���`f��T�4y�nr�%֗� dj���	 X�hT&~��%t�Z<	�����ӫ���⽤귐��֑���ŞE���5�]U�\���1��Q$�c)��"��#;[}d�����|v� �et�`�~��V�y��E>"[s�.�[��_"Rv��&�,ؓU����.��m���@�4� ��"�1�wV��*B̧��b�gs`�WV��Hކ	R|ch��Ɲ	C���2�gV~5��WOq�x<�Ĝ����C�V�\Z2߲� .C�e��zy�7y����S���b��O^�۠�-�l�=77����g:9UZ�R�$6]Ht�]y��,�p��
 ��i�o.��;/QI0�zl��ޠ%��Z!(Mrғ<g�f�M'�5����ţ�a�4q����AF�eW��F�,��j�0bx�/.:��}��0?�+}�G'�%�5�p����wu9_׳WD<���	Z��Hwsě�(�u�����,�I����������2�՛�N�c}O��	�5��h�����ZR DdR�Pw;�Ԣ
������o��d=s�s�$���[b�_�9�u�K�Q!�EA<�Oo��a4d=}'���U��A.�Z��mWA�_D�9��}BW�����	�3cU}~&>4�|�k{�m�30��P�JU��K#���3��/aO���������X�=��v.��
�2߀Y��N�j�ǵzy�G5%��)�{�V&�ɷ�U�����[��}�������|Ї7&(���<5��W	5���� �����>��C7��7���9T`�b!���������uP�B`��l�@�l ��p�C�o1�E��>�] ����#G�~.oI[�4n'�Ru�^�����7���b��0�[���X��yx#'��'|����u?W��'Qݪ�A���U|ȸ���.L)#��ќhR�MO���Q��`X���*W����}����w[�`{����6��eC@��")#z`��W�U���
�/�0��]��X�ś-:� �a��?��%`����,B�G��0^�ǜ�(XLB�j?��e�����bf��A�~~���~�n2��s�q^��B�Nr���v��_�/*��?�R����έ�Pt~(�ߨ[�p(��窊<��@��"��@�CWT8h��cK�AC/���7tL���9n���]��@$��� ֫/�(��-h������C
��F�y�0S0I��}�����?�%\���L���},	����uO�� y�{[�Ñ��l�q��ՒУ��	��[W�/FBl���g[Ά����W#��bw��I6����n
{�V�M��B�D��uc�(f�y����A�i��m��3�
���E� ���#��&�$�ю��˼�nV��0~&=�0��h1ߙ(�w��U�k�l�١Uh����f\4q�Y���
X��2��%�t@�q@Li8dk����\j���0w�2![G��Sm�Ŋ���J*eN�	f-ش��Y��
�2�ZPs�A�B�M�h��m`��@l"R���� x�0b3���Y�Wj1EB�D����#QU�U�2w��L���`�%����$��.!�h}w�s��7�H�6'�9���gđ�S%P���凬NN�5�u�'B��}�Z
�4\2�zfw�ɐ���	K���'���	,q��`�f� �YA�f��Y�߳`9�����k��&[O���wwZ�5�ǽ������j,�_�� >f=�O�v#��1�ɏ�W#4��J�y�����ԕ���n$ D��"�r���5(I�e�)~v�*[J	�c�83#�>P�X~K�,rC�}F�����H�,=��q����JT)�y�ׯM8��vI���6�40��Lh.��,�/	�_[-7=|��&�yԑ�'[{�VkV��R���F��N�>���p���{7�����aQ���Nk&����m�X�(��Ef8���rZd�ʅ��~�8&!���LA��2�Kz�K��;�;��7�̀ƽZ�I�wQF)Vx+ ?����׋���xZ� ��ؾ�ZN&�.(����dz8=źe�+��J��U��6�@k ��8%&e�Da��*R� ��^G/���.���y}Ĭ��*����e���=�A��n�H�ȷPOAъ�� �U10:?���:ƹ�@,��%X��W3�2���$}�wNKx?V�m��<@^�K{���vf:�/�u5Ɩ޷�@��U�u k��@��p�U�f2��-6SI���.�tL���( �q`��c(fp���nQ=u�9d�f9�I�h݊Y���'�B��}�,��6�R�d�ڇI�	�^,L��7qw�+�:��L��Qd���9�_�����^�ү`tu��� � |T���5녾���Z����
͂��B��b�/5<Y�<~�v�_`���S���N���B|�z����ف%�TG�ގ����H囨�J]��0�)'�e�Gؖ$@���N��wP���"�b�Bw(W,j1h��	�An���wL��3xbeD����ZB��6��y�ڢ݊Mx��-�����y�0u����r����`���s��'��9N��bju�n����T�@.��௢¸ 1�R钰[���g��P���BP);�j�����Xz,�lPN��x|sjD�~x��0]�Z�L}�"M�x2����� sK��dU-n^�&�<8�x댓[TӨZ�fJ�@�A����+3oj	�.��'������֢�%��S�!��pǙ(Cjr��x���I2q���2�>�ԯ��YYQ�@U�:�g��ʭC����N���Ǹ���q�4b3��y���=�(�����4ܔ+_GY)����(��릋���k����2	c��*����B�w��-��,���
Ba��!��^^[@hk3e�*F�ō��hS��G��I��.�G[��>3|SxV���m�[���}���`mC��F㕪�Ӧ������r���a���<6�X�����9Y;r�VP(*�l\UKf���*�����0�9s�y��2T�'Aeo�z�#���.PZ��f�j�J�u�=֕b�����i�e�{:��g�
�ui@I�'ô�<�����`f.a9"rC�Ttv�TC({
)�x��|���U֣	/����T6<�7[�];D&�7K)7�폖�[�IfV�_ě����dC�U���w>ex�~\U}<�Z��B>��{�l�x�K�Ґ������o#$��yI]�C��ɮ5AN�d�uG���Il�ֵ�;�[��2\M�A�Z/��c3fK|5
[�q����\.EvE�y|;okXf�~BR���*��"˹��<��b�C���P	�y\�{τ�r�D�Wfac�ԥ�_m�q�sx��П�=�#�7D-�{-.�E��3yt)��P��4�����J��.�wp�R��s#�<A/!Н�*<���]��P0n1�Wb����T��q|� ���{����w�.�� ��4=��������a&��_)�Cc�Z����4|��r!���3&���:F�ɆC�P�*��(ًRF��q��	�~��r��bƚ�KƱ�u�{\��}��-yK�%��,{
�x��f���׊��������4-wr�F(�W��W�U����ޤ�g}8z�x{&�c��ef���5k~.�r���	֥i���X	>���n!�5��n��2P;�D���C�d�[|=v#�d�(�q}m(YE.2�.�z��rE} i��u�m̫��=3�U�=�����:�B�K��:�]��!Kf�9kk͍T�9SW�_o����R�����*Z�����x��39�R����W9�g=r�Q$7<_f(��RQ��7��E~`��M�.�%ć����+��io�LI�ܟp����:���qm%��<2��\m4���Q��l4��sj)�sATX3�$C�93�O|�e���~;O]X�O�x�>������� �b)�����ď�uJϷ�ʾ����(l}q^�+��G�qT����_�ഖ>eM+�d��Jf�Y��+<1c�18�������-��r���|��sI����f]�0�L�}$�:EFZ3կ�o�b�K������+A2���m����=B�����![��{|#�p}#��䍻��>d�B>�M5��#��J�n�	V��W(��)ߵ:��������X�	\�	�t�u�9��oL��2dB;`f~�:���6����&Ƅ���ՄU����˃�_�/>�[�RN�@1?^B���G|Hc�DQ�(i���B\����fF]Ҡ�Ĺי^.��IgI�ǎ!�:^�gy-���O�N��}^���6`;I������3���P�>f�A=܆4x�!=�:͖��J+Q1Ľ�&�j��:?~@�)��L�f����1��|ç����8Mk�$����4�[���<��3���(�S��4}|L�����^"�����|O���q��؛�fz�wM��6n%"=��)�($��>�Ы&�Xh`�ƺ=?G�);�zމ1�Z*ѝO@��e�"A>��\�D-��M)�J4^ƅ?wi.L�o��2wI�2��%�H�k,�>���o03��L�wO�� Hl'��^�	��;��ķӣ� �g=�H�톟j|��P@��G<������%���%"�쀸��.Y���?>���/}n+Ti��ZP:
���ت�^֐���J���jZ\�1	L�mu�a
�@UL��c�������5����� �
�(��Y�����:�E.Ʒ1G�h%�#0�X�4��B�)!���XrU0�w�2��d���]�8;r�({XC1n�ڱsj���Ot]j'M�zP��A'=z�B����۱���.���X4L%P���qϣ߁[Q�KYߪ�H�:�KA8��m������C�<�� ��>�^|���~v��d��d|�zK�jXa"C\ń�h�Rxt�.1�R�@����fODtb������8F����4��zv�X I0���S����}�B4z��ո����S�˧�G�c{d0�.*���K<��5P1��P�������j9"�Z�f��Mv#?����Y4v�� *�%S���t=1N}�U<��͢Q�wC6�
�C�K����a�����Ȫ��"�%Q����D��BY�M����E��9����1���pSZ��o^�-A�#vds;�*0���$���n��k�NI8'�O�0��ю�Qܟ=�_/U�� �a�u�_
��r�v���s�/^/!:�"�̓������V�4re6�3���������@�Gm?(������.���j���<��n�����1�h�Z%�!T�FD.�e����<�m��ISsW��Rsv�G�D����0��F�����݌�� ���Փ��[�Ô�}�3�_�'��+r	Q�a��'����� �j�#�J�S�P��G�<O����Wr=���������&��䖸i�-�$�1 t(�����'���}������u :�p��MzK�"�#�=�՝5������ y�3����ښ�V��ߨJ��6,�겸-��gzE��g�� {��2�|3�I���8v-=�	���ǉ�h�{*���ii��?ӆ��e���h�����8�,:�Urߪn��f+�� W��\g��qBT`�Ђ)z��vբQm['�X�.�ׯ��g��q�cC�����y�Jd�<i�R���C���`�HaF[����֞�Y�pˋFY�����+�,I�A��@��,G���CS��Y��(k��C�dA�l�8�����u�?˼+WC�?
g
�0S���N��<�)a�9`0NK�!i��)�+����͖X�ƀ���mB�6b�TH��|��{ʟ3�����<��2��[���Q���:��ZY���s���b^4B5Vk\�k���j.���wU�=Rt����M̥�/c�5�	�FB��8[��S	FCX��1�0����͇�-U�
 {�Ҙ��6<��x��'��:@���I����+)�P�p(�/�ծ}�U|d��\Z1p�f|�/�����y�Rn�����wX|���(�-�t7�Y����c��O��@G�H+����;��p�Pf7���(��Bq�*����Ӕ�ft`k��~�W�7�ԟ�_H��37��s}�lr���N�ǵ��o�M��|]��;O�I������>z�C��L͟�Vv�s��I�<�"C�M��m�I>0��3���,�N��*Y�ź>]2�K1B/q��L�D���*�Jn�F�	������&� Q�(
��%�7�	nDh�jp�.���.a]60��FRE�+��]6���|sz<r��'�Ū�ÂS�*3٩��kڭG��;���=�l��22�0O�>0�j��63�賮�雩$"���l�����P=)��`�>:�eIH��oN��P�sݺ���m�Lc������ ��A�Ȭ,-���UG�~0ɢ2sO�[D&{�<���ǝ4�N��t9�E�����������S�����c��z�u�30V:7cW<�I�4��EΎ/,l��I��IC-�l��p��9E6�g��B����[	�0|�h�����r���A���08�޻2y}�b��4���ܪ�*�@@U��.I71Kx�o$&W�h��D\U���H �=v��Zz6'E�I-���Z�Ҥ�`Ҟ]%����f����-}Dέ�}�Ƕ��@�`=�W����잌��n��3�	���Uh,�
������ �N-����
�p_�>y|&�5L����9�s�
+f�K"y�.1paD�B[/V�}D���D�Y��� 5��B�]�5�mC}
��쥐ֹG),+�+�[�3Fږ�ST�4Z�!�j!�s�j����{Q�c��)\^�;���s���j�d�m��� g���k�%6��wډdS�&0����|#���6�mJi��%�D��XXs�Hs�� sW u���V�n�N����CQes'0WnՁ!�z��U1�W{�Wm�Xk�)������*��"���YO�M��Zm��a�G���F�D�M��^���K�c�gG3S[ գ���oa2J����/{��xVl����0�Doz��ڵ�=<��u,����єcd[�0���Ȕp~��bkT�*�!:W���T������3j*��Y'm;�p�����
w$Bҧi����2�А��_u\%��s��.�!}���Vm	i��4�U�K��u�SGF��PE{�����W�y�(��R�La��k�����vN("����u}U���Τ	�d���@� 瘳���������I�����n�Od����ۋz�y��܆+w2nø�~�/l��C$ӎ�����\.˔����$Zf����7S��q��ފj[�Ls�M�.gŐ�Pt��i��PdՖ6��0OGg1�YoH�Vǚ���C����E��co��흒�jZs�@�����ӏ�O�@����y˂�����.	B���>��O܌�뮐T�*G̓�x���s�q0;���>N��B�d���m�6�Hk��P��m��Ҭ����X�ϰ=��~ͼ$<Ol��=�_:���,/t�(Y��+!�2�]1�.�;^����!��`V�>ԕ^���rܻ	��n9y�W�Ўk|�]�"��u�o�?Y24-���)\	���XRh|R���BQn�C���(FQ2m�y�X��"�q���DW���Y[2��^q�Z̱}ˏ��M2�n^�5�0u>
5��*>e��(a�Ē-�S\��u�,�<���ʙ�6��F~7��H��L䶌�o4bSu�U��Yl28���'�#��-�,$^<mh_&h/'SׁmlU3�Aq�35��V]�Є�r��[�qٌY�|��1���������^#�s�Uh%��#�I~^X3�Tz��6.{�鷞P����HD~�?��0�(��A�h���&�4,��F"������fUr� ��s��S~�&uy�D�Nĕ1ZD2n��������0=Z��VUWzq�,�mf���3���Ɵ�Z��<Q��27�h����f����&;{�B�%��]�I��O8��*^o=��~��9�>�(2C�(\rNn;���0��������|�(8Q�(J&d�;m���uBh{�o]��ۓ�Me��3/V<d�w�b˥|�K��N, �YZ�������:�wn�9�N'N��?Y]�!��Y��̈cb��"G�9���HP�����I+b�Γo���Eù�کu=�6��ڼX����`��:�LN�t�b	jF��'�TIQ���X������uV�=�KZ�̓�s���CB|�z)����;B{/��,��Pr�U��ۣ��-
u�̂�gx-r�%��)��WC��RN�M��^��o���:�@�K�w�_��Pq�����5 �j06�Ô!��*B�S7�(�l�����J8ٛ����t�w���9��@�V�Ѣ��"#s� �'І�:$G
Є]����K�V̜c�ν��b�ah6t�y��N�:���1T�v�C���+$�#?��,F�������L�0g/R=��Ě,��^�a�~Y�sDF4I:�� �ᴷ8���&||3���C-��:�a���������x����[��ba�\(�x��H)���Y�,;uD��M=@/��٧%�*^�3X�&�>�6R$Cg�_�S�l�~(�;��i9xZ���ԭ@�\��<��C�{���k�����NHä�Vqĸa��n���`�8�������Ȇp0�ps#��t�H�v�x���7��[�e,�*�>���B��w{U�k"+q��Qk�=�>č{��_�*���
��?�,ؒZ�n��Z��h���L��n�'���xY����9w����x�����:AӬ�����&�E,K�dN(��d2]�� ���΋��8��}�*�d�~VJH��r������DIID�A棙���H���7A��$��p{�#;�xr��0�x��l�dE�kN�d�P�gb��ݟan��~��e�G��WH������ 
�]���zC�1���X4�ӕ�[��յ�F���7GY�{>�sU��(Е��?�^��r�3sS7H
j� R8�I�g����L�q��sB�$sF������Q[�ְh%B��j4���HY�s�(�V������d� ��ҧ��t�n��I�͕�������I�@7�c�&�!�����R-�g�Z�2��k���*w�L�"ء�V``����@i*|�-AX�p��U֙���(jƲy5�<�׶��OՄmU�@�6;�\��D2�K�(N����a���+�Z��6+��>�yN�(f¬j�Z��cc��#IfS�S���<f�1 y@��Q�)+�Sۙ���τ�!/E.���Ӿ�ĉ���rhA[�4��:dY>	����.�9^����Q���D�P1
C���kK>�D��+� PUx$tu$������_�/��{@^���w�кJ
i��kW�te����;c{�b>g������@A!��R����}Z�w�<Ժ���G#�R�<�`���O,�����/�N(æ�Oa���m�^�>l��NUȤ>��u��M���6�܎�p:�+�6ci��}>��`U
�8Λ��]$<q�Q��.+0����R�����s>tw�� qO����k �_�rʶv	�L�tc��*p�蹷	�4cB��]��-ZɎU��6������@�G�`���P�D����E.�χ�����R^�k����#�̮�e0�&�Y��GZ��t��Y̷�o��O��?�c6T��l�<]瑖���H8���0��d��!�N�K�����mz���ک�����X;��I�>�4N�E8!e�	3k��
�P��*0�� &T��6�BM�;����Λ�R��,�"��3i3���T]��H��Tm��_���ѿ�s�}����{�r��Kj���������*���9 �s�)j�V-��I �}����e�z��\{������Zb��i�G}�ȕ�2BO2����ײ�,]⢳�&2���R�Ke�.�P'q���]B���M���߶��8.-��ї���3���wCj5�o�E'�sZ��as����ae�{j�UC���\!����i�$��*�� +�d6ԏ����f0�BO��i�}�H�EH����	CCg!|P3�~��x���ZU�ܙ��>l� D��5���T�d���a�%���J��Z�9o�AF�#����խX�^ %��!��M���:���Y:x�j#?{�)ey�GR-E�|���-̃U���^���3?� �x�W��N����av���O���v=S���7��M����T��(�+��C���<XM��#�ѡP"������'ݮ����{-�+��<��ثщ[�����G���i(��F���ˀ���۶Wd��a�aeM�r���B�	p��
�?�e6�����`!'�k}H�t�Xt�C�X�E��NB�W�:��V�u�>΁�&�$�|h�.18X�MW0�c�1��?�؄����*�_��00��r/�T�!n��*���q�7�'t�?��)^�6\*�#���}�P�yCV��6��I&����\�����0�X�� s��@�f��j@N�	"�)t|"�x�-�G�ɳ��'7�+u�8n	�k��*P���<�|���NmZ��i|f��L�'����>�OX3F��=��V+'?�LXge��[�u8�U��!N��ٿ�r-0sK�DH�Z�,b������;1�L_<���������X�.6�����8��z�ܙ��
d����1�E�vq��o0��Kn�2(�����V���ѫ�S֟�W.��/K�%���/l>�N�
�5$�O�� ��*DԿ��佸����/$ϔ~��M� �A��� T]���ъH.�󔮎���I!Zw
�՞�ȷ�4�pv���G�S8�)U�d,z9����|�G97�g5V
tMV�Tw^	�֙�0"y{� +Q߅��&H�6�����mo.�M�Z�4�.%��m!eNRws���c��J��iڜ��s�l��hU����0#,#D1R��pb誊f�s������,R�0��m��
΄CAK����h�<�2�c�"q5�8���lITq'�ʀ�|	3�}�7��ZR7t˂�\��w�����GB�g�ȝ�M��
�S��}K��q��zl^iw�E��j��C�k�M�@���p�P�و��)l
.�c��@C��5
�9;��z/�~� ex�Y���I�!��
RF>��R�W (w����宜x`K�a>�UI&���H�y"�h�K��[�Gj��$3[w��8�~|슧gQ�K��o:<�L�'����ݧALfB�n��=�ԟz��Ne��?I�=_�X��O����QY�Ic���I�8%����
�1��B<��{��9+��F�|��\*mC �����r�X�b���ơ��%i�Psa䋘"��@ڷrrz�u�X��K������4OA[aa?�t��R&��e+��p�����O��0�	��YП08�N�n�nC6
���#�UT��eo���(�F�QXI��F��Ԇ��x�+�
�y<�X)!��74����?)�T� �h�c<G�_��"�>�,����<��_h$�=���?�1F0��� �kb\ �U�]$w�'�GQo����$;�2���?o�&��y�6�z8��� �ʌ����VOy�ޒ�̻8SA¸��M���5���]->��oƾ5/�l��K�gM�t�?J@�ET�5F��74:{}�/�U�P� |, ^B�Y��fm�]�<j:o�6cM[��ʳ'"����s�h���R
h$?C��E�=L ��-ɳ��*1è�U��5���{r���ѧX��s�@�����Ǎ���(h�0|"~��zq��N�<�Q�f��$�_ٞ]{+�f؉M3��m5_�E>@�"���9(	�Y������`3W
k���������D=�MY�&A�c�}�l�������âx�����NX�h�2�+@�$<��{�bpJ�k�AdZ��e�i-*�QRv�H˔�ӷǤ���J�^����b�ʆ&��GMx�j$�[߸!�e�"�客'[�D��H(�H���)���m� �J��$d�-�hR����D8��6H����+�pzq������׶�y���vꨦ)E�E;<�IUJ4�:��_�{���%�����>�5m�0{����)<�NjN$!�B�Ʋ���{��ӌ'�˄���Hl)����Ԍ牏��3
��q(��i�զ�)�(G9��������W���c&�E{��"ԞV쩆����|��>�ao�d}n�u���fㅭ�xO�O��{����9!L���:�뛧\���W���Ŀ��-���$Wu�O���Dz6�s���d��O \����z9w� d�Bj|�v#�wiԌ�x�͵ΊS������r��M��T�^/O"��*\Ba]5�� R��(���ë�t|]k���!�a�K���#����p�nWB��V�.%���8t� mf��a���D�3�28�0���y�q8���p(*@�=!Lt�!4ne�	j��q�x#6D7|�/�Ȗ��\"�]@eG3..9�c���A�l�Mt�@�-[1� p��T�>���S[���6��e�v�7��&#\&�3���Fܨ�E�?�O%�p�&D���$�MZ����^�0�}���z>e2�g���pQ $^V�����|)����Onl��mR׽ ���ĕ��7�P�i�E���; ����F�?��~�֛:xL�	����(�^��r��
[�湨�����-������������P¬B�k&D�#��@}L�HEUh��xF�H7P��,�/Plg�$Ǭ�� i8H�����N�e`JK�T�ܘ8�_v��͞�P�����yQ_���cA�K-`�޾�_�唚�����K-�x���?N��sβi��^��X��V틻���އ����
�gH�GG)Qgwk��	qܲ�L��<Zcx��1�d�9��a�J�.h���n�D-���o$�����a�d��wͮ7�L��&*�8n����=u���*������g)������v��~.��ď�w6�e"�&�
l�)��ڙ&�����KG������3����%�&��B��L�{t���DZP�|B���b��A	kx/�>mcs+>o�uy�*�}����3"m�L�!Dj,�vE4u�	?R�Y.H�p�28�.8�|BF	J���?��8g.6b�j-P�w�lK7)A�?@
�T"5����l!a����na�/�>�j�e��T��|h��Z�E?B�,�銔 �s�W��1��$ut�ˈ���2���Ɲ��Pξ��n�3m�l��t�z�Α�m���y����6|�Sn��D�����AtK�`q��^_��`��+��I�ރ�$� b&�l��?+C�p�z׹<�L��� ���e����.������5�2,S�!�*�`����l��8�&��5�nB[�Ŋ}²��Ո�	��yʎ7�j�a��roƵƙmU�Soΐa��`��Dv5��`/�e_�yr��{�3�j�V�`�u,�����nL�W�w}�HU���EE0���+�ً���S�R�T�;6��E�fj�y�R���-���m���U��8�=,�R�a�ҿS��vR'�8����G�V�X2ʹ�z/	�}^���; &	�Ы�&2�ȁδ�~.�.yxc���
*x=O�� 3u8fR9r�[��`�8k�~/�k�\@ʢ<͔�W�C}�Y�J���ˤ��2�g�'���"��>�|cf�W���U���v>k��0��p�.��<<w��,b�rЎ�K���O?��	pK��$��r~���_z��]y�l����:���Յ�@=�ރ��@6OEs�L��%h��S<��÷\Į{
q���8./o�w�7B���*�!UЗQM�w*�C������kl�@0iq�YT_��S����ਠ�U��CCg5+Zs��v�C,�f�.��v8[��GLM�Y�B:���&?`�3V���T��ӈr|�φq5�)Y���dN�ڕ1"����Cn��q��3M��>w)��p�3�L��M��v�"�^�J�bv#�ע�u9ζb,z̹s�D�o����w]"zE-Y�]?�[��=�EM�faw�<��g8fL�މ��=}�-�{��Sp�茵>�����I�r>��u T���r�Q��k.5M�ݲ�<�D�Io�f�����$Ek�*��ɍ�hlg�6���)*�/2h �x�?���* n>������hc�c��J0\<��Ѫ�)!c���l�`b��*���h����t��J��~[�,�>�.)[0�����	�H���*�z��(�1�>�S�HZ?��H��V�ٞL9�D�L��xmD�&�j��ӏ�f�c�������k�!��P���ŀ@��/~_9�>^5s���3.�{
�=��7��z�%.�y-SR�Be�XD�P������SZ��⛕�y07h֮<���HA���$<YY�	 #�6�<~�6�o�E/�hu:X~hC��\2��X+T}XO����0�7ϑ�V����K�+�Rk�	P��IVzS�%�T��Q�j%��e-X|r4�]�K�b��-_�Q�XA`
Kr,��]>{4X�d�Q�^6[�O�=��|�-Q�B����]e�1��3?�x���"�nJ����چ'վ[�8&��b9��T'�d��������kI�^����v�#[�����
�w�*A0����a�ޜ��n�M	 yN����:9!�t5?Z(� �1���፱����[Mṁ�̈́�~?\���1d��#N��&Γ��l���U��� � �>��Y����vl�"�B9�����"�R�%}O����[���A��,�<�5�Q��uB���2!͟7�{�E�ًA($,
ZK��Vf�<&�$l�$h�tF3�#�����<j�N��T�⾮l��=�|�{@A��;Y�v��m�L�,��A�D}ۄ%��a�?v*���:�Q%�N��e���z$�B���g�uedYG�*�>O�F*COye��v��~+"3���'�ӣҳ��@��2�(~�!�le�&�m���Z%�ʓv;*M�ѽ�N�)���c4�,[(��0�;�p�%>I��<�C��t&Jm�4�`�~D��B1�X��0�N,/�Bw���B#�]TL�?���(�Ѫ<V5V-~$گ�����,��!�U����K��V�}����۾x��5�y���Ā���>�!*]�m9O��Y�4]Vǥj$�wb�n�y0W��%Y�*��v�����ãm��tº v�l@P �����Cܿ�%V[#��x��"�68�P!R�6��J�[��D�)(�х�	��@�\��������od�����������=չY��BS��i�)�p����T}��?�c|�=�G�)B�ؓ�
�l}��Ž*
)
H��Ꝛ>u�ds�W�ئ�b�D���R{ۃ�ʈ���@r��Vkg�A8�tI���L��K�}+%�`º.Ya���u�q��<e8|��6�m��y�z�qpJ��y��@�
���BY�xڿ����������m�m��fAc3��Pz�n}le���[���`�����S�/���Zj�81��T�u�p�Ny��b�5ů��i�N��30��Y����o��'��{��K.���jG�G��Vv,�d�+�P�#�ƥ��O�}9���Z�����q�3�7|蝰�!��6V<02�XiA��1�	�-�]�be��T���rW�5uEd7a.m��1}�%��h�>�#x��\R�P^��궈�z��OD �<`w�>po�j��G��oI#��k�s��-��`����`�ŬH�Jm����1�LT~��=N�.W^R?�c�m����#�F6�JBx���Jg+W�<���Y���TȘ��/F6����'7�$�"y���m0��o��JǞ��5��R1�;���*��l���}�A��l��:F�4�Ƹ�*�v-͙\������q���ja<�/M ��DH}��B+�YA�J�4�ǘ����{�t�H�j�����Y�r��n�t5bh/yگ�CEL�/o�"d��8�u3��7qمGd������!�df������æD}�(#;s��|�4!h����FɯJ��	���Y��	�BY��Q] ��(|�|�c�M?يk����9#+~�#ې�O3BU'%�tsN�ŝ��Z���qߵG�)��VJQ��&=s��L���(�����I�0催o�v�����8���F��[�Y����mPe#l7Q5{�-F#u�Xڋʹ?l�y���?�圣#�����23�����M���OÔ���-Ƚ2}�BEA�u��K�[�P� �/���M�"�"��fm˶����*��uw��߫X3�Tz���yǠ��ZkT	�#.
+�J-~����mE��e h�>w`�>����"&ڢ;�p�n�#���I%�ݧ��tNl�7�y ��J�R���'�ư��E��'o�\��P8Y�;+���I/����.#�π/���'�^3��ol����$�t�Q>�]��Hv_.�����&���Ƚ�9�bm-��/Èt��S��e�%�c�
�s��|
�:P�U,]��}�9��8�E[���|�N�p?���V���w	��ɛ����>����� �y��,��Tb��f+�vvPP�.��tR���	��43Gʩ�]�_>�f\���{?�a�H�Ot���♨�q��
gp�\��W������#&���8���z�J�eh
P�gI.ⴵ���!�Ke���J{2=�Qm���������00j�w"�3a����>#x�Sc���do��pc��!��BH������yBޥaga�0EW��c��`�y��#�$"���P��RXm��w���Z�-=78By̝������ۂ����V�ߝ�L^bXލ���6;
��7>��;�=�]��Ɖ�����l�Y8�RB��Xl��jQ�ha2�p%�������
ǣ=E��J'&6��uP�M�H�,j6x5�/���(Q���\a��a�!1�soL�ci/��v��[�
��EN�bL�
ęta��^�Rbm֤�u�CEM"��M�u�o�r�U����n
f$�&�Ã���4}B$ þ�P�"n�Alr��ޓ�zA�ո+7k�y�Fv�=��9��
�,V\[o'��ACwQ���8�?v|,�ձm�=�q�_�Gi�b&�ȅ�m"�d7�x��<��s�L����j�Q�� Wj�n� i����zX���H���Vc�M�F�qr��g�$��_3�0���O���(w|���[�����9"Y�58%��L���s�>ta�\[Y���W�6KP���d)ϡ���D�=��n�5�ը�o��������"y8�:`;ב7�~���x�?����!佇|� �!��8�=�!��O��h�X\!�
���;�B1�]y��ՕK!�_�7Ϲ�II-�B����[��:4/_*A��Z�����#�Lzm�1B�V=#���S��=;d�\\��z�24��"U;V��7�Eg�i��۪�xд�2��Su2ͳ��3k�m�˲�k�9�iǃt>~=�ϓP���2���'`W�G��A�&�Wqd�������ݵ��s)��@���X�K��E [�d%M�R�
��*AL__FAqܵ,�0�S��ptZ�xqd���9�2۷/�g����y�oLV�P�|NO:큑TJ/�=4�V�M��a�o4	����$f~�y@}�@z�{b���պ2�6=%�Fi��?��T�<��C�X�-��z ��Sj���-���d��7�WX�����٘ȋ�&͏�W�[:t�� ��`W��G�Ru���l� g�	��[P�w��/TmE��:�?�A5���}sT�-7��A&��b��A�E�ɍYal�a�h<s*5��p�-~(�5���2v>��Z��3�.�J��hv��uK��ϢeV,W��dI�Y�b��H�����#_���v�?@w���_�]��1T�̤��j�'�]�qw�믾�`���S4Gmb)}lafZ��"�J��<^��,���G�˿�8%��o*ZTuI������ ������=��m6;2JJ�֍��l(&�F����J{��9	=���<��Zˋ�^�kZ��� %1�pv�SQ�D��*MCp��$�������1_\9ڙ'�X�����H4)=q�e)[a��a�a�K6>�(;��4���9"��=Od�p��-�`uL�p�B1:'J�}[�D'�.+��/MW�~O+��d�n`0��d���e_0v.b�࿁�P���Z�be2��L�e�R�_-]����H�v�>]!�\6���(�w$`����-�v&�=έX*;��'�7@.𣏕@׵�����|oސ����٦��>�	��w��cMhf�uXHI��������B���ZX��_3�v�d�;d���7���t�f��l��pN-+��t���x�Yi����`	^���K^���{f-� �����a���̩�Οo\@V�����dy|5J�T&�͝[���k�	�B�����┬ܣ8����R�xY���s����t��ݐ�X��Ͼ`�7�G�D��I}�&ÊK���6ș��\�揼�d�B7Y����b-{c�nq�g��ǷD���4�Q��֒��n*|h�G[ Fl��;�~�"��Rj��.�>�H�0<�LD�����+���,꿵77�ճ�5�\ͭ3 ������h}���8�\o�����N�Tt�=���fUD�0+��������[�a�nGU�(~�ձϳ�%Z�.hsAtO,�0����]��Jk�@KEߗ�@�2%�
�3�����(>�M�1��HX*�	Fq;����ʹSO��#�l,!��UP��ar�q^Z?�G6O�ޥ�y� krNA����2V�x��G�t�~<Q��
� B�iL�������y�:m� �Y��I�X8�=1�T�W�'��h6�`R#~�D�k����Qa��ROR3,���8B�Q��<5\?�͓
���( ��Y1�X���e?� �Ѭ�+t���#��,�,=�<�H�\DX�bf����Vs(������
pn�"���8eʒ|"�U�K����� C�LH;9'�am����ƞ.`�w�Q�����d��FG��1�Æ_�rH��
WťJ6�5Q���R�-�q*�������JF���D�_�r[:����Gz��D��Y�I�g̒(��I]���=٨L�\D1�4���x�������9�8I��|�OR�Ю?m)�<#S�W�snD�!?�p�%dMH ޳���@�QB��ȗN������|U��S�p����Һ��0���w����uz�O�4��Q�}u�
��0�a��0�� �N�1e�vSx��x�_Y+�t�;�0�88��)�-Գ���-�����9���R�bb�ό8�X�(3�ba͂�5Iﾢ����&EtU?2����#�K�~����%��G��t��g�Ʃ!��\˛\�F��0 �I`!˽k�Ǡ���|�#!t햼D��u����%�[��{]_$���u+V�{\u��T�d-��_�?H�f�7�"��s�� ��L�I턭]xD��!�s=�:���ה�kԶ�@�}~j�E�f?۳�إ��~:���}j>^o'\���v�h��׼WM��*m�:����-�7�'��OE��d_�W�%�)�!�,��ՁW&bh9��(A���߈p7����S��������MW�Ui���N�c������ϝ�"L-��& Y/F��MK<��c���EJ�qo.&�5�i=po�g�Ȏ�<�5+�D.#tk^yZ�E��Aّ~u\��2�͎"����N//^x�3k�+O2��h�-�8���!ZO�{g;�c�8t�#�/EΙ�O��dz�W������ۨ)s�li�/VS�
��C�j+�L<��E7���:O��������<���0Ja�n�ݏ���������}�T��Pe>P��TDR&��R�9h��#|+1Y,�?H�l����\\��1�D�j���x)8��N���r2�=R��t�^�z�h�ǽ�i���)N�L(�	�8�2��MΌA��ՂL���cR>4݈�h�qi���h�o>k 9��uKI��Pv�4([�!+"���霨��	�E]@#�|��ڊ5��7lTTX{5э���%Y)�=�Lĸ� �Y}��Y�s�-p�5�"��#Ǔ��܇��_Y;�)���(��g}[_k0�9	�� �IK��u�4�r��]�����H�����n�MJ�$�\��	"�^����w�e:����w�@~t��������gmu���l_��:���;�7��
�#TE��p��Ƨ�8�wé�D�gȗ�3_��ES.Ggk`��K����9�
ϋ����U|�k/�/�D?^}J#�ZI��q���ol���d�ҸٳM�"*�}��V��|��;1Φ�;n��ede�6F�~�T�K�+�N���ۂ?U�'A���k#LW8m�OIA��M��i}��w�]g��,�M�-�T�\��u�#�uY��7��W�So���Sa�8E��(��Vޮ�����d�%�x�Yi��`�4����VY�[��Sg�A��`��d	�YcjA��1�5Q��͝�8�)�� 1��b���nA����v������yVÄ��i�Ewϵ�'��}ɲ��.c�m�K��Qt3i���)��*	���8�g�)$̷�P���6��t��߱%�����>�w߶��/rU�ȹ��� ���Eh��6N_5�EՐ1�@Ą'T�V�:�e��0]���1@x��n
���T��X��	��,dޱ�@
L�k7j�ڸ���)ё�W*�#��_-%���٢�.�Q��u�F�qq�~e���ߔ�׸-іĬ3�#���sC���*Л�m�O��$_<���K��ya��m �\x�R�_��ڠ8�u�����%?�[V��[tc5�����&�_呇�4
*^|�^f�����z7e�S;�9TT�4^	2�t�y�z �8�gHp�!y�D��=9�����m�d�H1i=��&�Aݺ�-�� }v%��B�����7<�ٍ�*�	�^~]�^��{��bI%2?~=v��߬C�$M�$e���Ϲ|Ձ�\��T�V|,2@gbC�9�L��'�֕�"%˔`�l�H�f�ݺ�4���q�L��>N�뜵��KJ�I�*'ie� �3Y����CC�r@	(ӣ 6w����+��c˟{��s�I����uK�FD55����E~�}��;�|.��^�h��s(p�e���މ���/�D�[˗�OD�����zq:��Y-��3�ÃI�ZU���Wd�5P�C�/"0^�J�^s.��jn=Ð��Є`[�tk��_��5�F�&���Ԭ�� ����k>�Hq%Q�w�D��o'��W�hs�A�I��N�A��t�v,�����,�y��ʺ(��y�	�v7ݍ[�A>��>���nvZ���ء=W�+��U�z�9?>[���,�?�wQ�b.@ː��ǳgyA���wA�'W\ߡ �״��C�	��ӣQ쎦���#т�ա55��� �YCM;_K�[���N�d���d`~0>�<�%��0<���'=��A�}�`"��^m6È���ȱ��v�PHR6R��_�wß��
�|���3�DZԇ��L�%��8�[�V��n�ĝ��z��[�EtQ`y��䁼��xP��k��va�x+F�8��{�_Ӄ��q��x+��jO�<����T�L��g�;�Ot����D_F��o{�6-z��-�r8XB��/�����$���vw��!����Bڠ���\a�#Ǉ�R�+�N�)y��Z{���$�qO�G�r�S]�o�O&st��Y�<��'!ヒI{g��OȃR�<b.�2D��XZo���kq�щRy�x���k�����4	�/r�51$���nX�s��"O�HB&T>f�aW�!@�2���.��W�ڕ1��2aVcV�Ӈ�"?`�Fd�sh4��=���1m\t1��O�E��n	��x��qE �S���W;5���ESU���w����XN몜tx������_;	-작��\���m<�Dh�7d�-�Q�E��
ε�}{��ue��j�l!� �E3<���ԋ���01W�V���{��H7J��ΥJ:��dn�W��~(�h��=�.p(H���u���k
��bA��Czp���?v�?LM_����i;׏�Z���ffy%"�6і�c�:��It����c�k�,Gr����T�Uq�se�qZ�M��߿��'�箪=�b�8I��I�p��E(�)�d8�a��
B�]�E�e�i: �3R��]h���z��CG)���jc�7#u9�ro5~R�'�XZ��&�P�|�� ��]I�x0�;�?��~����0��Kt��\��Ψ�;�����[	I��K`�)�..��by68�5M�kw�q�m�IV:�c��rIY�b'���i���U<����h�s���R}��I��Ԍw��������L��"�C�3A�-Dzuh��7ӋoL���j�硪����������d�9�I���IgvP�r��a(J�'uj������?ch�Ug�v��O6�s��@�/�=��x����'V�mdaLvx<�g8���.Ѻb�L�%���৐<Zt��觐ae��J�pŹF�nY5�#hC[qF�ᴧ�dʶq.:@qi5+�����ٍ��%J�1�������P-�2!�o0l8��2Ԧ{��<lZ�J�s���&��H޲�Άq�>�%ͨ��PA�U�V�<�;^F����ω�|%�9��Y��	ӾNWn���_����uo���#���W�q�����:���3u4��³qIe7�v#�,��r�M�e4 �4��%wYB�O�=�v[��:k�sN�&�#�Sf�)���0/�����o
:�``~�/:�����kw��8(M�g
��U;2�AeG��gJ+cr�Fa}u��D
��� �����3Q���l�ho��8�M��M�P�@"�5���:��� B�Vd��P���+���}���s���f!��h4#����X���1�����0c�x7}���oW�r|f�����,�C�6���%�8��U��U�Sᖒ����V�uݛ܎�y�N-O��o%�����g�h��+�yC$](��Y*��2D��ع�]Eت�kv	��[)߱�������~�'�*&��E�����۵|f~V���T���t��& �%�7� V��6>�\���&�6(��f^�Շ"d@���%�SN�	]��?�͒���O�A����m�~�'�F��z��G��~wжB���R���{�z��{ru`�q%�������[��y
�h�ƣ	\���G�4�{Z���8��$Ɠ*W �I�ea��L.{���e�Y�	���<�pK͡Q@S;Ȗe��jI�Q�B�ʎ�*�9�M���zi�9 {�;��o����͋هxo��g��}��:�q,�r����9�y�&6;sP^�a
>��\%O
�杊�-�[�~�ǘ�|t��)�G��1V�˩�F,���������c2�����Fs����� ��v�:Qv�t��o��{���Q^��㾒�=VC[�"����T��Z�E��3b����]��8u�DԴ�=qrD�9VsJ%��@>��i׍��R�6�S^p˄�-���uhY� 5��r�b>���#�d?�`��K��Q@�ot�ol��N�'�aU��9�\�-�N�gTVN{�C,����l����yRUb4Y�VL�%	���wo`r��i>mde0���j�~n���KX.����@��㓟}M�K�JS���r���/a7��,]���&����x�Ge}خo�К���k�Ed�k #��R^�J�jC�2�4Z���PJ���5��'�����Ė��򖂹g�-mht�8���$mA�غ{LD�?���w�D��GA�S��,��k�г���w��kN�v�m��u�PԈ��z�Q�w�R$:���b���ٕ�ט��F�7�7��/<&�G��~zH�sy��Uӵ�ܦ |�F����RpF�kSP�	�0A��kLM\	��	T� ���IPet�#�!S}���yGJ�ɾ՛��c�V*W626�r*(u��*e@��s��*<�yj|T���g��?���A��0O9u�!�(�

�����Q1�Ke���CZs��8����� ܃9���bǭ��9{zp��*2����_�&�^�m�<z�/���
\�M��So�N� 4�	�H�� \�l�H���FR޲�So}(\�����6W9)t\�+>�F���Ǭ�6M��_�*o���j���M�z�/!e�h9�5�d�z^��� �U�5�K޿pcoʉZL�KA�7h�.l�4잮������Jܿ���	�,i���@�]�9F�`�8�k7xi��k��Qa7��4���vB꣈B�֮�e4�;��0���^�Qmާ�<�����