��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��nͳ�R[�ظ�_����Qq���G�]~��\�^�W.Z��ke��X�?�I\�zA@���Y"���a`MBl��$���X���/~%�cg��OU#,��;o�w�F�~�wy�0�Sa��qC�$�_됲��ݗ� ���D��.����v��C��k���<�$J��3��I
����<[�P�}&ʁ_m3�P{�
A���-X'�H4Eml�}-���i���[�f�c�:p�D��oC�b��ˊ\�b��~.���������m4�G9cJz�@��&��q���:���ѹ�Nnk+����iq�ڥ�%ca_�P�e%���b��d�C�yi���&�ܧ�A�r�}~X�du
�e��sg�gF����x�o���Χ�xf��U�'^�b���S��	%�u�������Tj2"]�'4�ևA�q�cw4�#��Z���g�UAKF����zq%�d�߮�E�e�M��B������	^��"}�������%תddu�6x:tk[�	C�X���@�#�9�g�0^KZ/:٩��%�&S�$��V	r�M�Ԝq1�ڒ���7������n��T��g�N��]�A���d�r`�+�`i��%�Q�逊A>M�â�h-lf�.j��d�gm�W��v����%z�C���HuC�;��8 7^��v��a	�����KlK&f�	HkNN��Q%d� �P��3�vY}IA���^����6[N<s��t���b�Gύ�V�9�q��GhQ�j'`��/�G@�^j��i��=ì5�eC��/�뉢<$���R� kE�1��C(�O��!�`f�2�WD��\����<�p�bl�p�	9��W��č�h76p���%�Y�m�S�u:d��qŬ�w���##(���n�uO���? N�����d;��QJp)
sT���1���
3#��J�q���Ƹ�<�"���I[�<[�ENk`&3&�mL���b6/�o��\܇vi6Ezگ'".˜��W5��K�h,w��W�����Tr�^!�}�׀ȓ�i�ا&���=������)۾���4?��ª}OÆ���ږN�}/��˶��K4M?�F�r�-\��jY:�����J"��gy�c)i�����_-�ݹ90nT�B���u��1L���ۭ	��
	C3�EJ��x���.2���W�~��GW>�FN)r�,�(@ �V����
e7.DK�KA! �$I\;�x#M��͞.�=i�C���ω ��|�ƨuJK:�ɯ�_Q�^�4�|~��Z�s��8v3�`T���@���n��EF��U$2,�5�������E� ]����.k�y���FPZ>%�'v,!RpgE��7|Pqbj��x�mF��}SU���5r�OB8�PQ-�|E�J��Qdy�ظ����EM�TZ�1$��'y��}��j?�����=G>��ZT�iȨ�,�n�j F&�����Ü&�fRhU<�j9���MbA������Љ��0_����#de��� ����Ta��o��a�#�#M� 	�a<��3��Q5�8� ��܇��CoA6ic�n#�[Y�/�Xr'q@_�m'Z�y����6��R��R�[s2�`׏��=p�I��Q2 -!GB���߆��o1L��D?��8����i7w@�G�yOR��45�+������V��e>�>A�����q᷌���%������R�Y��4tt2� ��۷����Oɵ5�����m�A�#*)��/dEX�I��������"��q?�	����u �4��p���8�nk\L#�C��[�J�*v�������V��0NK�q]��c���~���K�a��%�������);H��8����᷷I��q^ӕ�w"k:Hz1	�9J����{d������@c��i��Ջ^k#�3j-%E��Ӹհ]�%�w�� "h2��G�@�WK ���%��Zc�ȽU��]^z>˲%�¢�=B|��\�el���^�PS��`�A�o��*i���7���d�:o\z��Y��_'R��YX3c%�H:��N7�Q�]-��n*oi��٪�>k��+r���r�� �y�^b�l+1c�g�ѳOQʋ�Г%�4��u���;@��p2Š�97���d�g)�N��vntH�e�X ~^�X"P�y��w��Qٮ���=��ֽ��	����Iy0P�m�{R՜�����Ǒ|�hO;��A�)� ���l �n���.�Tt�p��a����sN"�B�st�*�Ɏ���$��G��5�ɒ�S��#,��:@���S,�̏�\~{��Y�4sv�k��^��5�?x>�F�(�.=EՈ_q�#&ÿX��.�.�=Ǧ���� i�ҙ��!�� -H��@�DR���|��Z�|�/L ��6	�\ۚ��K�@�2�u��h<� �����j��P�w��b�"�ݾ��K�TN��SGXS�n��J��_Y$J�"�����ܬk������(��`@d������uj��Y���a����,lj�����d��hW�֥%�)��b�ڲЕZ����c�R�ߛ�I��w�CvP��;���d�0>(Ď��giC��Tؐb�Ŕ��^ޞd�����T?z�T9O����
g~��X~$��Q�8�7�u����kBj��п�-F��7��i��<�EQ�j��~OS ���~7s���t�]���v7}׌Vvq~Fm�%�n�~���-b��|����6�F
V�&y��5�/#;|Ɣ�������K���7�q 8�ܠ��!�/Z�b��R�՞�Õ�naZE�&5,��tK���Z֍��.�shⰜ��ݣ�َ��G�+'�������\h*��f���Up�5O������5�"���h�/nE����W��y%d�#�5M�t�rr��<˝CН���&/W�����7n9QT猏=FH���6�Nd.���U3��ueuæ�{�}6�Dʅ�9
�/�.�.ߪ����*�_�o�lhSl�S�y�A�isg]���T?R�w*�~NgH��c �˺Ķ*�&'~�&��`��ί�/
�Ky��й�7��*�]�s�ag[�3�dt�Χ��i$A5T��F�U��5�n���a��d�u��P
Ú�aT��3�[;l�޶5�&�j i��7�U�eL�@Ò������.�#A�m�#	�Vy>C���Ɲ�w��$����#$0�H�sLК�B�=id�CJҎm˴�X!C�<LB�n!|>�>sȼ�pr�8�����Wʇ"7�i���c�Ξ���p���9r<�r|�w9���&H?�ܰ�R�?�T�)��Q=�a�g�{��lዟ#qA����NC��|�0?P���T�M��ڻteA� ��!�O�t�D��)U�3MNp�#�1��T�ś.ղ{�.��3�`�'P.ۏ,_:fu΃z��#�R�PFC��7A�SLAs ���{�t]	Cv(���7l��9v��&05r" �pӊ��g5�M7I�QT+� �����P�g���� ��j�hr�c��W{(���H���{����XoggNn���A�Ԝ�p} ��D��>�������	I-�z���B���c�g�~o&�C�@z%@N�\�B/����/pdj��L������I���B���"*x�#�����4��2گbf,Z������LƒF!��rx�x����>[��������H��C���\��1�Z��w���C<��xڎ_�n6�ʔ ����]��8$�ۀ�A���kk	lik� 	e)P9O�1���6��k�x��b]�>���p�S�K����0�u��"A�c�Um��P 6,f*͙SBS݌����/�f;��<��$)�֝G����zw�z�ƕ����C�2͗���"�M��ka��a��Bϥ ��E�'ti�9�2,�����B&~�˔#�e'/��s�##[0׶=�����	an�l�j�9L-ZTFpk�	:���""o����;a﹇eL���[�Z$RYO����V`�9���׍%�[D�{��Q��N���H�]����7�x��Ӎ��,X��~D�+7�O2`|EK�L�=���O@ۏ���,�y��f�N����s��&�'�!����נb'� ���%B�sb	�?q5� �@�>#��q�_� �Ԓ|΋��#e!QV�vk��˗V��ܙ��d���;��e��Ћݕ�%��%Li��v1F��~�3t�M<Yn<���j<1�s�