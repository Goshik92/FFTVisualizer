��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��X�O��v��y� ���=%;��(�Ͼ�����6{�R� �5�!�L�q%u��r���K�����u�/��9.���c�Ӵ1�:�!�_\�P ������ep͊�Dɭ�}��U\��|1�[
������	.B��8��&[�$�)ֻ!Wۋ�Xq7�1Ƥ��+b��@a�Gѧp�s9��"K{��'+q�H�����*������\vi�?s�2������$G�A����n-���$�N`(9I���Ty��)��-��Ə�U���Ñ��^s�m+E.f��S�{���I{���=���u.ٱ5u�P�8�(��$�V�����`��<�eI�_��W0��\YN$*E�i�w�|0� w�5H�������־ O�/9ܸ�|�s����#�?�����QÆ,E�oW�a�җEt_bؖO�*^s���W�tN��_�}��s��M<o8�p/۞k��Cy��l6�6j���K&��q�\���ܮ"aW?��Sf2|�\�"�wT͕��^�w�xI�e����'^α����=�����%�OC�������a��GwE�~	��Lt���R:�q܆�v	�b�`l<��?�f2pf^K��^j�#;�S9obջ�+����&P5p�j�T�'�Lؔ!��z��c�]��cS���Z�e҉�G�K�8�e��]�_Xd�o*t4������-�~,jHY$����.9�c�<��@���G�`��c�:�5{�t��IAun?uO��_�|UvU�Ei��(!hjg��-99�
~�����,<'5� �t�Ѣ�d9��g(����A�Y�f��qL���^��S��sY�p1�n�K>���N��X_�!H�G]O����,ҫ���b�(M�6*�:������+�"�����gO���-���ʕ
��/K��(����S�A?�L��������=�;�~�|%�t	\6��܍:m�����:�}e␄� �"�C0]��Rt��fX��R��"����a1ɳlE��z�p�߃=Ϣ`�
����HCɣ����	�A��Q��Ϧa��Q�A���[�Fje55�.�^�X!H�WRڬ�A�����ףZ��.dD��r�:i#���N$Ph>�)�����tv�&���C�;��(�sI7��}%��m� �JzN�<��l�<��3,�i�Kl����"�P����*�6�rc{�l�� }��J.���ܜ�O���x�=$��Ls�6��*�)�"��[��/�]��'�>�^�&�N��J~����W�:�������^ʔg�Nx=�w}5�JN	/���A��@��i�`짗�.ߍ-/��W�����<�$��C[��Z�qU�(>lS�ы�e�j���xz��E�眢�H)��!�*BZ��{�,x��]C��L�P�CVM�Xp:���+:L��[��D;ڒzD��zW�!]��Yp�)�8�n�>%��v씞������j��7���	]Z-��'`���b�sS4��\��߃�g���5d���l�^�����S�k�ڪ |o ^P�pG[�q��؛��v�mAU�Nǭ��JE�p�Jq?�HZ˗�_ W�J	�G�k���Nԝ�7�8�ޔ��҇��Kqh�0�8V�l��|v�����s9'�)q&�V���w�A��W7]o��{�(��o �co�B�e<8���"��N�'�c5#�qf�~`|7N�H�V�T�Ui�2&I���x�2�Z bk��iXIQ�	�A�%�pJ1g�CQ�^�g|�Sl��k{@x��żދY5�P,�M�~1�I�� ��%*�ir�:�g��v��+�e`�O��m�D?��*��P��$;f��b�'�Ћ�Oe4${���iٌ�������\4���n��vA�A����];���Ջ��C�&w�k�|<^V�8~�M���[u�eI�>���x<	e�T�C�����a�[���cw9O|��M��,���EXw�I�x�z2`����}�}P�����hQ6���������܆'�+m�����AȖ�6��>�I������ �#��)?��f��~���`��k/�;���dh�-j�J�"��8��xI�M��I���*t�7~&V�ej�Z�NqKýM�~�[-��ɠ<.)3�=t���M:˷ʔ��j�)����Ž���:D��G&��U��Ǎ�(61v.���*SS��Kw��&u��)O{��u;��W�a"1�ܙ�m�/iV�/m�K?ف�^B�)b5]4�)#W�rwŗ��S� �-���]���B��L0$��5L� ���-�f�ٯGv�����
�9�De!ږ�������6����M�O�h:U�O���փx�?U0%��(FZ�M�{�>�ܵ�H,���;ڇj*�=B�>#����Ze�I�*x�$畳b���ڔp���%�����	"@d 8+#�{�E�q�*SA(ζ�1�ǆ����%�ݠr�.w<��:�!�
.3�qJ�ǦI_]>x�x��6Y�O� 8 �*Ⲫ�6v<*����2j���hƴ�y]�֫��"�Ȍ�>��i��6���p��AR�g`�e����Cb� C;��Ѩ���Kk��{P��J]�؅E�z�������^*EE��>�0����3#�q֟r�q0��C�����xU�u�R��?0;����PS�~|�r]-�䤋;�WL��Q���2J�D������"���z�{&{%"o�[��ް.����h����+�:�I3�kt�=&ڌ9�G	U��<�����S��'D��{Uĩ	y����k�� �8R�ݤ����y����wұ���q?j�BI�E��%���Bdb 8�ٰ��^%4L8"g���Թz�w�&�5LfM[U��2����,@G~����u��8���%�T�/�&�̱���g{�� F�]U�(R��V�ys,R�k���h]U�|�E㢬�o?/d��y�c0��P�!ϙ����?V�c���G�J��l;�ݔuX�����ϥ���,�>�Ӏl;��zb�ӄ�fάɖH�����mQν�|?���-��Tb�K� ��UbO+��� ����.+�̳G=m8��ꖭ,���~��k�dg�o�P�f��`7ox�{`09`�V�7��|��[� p��ljx��AإODWT�u?-����o�hfTV ����ޑ����:$E�O;��,,���
��v!9��� p���I�9�n��L�-�|�wv�͙ȭq����zf���F�>u/�A�� UgZ�c���u�-"�<����+� �r!-���F��-�I���D���y2B�5t�_�v�'X ���o:�¹�����"f��mǄN�f��� ���Y=�d�$����Z�Y�?��1�N���_���k|c�k�_o3��&�v�����Ll.H�g�Jē&��˺��
�ū��綉L���Hs-�.L[����7�;[.��9���:Ǆ�V^4&P����p���k��
d�r1�M8+��ዐ"�n�σ�>�iI��,]s�>�]C����!��͝�f,�?�x�i<:l��q�-C)�U� Q��:@�J� Fg%W�l�L � �)ߕ�,kv덁R�'�����n��.!��ɩ�LC�!��*��g�7��N��$���|�y5^��C�7��ԕ��`D�P��g5��/����K�[�{ؐ���3��y�1NQ�X��9�،5�6�h���~�cԸ��r�q�8��a��gz� V��2�~~�mm�20��mpƹo���&Ox�_0��A@��446v�U�	�6�[	��?���M'�0X���B{���x����"��>u��a��H�P B6⨥`ɾ_S�8�ȕ��ΐ��O~��ы�PWzi��"߸�����j�pk������#M���?8����O�arxu��}�����6mM#O�����8I�Y�UT�pg���{m�_�=p��2*g6v��RR���J�|t.ʏ��~p�8Jc̓���v.��f�����?����|�?���!�I�T�v��>��c,�&��H�=�If�;�<�yX�G�S[o�gm��k��`�[��h�4%���,�r��}��<�눏`�h^��W|��g`gs*����{�ǔu�0�Rv�?�]8���À(&�d#\S9�qa=
?8��L8O@ʩDY����r'?�aa���(�^k�:y��T;|�c�UԖ��J���oV���
��Lv��b���>_�,~���U:�w�\!�-����F>�z.�m�lÍ�EN�bh�X�^�~nQ�z���0�t�{*�Jt�Pu����b ��}��D\_����pD�R�uo��ݿ��c��g	���_�q5	T`6�.�R���R7ꈡ��@y^N�뉆!�T9հN��������Up5���*�� }SM�/I� a��F�V�&���W��=�2Q�� ����J�[��{�e1�;��%��zZ�KG�6��qY��Ռi�M�|���m����R�DKGH���̴`ҕp�$[!�5�]0��L�z���0�Vl��&՟�e�7m�g[!<�P5*�]fm�d��ϗ�ZD� >w�����cUab���a����H\˓N��v<sL_�m[;gA���a ���Ǹ�ˌ|����E�\���x�/wO1x� �R1t?�$v����i��l�(6r_�
OxyUfZ�������`LנT�����Հc<"FFA�����
?_8TX9�Wu����f�(��K�Dp�&���kL�&b<8�W# U)|�=k��@������P�]�~���S}I���1�7�(�_�\����M�7i�w��EG���!s�N��m�w]�Y�}�洹1+��u��O|����*Yj�I�;��d��'I���z5��WmZ�΁����ғ�t��A�~�m��:�������^�!
��-��֒%w�u���q@���b��[��SB���1ϱ8�i�Q���ÙXi��M��0	���:���]h5f
U��u���(�^QWg|�-Ԫ��C4`�Ao�x��EBE�mH[�h5P�S�#�����P�Sǽ���8VC*�f���Iyƾ�_5=�I(�՞y����ֻ���y�0��ԥn�����@�]AoZ��j �$lӠ9�����-q�k�^ׄL�[�5�tU?{.��X��>bt���QS�fq5�%f��}c4�[}�?K�yO=�%a�AR���C��
�4y�����b(I�!�\��>�~Ǉ�?���8y��Zp
���7uc=��I����#C"�֟%���$�N�KRN&1���7�^�-Ϸj8��-I���>�އw�.ޏ,�樵3��(��}蟴�>��[)�QX��Rr ��hvep�������IJ�.���1�z�)G 	q���<�ƾ�@(ڤ�A�TM�E|��7M6>��G6�>��9�����b��J'�6���ނ�q�	�#�brP�xiv�cJ);W��j�tf���7ӷ�w#]�ab��L�0��Gk�i�~�w���΍���	P0o`��Հ��i�,�5�؄�]����<w�b��r���@D��ͬ�m�$�$��g��g��ڞ�JN��%'&G�Ѐ߸�[A%�D��[?��y]��ϖ���=���FPc�ۧ���!�J�g�$a����'��Nw��z���kIND��ӝX��k�4��tc����I�Q�{\i�^c3���0�.6����-�)ܧ8��
�j8��Gv6?y��
W�y澛q��9�C���4�;ZU����/�ek��;��/f/��c�S,T�7ǖ^a')�ԑ�`͢��eJݕfv�4���O+�᱆J�ro�|�#��3�;d�d�cC4I����T�"�i���Y���{D�����30N"��f�ǻi���O:�D���~*���{������ݱ�)�V��N��@���wQ)g�#�ozA�ޤ �߽���4�fw͊�ø�Y"�E(ե}�7�5���-^���P