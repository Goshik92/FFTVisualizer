��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8SjfSު�U���K��)`�c����P�k����C����׻�U�(`�-�B��H�0C���)Ck�i�ο>mY���w@�^���G_�_gJ�t��$�\g�L��Һ��st��J�R=Ϻǅ��S�5��E�2(�T�!�����;��
f��W�(�G*۪b�r��ٻ�� �dc}�f���ue?��=��4&d�Ѕ���� ��C�f)�Z ]<���ڰ@��%��j�(�"g��U����n�E�d[�+�;���g�L��6G`.Sń�mZ�S +l�a��b�z�u7����q,���7j��]����Syx#�E��h��x`Y�����/��r[4;�ϝ���/ԫQs/&���f� [�G�W��=/RJ�B�0�9l�$z9�Zn�;6����{Imu��EZ���l�/�Vׁ�(��������MX*zk����e)����zZ��Ψ@���Fw�]�|��c_�i�ϛqği��,�O|��������oV����%3�$���I�-��"�ג�Jc�xb���Z�CS�x�r��u�ۜ�-P��S�Fv��6�.�v��
����j)n� �g��;��x�Ӭ�˕�\�Y�4�#�i�f!1��vd#7���n���oh�_�����NT�^���=3�k�#�Ќ���X}�gܻ��+�)���̸v$lK:*��o��g�T\㳲O�⹋ �Ï"�1}R��#.���Fh�0�6<�c0��1ޫ>fTŁE�MR�1�VO��f_J}X�6 ��6FI�V��C��e��O'�6�T_��n
��m���<m���ǘ������`l23��g�'��\����fʍ.��"~4�h��v_	n�k�	n�
EL��WO3�|&���a�����Q�5ԇ&����S�dԮS'{��[�'�ζ���U_��:�p�m�
/d���������Q��tA���^�9�>��h��S�����B����E�����d<��e����n�X{2�y��,�n�;"3�6Mi���X��ֈnn|�j\X�&��M(G�2'6�qE�t�W&���5A}�����~R5E�w>&��.�K
��d���|�?�_�x��"��cW��Lo^��f�� i�����?+�-�8�Q����E|�Q��<CF�S��PR����?�벵�؀Ć�o���?�t���W� �=�`��E�yF��1�0���d�V[1���a�|�a�6�=� ��BN�F�zؚ�fDt��L�g/&��P���҃]�5t�-�=��CM!>]����0t�:�:M�t�Tva���#ػ����`l��Р��!���+���C�ѿ��O�1��b7׃����O��ӂ�VӃ�o�?]!���c��v0�_p�����Q�,�}y�)n��r�U��;Jk��	~��TW�o��2�?n)�|Gr7�:�N���<|�[�E|#��?8����Xl���W�2�U��^��Wg�2��Gۚ~�9��!dg��Мm�5�p��@w|/��M�9���3���VU�F�e����4چȫ5�4b�W�"��`�wMO����w�=Va$c�6i����2l�$�~�G����L�ď�	m�BrA��UU7��w<�ںGC(0akg�ɨyF+�K*?G�tf-)n�W#��R�O6�C���`'# �\�UO^}����<)����o�l\����z���޼� �ֶ�
%�a��;|��kk~�5�4�,�Gt�����+k��J�z�r8���-$8V:gH��(�-xi3����r�Yg9���H�����M��*�䁢�s��t�m.:�ZUW�*2�4��t�nq����E<N(������^]y�o+
{�	;'U��st`(����l��8_�B���;�2�K�d).��Ilq���^�D�;7E`;�&�b�Q��1")@����PEU#q���.\���u} ��l�^���~�R�FS�$���b�}�>�v�3]J�AkA�Te�?UE�*X�H���ݺ'r�2�,0^��xM��l����&�8`^������2�r�/��nK�d���YE�7��(�_��⏏�`�×�ZU��d�UZᖞ:	�Z4T64�&�j�!{�]��KU�*H����zp,�z�S����mƦB/�$��Q����M��-MDe�6���D"�B������3�j_#�'_w J�l�4���󁢞������|���Vt�%��C�m$덠��Æ��G��M�'���t������F;GO~|�<���՜��`��&�Fs�AK�w~^�BN4�!ոwAVgd��$b�+��8�"|9 HA��4D� BﵒJl����'����H�I��(�������|����|&t�F�O�1�Z�������׉q���C�������Bv�4��GeC��a�����"�V�D`���G��7�=�X�1���FYX��k����I�iy�fɵ�����:����)�a�z���K|�w�i�\6^�o���_ѕDW7�h]����ڲ�������4*���?l�=�t ����Xcw����Я~	�LC�LW�'�J޹1q�&kHʠ��9G�ޑK��2�f��ꘇ�#W��${ޚ�q~뢥�tnE��b������� ����l�Pn�Zmq���irM.VmE�����L9A�k��Ӌ��*0a&qat��RZ� ��	���|��p ;F�?ĝ��%�����ϝ�LIk�CS��T'�n�m��S��xD�����mK�]sUG��#1VY�h�W�ԒAONa>E%�����یl�[D-kl�SO���
�z�4d�2���<�+�/(��A���&�A�vo�x�x������n��eH3�ɼ��* �O,��C������Ƅ�~�lT�@��;n���^0D% 
�U@g\��ݒMNBQWx��<\���΄�I�FVFŭ^��m�O�V&�4� ـ4��rx���Z�d�NI5y����H9���m�1Ƙ�I0��S�Y��)L����aDd�U�����_��,�;�3�T��V�ۿ�]	�_����yC<��ϋ��R�Y`��X�k�t?���F0	51��5��o���4JPZ���v
>�^;���eY�-b9��+.
��j)upʄ�U�&$��n`����6o�wtL��^}(=}��Y���aB���7���5������Y�ᆩ�Zg���7	Ԗ4�,���E�^x��"ާ1�!Ȅ�K�s�`uNvV���'��(/�(l�Z���H�HJ�Ph����_��`L����M�����)6��GҔq+��=�:���Y�hRY�5�ʷ�=��G�ף���(�뽠hp�I���?���[�K���%�S�L�:����X�l�Úվm2VJ�f.u>04���0\���ѓ�ůΞ�^a����΃���Ǜ����A:Zo��S�S%�s�������� �~ż=i����W�$75-%�BQ�Ѷ���q1�n֧�&�.W����rl����|ωn0��t���K�.Goe�8��y���ϓ�,#��*��k��4��^_�[�͐w`�g�hby�c�^>��[o�E�� u3�7�C�"ƈab̹���ͅ��V��Ji�"J,	)@C��d&��A�
 ����x(7���`��$h����x��XBfK�FjpԨ�����) �o\O�bA{�Q�Xv@RA�.��������\�H��	8)T�d,��V�8!�k��Q�ǁ���H�p��l�[����8��w��X	K1��`a��YF�H?�߯:�Tb9 %3c�W������vPt:=w�I7�s�����N�G�L���;	�}��tA7�F~�����25�Pu�[G�Nw5x��3<����
�����P-]��aO����*9��B�Ut���:�D�֣B����)�6j���}��T�����ϡ�S��(�7]��5�%I��CJ�W��n�2�FQ_��V�M��F�M��u铈f;�8i��t�A�,�����E3��݋7�\�����dK̲LnkyU[��)O�z����h�(��C�<���A �}Ձe ���ěT�<{��GP�i�m|{v<���t�SN�LI϶�ǴN��ҎR{ѱ���J��j���W-Z��e�!�5�쇀���`I>�V�8c�@,{�,pԕ
Q��{�E����c,��\h%��Wh��=��(��C?c_��.q	�d�u��N�6~8��?b��{se���;�ےK�*0�A��95�d#\坖�WFjP� W$����<ĉ��������z�'Ϊ�:���r�����FH��i'3�Щ�>�²c�F��f�5�r�\ #��ÚU�>A����s�ٔ���Ul�GG���!�&Y?D�v׶c �z�?����v@��L.�Cf������茕4m廭|߫L�/Ǣ�D������ �΄���Dbm�����z޾�1w�q�Q�G�,�t�R!]3�����z!�}��0\��H~J����R��v�m�)��Y����hX�������qؿzQ o����E0��z1�w��:�̿��&���˴ ���,��9�b��h��['��6%�5�ꊼ��I5h�˿sT�۞�)��u��1��O
��Ѣ��:��	G��;�!�ң�G_��ˌX�a4�-���v�⍒�]Ǘ�Ө�H:�a���jU0z2�Q呡`�%Ɔ`,g���=|.6�&>:Nz�O����B��"r9L7BZ �I��:E��`�����\^g���}!r�c��!�sS(l-��xD��ģ�1S�����6#p¼�k��sgLZ�6Y�O�w�O@�x[rTd� �pb�L,�|u�����c���g���4��]	V~څ&{pŲ��P`Bw���^��=Q��)�z��v&9�����d̕�k�����{��>�=����$���1h�8��?��hMj���l$#b[��/�X�Q�e�HP���ʬ0���?��������n�٘5��o{ǌ�yB�pFP���:��ͫ��7W��U��RΣ4���tiB=C�WY�mγ_�~�)5Z��H�P�3eg'�ZN�Hn��E�I�a�=±����)RoO)fD��%F�"#�Y��E��g/�8K'�I�)�� 6/K�nm����Vb;���(���;�����d��_������l�O�F5*FD����[F���F�{��[�y"8��X�'�B4��#n�9�D���f��N�9���eq4�/�� HW��j����~�O�j�{_faB����z'����Y��d�ֶ����v<�:ND�Kcb�S4-b��4��?w�'e <)hkB1Q)�:�d�Z�R�W�J[�qZ�E�o7>��R�z8Ч�m��hCQ��۷\�I�5�(e�nL3�,t���U?j�NDCuPRńΤlYXN\F_I�A�=�
�m�{R���!�q�W��
u���	Y��n�=�q�G�޵:��:�2��A�@�_ [�C0��bW젙_����f����D^�L���u4�1G�F�����{fvVM����z���A���y��a+S��a��p�!�j���H��06a���>o�=�����P���
<W����˽���#MQ�T��I�P��&���.��	@΄Ɨ��>;O°c��]Pf�:5���r���|l��z�F����^����
;��E 5�Zu% ~f���[�J�.���5���>8�rH�^�Y�i
S���i1������+�+#"����� ډZ��#���'�\�'��!��!'�2>�`3�F��lh�R��#����/�0IՈ
�1�k���J	����12�:B��
�*�Mt��vẋ����y�P@��l$e :8֞�3��y�����9p�#U(�˕�3o~C�C�7f��vD�ƞ���Tc����4������S��Q�&�4r�=�\���������#_����ҕ��<[%A�t������e�hU.�SY��. �����.�0dJ��1ͨ�.�Ln%'���n�V��9cKI�R�����;���bY��5��\�;b�����>�]?���5v+��^��N�\�Y?B����p}Ԯ�ŋ���DkQ������}�����Л2+Y>��
���<�Iةߺ����'���x>Y���h9@�@� ��S��a1���QjB�/Ґ�;��������`c�ד��>��rC�>"KZ�����+��j!0G���&�j��W�="f}���{�ArF�py������2#)�sNE�!��"�1�"g_oG�Åe���Ƚ�凐�j��m$u���Hڀ)ߙ����Y-ʛ{��R��0��uY��fm�y�ʱ�ȱ&�np�^X�V�e(�kY�轸S3�Ω6C?)zv��L,\�n�p������c�<�6Qu9kI�&�`�9�2mK�^�܃
q}+A��9��~�����t���>?�c�r/�%��]$�{Ȋt�9G��~�#��N�m���ݳ��T�N�k�*w��Q}=��_���,B8O�V�ᕭ�x4�O�N�Zw�®U�;���E��Z`zC^"������%k!v����=�������<�#�	���XaOo�f��CR�@J��c�o�l�',bG_i���|R���4��])(�Ss@Ƶ:	���m�X����rI����^n�x��F+6nm�3�:M����ݿ�ļ����d۶�����ث�a�-8��J�7(�������^��o��e7��'aZQ���u�Ƈ�_/�y�Ё�8������7g~�x�Ȋ�՝���
p"�{�����q�Ŧ����D�zi�3�R�3�\}�J	A�W��|����i���[�|�"��A���i˛rn^���}S������j+ntIX�p���bQ��N1��.\L�ԉ�n�$u{|��(�
4�?�i.�3q��%�4� �b-R���?���e��k�t�|k*҈�/���&Uj�"*�#� ����C��,�v>���5�彥�Z[g�3Srܼ:�;���\�WJh R���:U�pd�Zr�z���䏉W�����0ц�cõ���,���T<�+X�]�'hc@�F��&|��F���-���"ȏ�F+c�>��ρŴY|kN��\k��[�M�n��xE{�ł={��p��WUr�e���@�H��5�=�0bg���mͣ�\7�D��Ż�2��+}J7�c��S�o�Q��!��������{���pQ������qp�'�lS���[�PI���r��cZY
ॗ�Y0��
:�;��q�����Bda�ӡ؄�?V'n��p�_�0>�����8�ެ	��\�ݛ�t7E�/W��4{}~c���ii�C��^�+I*~S2�q�3�@h����V�R *���*m26(w��̧��X�ɧ�(`L�	��򚒒!E��h�/���Ci��Hr)�̺��[ؐY%�!�Z)"rO:d�ö^#7ָ��	����g=�/�EbĹU��	���H�r!Ml����}$�gI��h��e0��c�����8O������o�zUHQ�(I�o�U� &Q0E,�O�C1h�@j�M��t���O��{�\�Tt�����^\��xN� ��?H\#;����ت�^�h$�"<���W�pd�p=��Jg�O�L���5|NR�Iʂ[���Ŀ#Ϣq7O��}m�F��t�1������eZ}��w�.���мX!$�2�U#C5�c�릉�����ӐֈD�X��>&�X�|+��ء�u6�;��Fd]�����S�� !Y�g���P��fU���xm�>M�y�	0�#�pe������c��'�uO�B>�M$����dS[xE�.5/�Y1�u�0
z�B���[�
N]6�ޫ�']��4�To��D'��`��4:���Q?+���e��Ӽ��Q�QIUg$M�a9T�޽u����1��U�-���K�]����ݿ�+g�/̹���"���L��������mА*��\�I{�[7����OYhF�[3.�0L�i�Ntł̤j�)_����Y�l.��	R�A8Y�[��0b���S
�ĳ| p�s������!��=C�g��e;�oBI<��[��nrX�L�NĮ-��"��y�3���]��D)	������4���6�&֕Q�*�;��~�H*�&g��K� ���KqQ�p�$z[3�:�8$x��~��X0��]���
��P�UK�(F4fr2�^|c7)r�1�#G�c�ߏl���ڋQ�$Nc���jؒ|.
z��٤��:-7b��$�=O�H��i���F_\:����E��N0�{�m�	��ω��0�jY�8�H��%��J3&�>��0Z*��&D�$�TM>�%a��C5QW(ʤ/|�o�oО��KO�O�́�,��z���,�۝ ���+�V<rd>n*�S����#e�qW ^��ǯ������!Axu�'_�x��Q��E�n����<�p^�~�f�ψ���08R��/Kx �n#`45C�v��/{�݌��Қl-��!�7���߼�!��VE����2q�ݛ�G/����T��!>�G��!�;�����I;+��M�7E텿�5v5d�p��|N�������q�ˠ1�wIx���$�4v�^x��j�nw?D����/zR�=P��O�=t���?���*<^���^�iX�@��W��
���"��8{���K���$R�~���l"K��?F���(: ��BX�/e^�l$�r}JM�)B���2��G�ɔ��A�}B����U,L�5�sK�2��P�k�W���-�����������^�P��"��]58%�[2����P@�!3�V�7�9D���C��ꫧiO�琞Z<h�_��P�|��<K;!�}���pc�(�
T���B��(��Ư�\����s�0�&�%3����*�֒H�q�^?%����]=�-"���jj̴ɢ3C�u����k͆�a��J�t��}��lgp�a�cJ���L�F�2���Щ)���� �/y|ZGy&C��`oIr����$8V%���Po�H�%�]���1�2����J�雃6�6��:�d9~'�5���k�����Ʉ���NKZ����tuH���� �]G��<+��J�8F�Sr��N��)�d�HLѲ���?e����b����~�c���,/���-�=$77p������敐���Kn��8j� ��`�Y�:;#&iA�{Jzwbkl>���>�3ù�d�)����f����|PmeR�Ad�k��	h)����5NAzv�8a ���us9�Z�D�!�+5ӇfҸ}��?d��?}\�]̦Z{����7�S� -��\�Ob��O�������,K:Y_���>�fBN�ɀ
�	�l�	j���Z7�u[KJ����@fJ%\4.�]��(�� q�o�l�wTD�*�a����,5�>�Wo����ȆX݃<j�?��l\��2e��©�S<^v�J6�1ы"�3\��pϮ�HXg2�w���{�Do�n�U���8M�l^�Kk�*�tT-�V#AhM"MZ�el�&n�Q�+�˫��&����R��(�/�y�}�%!l����"�CE,�V�A�|#��u��0�} ��A~�lY��3���0~�l�w��[C�7�+�Ԣ����@!ϡ��d;BS=�0���#fr`�?>rU8�Y!�����GxZ�=����XO�wL弽6�^�H�q��uI�'����fև���Z~�w��I�"]�Y��3sc~ ��e�+�OA�.Q��|���i:��(F��Z��Y��1�8����`�����)3�%N�++��ic2��KӐ!�ȸ��_�R����mg�h#�ҿ���������/�����)8B�\a��ٵ�*��D��E`�O�����CrL/�Y���9�挮���ԑI���;q[f�SO�O�C�|/�AB%mv�|\^�,���&��ku����Y��=7�1p�,�Џ�!h0���H��'g%My�'��%��IS��4�rt�?ep�;���[����ɰ��{���g�vK�-�A��q��j�\4�b��	�3]IhVZ z]t��ݪ��W��
��N��������k<f^?�^�N�Է}��*�X�#�#1&i�2f���JW ��eL�{͢�v7�rM�(��� ٨�y\�d�"յ� ��91H*�"a�>=$�-�=�֯����kKn�Ӑn�5*wlD�Ќ��XC	�� F��$������c^�^%�DN:�K�}|/���$�T����ҳߵ�HA�����h@��~[�Uv̐�#�b����R�����!Rl�dU�bJuz�G(I\����%���!�B ;!�d�h�9\aa��ٷ{�"�P�D�;V@�/Ep�S���>-�Y�B58q¤�倒i3P&�iX��NZ�,\P\��8�}Y"<�1�V�3�쾛��#�|Z_��g�����3�W�5��|_PH��9���"��iB0T# N�Z7^&���a�O�9�)��/�|uue��I[j ,��Y�rŃ��s�,��ю\r��6ˉT\4c")T!W��,�5�6�;ˀ ��O:߬ps]�e���=�ኚ�D�ᬻ�\d�1w�l+�q|U�ȧ�dgGl�����<����zn�6 |%h�߸1oA�n�[°g�'V-�q�;:�Wk�H�c(��st��b�9�3NI��Ax�R$C�z�[�mY'�ֹ�06;�7�a�nG�o�`M?���s-$s9g��"RiL��I��ť�L�Z�Ϋ������<`ux��H��O�n;���g�=�2��mI?w-js�K`L�JO/��|���)��x:�+���(/�D�,�ֲ���7�^NT1����gK5A��м��~$�٨���}���\(O�]�����&Hp��ҿ��Q�/�;W�L� �ꇈ�r�W�n��%VF�ӰM� ��UK���+5��MA�gy��ꨧ�B)����=<v#ej���+�0�m��T��=2[����Q&��W���r �snp�Zvh|�@Af���uBR;�]� ��y��3r�TD��Z,��熾x~hd�<Ֆ�[V����L�T�$�q�`Z��uܨ�k����u)���,�=�>�OX��k����a���!�j���Пd �m��j�3���
�p�� ,3'�þ��l�N�̑��[���"d��zU���kjxΓ C�j���ak�[�M;L���O�AG&f *�`�,gD�:�C�ڲ�VMwJG"����B7M4��'�f��P�M"�\����ܢ+�K�턋�'ųS����W��%ɣMn��A7+eŧT�p�Z�]����s���o����R�z���ې1"P�'<s]+SP�"���Z�r�Zr<=���G٬�	Jt>Η}"�5�;@�x�(v�[���\� K��>BY�ј�Z�r[�צ�v�I1!�Oh@1v���8�Κ6�;Q���%F�?�_��.ŉ;���V�ܜ6�����a��w�n��x����9b%G��e�~��O:p$}i�(u- �ň���m{eM���I�6����N�	�+q���y�]�7��Y��!���z��Q�V��W*�0�~�� �)���h*����c)@M�uJ�d��,�ǜ����Z�C���z�D�茼���&�\�>h8�z(�6=>��,�z����n�:�A�6��,�<x��+V��1�P�{7�]�ߊ1�+��-���.X��ZXc�v$��������=k�p���\�^���jFj:T�������`�Si����tT��g��/�"Y&�&&B���ϩ��#��<�p))�Hgq4phs�gd�h�8�w�IM���C�+z�&C �29F��I���6�4��+谂��^������^5����#c�:9��Y*�[�j�j��Ĺäf���H^p��
� ��3�y�y�S��ñ�Np)�-�� {�ώQ��7Rc=����ex'[�����I�x�� p�q��qi2P@6�#1̅1gX3�J@��$��}��l��Mՠ׶x-�'cMƖ�V�"�\l'S@�Mq6ԫ�ܘ�})O�CK��0Ux{�Ҟ�F�0�o�w��1-����h�t�g~��>i8����0�Eyh�8P��ezy}$�/34�ha|gx�A	}[0�&��%lO�LTFojd	���NyD���3��G��� ;r�"8�u��N��Lf��+<©p���	qsGv�$��Adk�֦�)��a��Zʡ�L�;�7_\48!-4(�~Cu��@�X:��7	��U���!�t	��j�:�^78iG-�L�
ß��j��ҫ4v^
ËF����UU+e�G��y��;D����S#-
�*3���茕���"�%!��s���0�C����J[%�J=�X`�G�����RSE���_*d��g�9�%	c�Ef6��0F4jP���M����`�W�A��h1*�̢{Hy����א�˔ U&l��<M���>�Ԭ'%���ğ�l����9t3-|��d	�>-�L��f �C�L��jD�XV~�>Yԫ�}ؼ]׾�y��sz(�HI��w�Z�g؝�5і�|��	�^��Z)�E{I.ղev�8�y�+������{9��[�˕���\���,ࢊ��@H�7�s���۽TAe��t�'"&r�b�u�1�D�u�����g��S�]�#��W;�U��s��o����~=��b�-��4z�I��Y��@5	��) �;%A̳�}�/�8�$s���#��+ �f?�,σ`,s(D�%~�x4�N��3���<�,���k�`$��܏g�=����n���i�J�V ��3�Zqۇ�|�푒R��.��g����I�M�wr�DC����P���x� ��R��)�^i*�2^{����l�#H3�I�.	��P���M�m��γrd{�����L4�C�IL��\n�K�]b��s�jҥ�6�3��=����R.f5]J��|5��S�+���3]��S4��e���yF��
4�i��0g/y����Տ���8!�ol���-�@�1��ǵjvi��Kt������:�.�mY���Sv��q���᳙2$�?ktS`}=�`ڝ��i`@֤��%��c�5hp�M��6[t��];��;�����s��|&�ڄ�
��!@��]�����5ڜ2H��0C��1�ݎ	ۗ�2oB��C�@������kx�\��/918a�P
���0P�� ��=�q��x~N���HY��_�~>3x`l��'�59���S����i��pxe�L���}=p�
�gq�2�A���.�G�[=>�ҥ�0E�r�g��E��i�qa筰��%�W�xҖ6HL	1�N��h���95���׶�eq�B"��ږ�+�86��B��N9o��=������ֲGe�����7p��w�lز�].�PZ�����f�i�����(���D�2R��][5A�x�B�d�YЍs�&+6:}[PH�o���'sK�������g�(ipͰ��o+�i�/����8�_	���f�/� ��V���.2�~,��su���΋/�,�<������d�B�����Aآ��K��)!G�k/�7�ě�#*;!&�L�ܩDk�|�����T$�F8R�'���n�bd�S#�\�/bE�ܕA,܉.u�:C6e�WpS��T��a���/sALo�>���[�f���6.H�
u��H�U��M"�J��_*,	�Ogݗ�=�?����$E嘹On�*ݚ�<0��WH^�r\�(1V�!�o����y�bC���P)'�Fu[�C:`K��>ܤ�X&��T�hm�ɇ�C�$ �ᦅi6�^�ȫ�_U
�ۅ����= ��Ӡٱ�e߭K�}7��#�!��)��ޝ���������B�w��),9P�?���S�����U��W�o+��������%@�a#��t��&(�!=�uuX�q�M<�&�)[�w�����}B`dz��A�(d~{�L�mʓ�޳?��u�4�m�O$n�lJ������&�;m�� �
s�n��ؤ�Hoϐrwv��C< ���=�nv_T)������?��̋�y=Il��G��9��0�~�(�`b�{��I�5������6t�