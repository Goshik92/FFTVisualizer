��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]����
3�kÉ�'gP��o]BSt<��(:�qB,]6K�����Ц���0�ݐ�������I
��k�:J��N]��} b�w���m�pR��-�V�j�<�� (��fWF.;z$|�{���WvB��&�\����"���la�0�hJY�YTר�FZ7�r<����2�y��D�Uy��?,�<����jN�LJ�L�ǄO����
�F2���KB�"h3�RU-��p!�ɱ	x����2�-��3I��@!��O�Ia�9B�@�����{�qq`�������o��éJ�#
�h��}Y��q0Ě�ӊ꺙��m����������o�܌k�4��QmG8�=~��{�7J
�<+X�)�GWQީ! �{^�a�_R� L�Z���F�Q�7@�-I����v&�R<ۓf&ەbԘ���i��E�3�C<T�F�@G5���!HN����D~�A%9?�+i��C�G�r���r�`�<!��n"p]=�w�K�JqKG�k���{,�9�� R_`2�S�|��p�J�ɿ3��l�#"�\���}cP���=[�Ɍ���4A�h$�;��	��3��F"oD�"�Wm����W�H��,�jl~G��Xv#��g/*�`��y���O`���¨nNj�T��;��2t�FjA�0��!����F�ع��?ć�ȉ��h�f!@�CEBJ-����L�Kں��S�<η�,K8^��3�"R�(�d_f*��<�E�t��S��k���#`*4]�	�Fѝ.�g*���T��(���~{Z���D	�네�\���A��lz��@wV������n�wt`&���k�}Hk��k�.��\��i���8pw��Qlޫ�>�R���7o����dj�k��>;ې���u������j��1^1��.=���/B������8/�a���5�X���M:a�uSV�d�i;/Qe%��#%�@Z=^6�:��r�i���"�偱��B�����>���Q7����Zs*�6{�֔j����av�r(�4�+V\>�o0�1y8�w������&aP]�{O�骘���wjIUYQ��n~��}g1m@3���3��oi���jL�������,�Q��|�lխ�_p���u}�i5�H�_C_�Ŗ˧=�-�Z�N�ђ��*��2��.u���L����H��f
,K/)�c��M�FbM㡒XF�60�w;e��x/�M7��!ez�|��x�(%�����pjA4����t��(mh�#ҤrS"���6�f� ��q8�of��#
(`�p��z���X0���$�	̠|��`���$d���\u���o�k���d��PV#�QA��,�Lbǭ���wh�4��,+���qo��Uƒ��]��ɴ5�4�#�+�j\��0n�f�����V�tMYsohs���8��,c�N��NT>�7�I�ѧ�ښ^�0�c\�`���N��˧	ɟ.��Q�v8L(�[����۸Y̴<����C!N(�W��˾�_���I�l