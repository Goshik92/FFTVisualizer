��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��do�F��ĈMz�>@\�	U��f;�m0P�ѳ���Y
��D_2��F����ݨ�4X�J���̓36E��������m�3�ұ�E%�?�5���U��^do�1۰��w&��B�<I��A�,��հ����aR�UG!��@cC���4VO)���P�s�[�ö��e��2h�y�V{�P��W�% %]m�u�D����kӌ���9}&<��Q0��/��_z�<!�J�BtVh���$�G���⺷Y2u��"���>J��BAC�������u��٩�>E�b��5rQ�m��"s�+đ�z�f~��#'y�!�����˹��o$�i�"��RB��~��8�� �	��Z2�~`3UH�;.{�_d)K6-��I��+-�0�.�Û���VT?�Pn|Ϋ�g�~��:���N��']J"o��aH��?]�����3v($���X�9;H}�����8�.�tE� fU���D���|�!%�����!�*�=)�� >���8�eBf҃߹\=��!K9ܜ<4���R��!^��� �a���]g�]%W�rU.&s
�z�;�۽I�r�L�ip�m�p �~����V�Th���)��l/�	�-؋��re�?6��\H~q�:1»����8�Qc��V�p�I�i�VY6���k�������x�6��3��4��%g������\0OVzɲ��yIů͖��-n�!�L�4����
�mӴcU��b�R>�������
�J��6J�Z��)��2���dx~Z1�mz�0^�]�h���Cr,��aQ�A,�N<[���-��K�y�� A7���NWU�y_���]�b�oh�ċ��gR�}'�Џ�I |挥��0���/^������`���e�Y��Q5�п[�DӬ��lC�$+��]ˠ�������č����Rk(Y����"������`����p��P:��9a�Z��,�M��'Lú����|n��fj&s(�1gx\I1抷�4�8[k��oQc�A3�f�<��/(����@K]K��@��f�!�4��&�V��7���e�L����n�������G���W6 h]T`9�p��9u(�"��$5�l���� �{1	U Cx
�wkG������9��f���O��E���� �kG���S(z����#mq]��R��S���;ۏ;�y责�+�p�s���G���q�fq����DI��������b�?I,���wZ$�$D0�� �����8x3Q��x,63-�O�Y|�,��-���t�������V}�m�t���QxQ�,��/Ŕ��v���O�H�����i�@�y�dpғQ�@��KL�Ɠ��f�T*�d Ʈk��7(7�,�*��֬m�B�S����qtSXo̿Im>A-�f1���������̸pD��[G���(SB���ı�B �� �����1Ч���~�N	�V��������e�+S�� ��Ƽ)�W���}�=RּO�E����\�4�� �@��/��QVF2}�dYt���G��܁�b���+�)�BUm�W������_�?�;��Fc���Ћ��ι���H���Z��+�OS���TAL�ұ�� W�-�{���ǋRC�b3���.�{�4�J����y�M�Yj�h9��<'���o�6<=�����>�����4���z3�����Mց�D�E�eȹv)G�J2�!=nk4�~�T��_B�I`���rv��#,���0�g���Ȍ���n�W͊��U����� ���MW�K
n*4L�P?H9,��_�5"6bѺn�L���􎣚���q�R!R��oY����߅�b���6z��0#�A��,�����ʽ7r������9��dLHV�'���J[	Gp��ue���.|lֵ��~���
����P���̬��5w�V�5,^�Ң*^�+	{�=��[����P9{�"�2��dt/�"ʙ��H,�������%\.c>T�%r�(R�W�Rlx0�A���T8.�"�L�es/5�W�uW7I�%Gf��gu�1)�T�&�,l��/W��]��x��������hނ@u
K�l��%�&�����C�W�e.�����m��+�@-�10���da�r��\�/�=F�?H��V5�m�cM1�6�s-�St'%��?�b{�OK�f����A�����\��N3d���΍��Ǎ�uf�umXl)���l�p�(1�3P��7!�'�Z�v*dQ2���T��Xᇲ�M��AD�*c"��n��g6��g�Wb*7kd����D��xdsp�#1^!熠�����5���R�4I�g���*��M̛�rLc��Л������ט�D�&oɴe�Yi9����H���GL� �Zƌ{����� ����}� K!s��;�b�&��_*�Z�#��ko���_r����Z��A� �?3�m�>�����\�K ��'	�4'�q���]��0y�k��y-�6����+���5Y�=���\��: }31_�����B1�ĸ	
�N�۱N�ٵNퟴ�O���L�A��>:��*�ʼ�q�F�����B3hW���m�~[=��w=: e���v$:�M'5�i�Ҽ_"8���� 5�mc���zl�eճ���i�f23[���3���cb�7�]�,�n��F�V*
s*hG�̇}u�Hس&�Oȩ�秴�3"YXG�Ͱٸm�c<�j4��wv�#	�X��P��qi��h54�����;K%y���?j�(��BetˑNgm+�s�:�����½�?���s;Y�8��	,��v���Pׁ� h{���JGl���'�QpV�9���|�D��f3����:�1豹�j��h2�,t��@\G.�U�5�~�s�S�3�vx�r{T�p>�@&��W�E��_�p	?��V��|�wL���t'�`��Ľʏ��i�3���}F3���.{؉��C���]��~��rI���H��,d��n'{�O>�U.�9}����ڑ���|�v�jߣ�U�ֲ��42����&��2$T3�X��>K[�S��1&�S��[R��cbbϏ� ��l�~��x0R�MbF�`�Pn�T��m�����ʊ:�b��t��_�)N��3L��x�a�;�w�ۛyR�J?�ŇN1�J�LQ��!߅�q|}ؕ�+!�8�M���a�{&j�+����W�>�o�I�!N<2�M�@/Nkȼx��}rFy$h����2 �|��V)~C�kr����.��B��l��IR�,8kCn��)��aE;�˾�4�}�����?�J0��M?:vQZ�Rn�hd�.VTP�Qfдx7c>�G����x{T�!Dgn�n��\���Z:n�d���%���k*��b}r3�0)U���Pؙb! *�>W3sZ�j2���Q�ߟ��"w��W}�Yr�u�oa���?O�� �ϐvXuv0B�l{V���t��
��r.��7ď(�֋����0#7��(���(�C�(�O!1Xc5�v�l���L�,ӱ�/��"iF3\�4�Xy0����x��� 
������;�!��uybW]�%���G+�7�!��i~����S�����X��}���D\�odt���+\1�%lVZ�)2�=p��=�t���Ї'S�C�hrӿDM�u5:�yS�I�1����d�
< ��i1]���̍���⤘FM3�U�������ֿ��e
�NZ�f�ʛ�����Q葦��ie��` �k���B2��x�v�[�ի�^�)_w��ۥ��QԳ�{�*����q�|3'�������_�ȏOt�n3��.��|�\"�H�����At��-I`
�|�Lk�Y8�JI��w(B;�\F"ӓ��j�����Qxr�V�����f�A���W��?�A{�4�T���&Pofkh~9�K����������d�Ė!��vj�x��i�%�!v��e��gV+ds��˴�Qk\a�������esl�+���_���oF���M*!�c�̈́�\A)Pe3�8��TTIƶ�L�?��l"c�,ze����~D�����d&)���Dd8b��.��|�tej	� W�3���wv@��r}8��r#k�7b}���tO�=fnDwn�<��B����Aw�s�w�T+����ӓ/����/Ϭ���zc#��ǥ�\���e`�D�.�*�p-�79Ҁ���z4��n*�4(�����V$�I�Uf�	���WuMr�_�2�;�B�
j���^���t9fl�C`'�H�rt*��Q' j���|}�0����k�'E��6�TlUgd�"'�!���9�����u�3l��8F3B!�e�S��>�ǀ�!eڻ�,���H-i�,5�N�����������>Z˭��@�������.�r�D^�A��,��ފ�
>-`p�JQ�oC=�idI� ��i���C�nd�^��A�J�e�����T���3�Kz��%�FoQ�J����_���-H���� ��t�h��
F-�V��Ϻ�/�{ck���c�Vw���C������I� H�wZ>/U 
�]��P1x��?+����r^�i@T����i�T���y�&����h%v!)-����/ ��q,ړ�w���)��?��ڀ��Ͷے�ʹ�7�q�v'n��P�(�0����i(6���G�Y|֡ipG���niT��´�ˢ����`�~E��{���:�������~��r?���b�qO��Z���#GM�>��6x1r *����}����H!Z���F��Lu�g���4i�<��G�E����"�_��(���u��X��w�E'��0e��������i�T}.��_c�m^"�¬����)!#?H���"5B����M A�|@�;��n��֭ы�Y?�f��*�=8��*L��0f#�YIn���0��FMe���
_���R	y�f��}��KR�r����gɪR3�1�M?����:jFz©P^`����/�H��˷\�_n�^�xdl{�U:�}]��5��'�RA�"�@�s0�"��P+�r�_��o����7� 7(u�XRwb9�,=�hH����Dk�\�H;HH�#��6|waR�ؤс�������ӫ=?l�fݱT��T 1��6z�w#�"S��+?H�E�(9���zM�˸�G�evE���_(����2��O&0ͅ�T�c5Z6���PY��g�-���@��[}�w�n{Ӈ�o
����%�6��E]�l�v�f��]ةu Ң��k�P�����E�!4�L����4��K�S����w:�e�`�s�S��?��6)&<�Ni_3�_�I���[
^��Xd׌2��/��0�\o4#��)H�OtsQM�̋g:�i8��L�N�.4 ^l�H9c�k��֮K{��iT�̭��#���k=�CGj-rf��D��7|Ui��[ E��G�:N̊mT��\U�E(�R�ދXd�U��!����ۨ���ގP���6�bW%��iz�D��C%�i��8 ��a�H��, �"h����Lý�z����[��p�٣���~.ȊW�1�Ef��} K�����(�1�  ص�u�Jϔ�q.ž�:��i=��m���z�Q*4O*���&�VM-�@l���S���N�����P1��%�B0��r�i���"���m�Y���Q�^=`�@W�����y���a)���S��q����_���j���ni8ҟ���ݘ��+fL������p�< ���a��=���kfI�V��<��B��|\���s�90�����C�����7<�H�L]bQ����=�H��z�ּ}����%Ў ./ƼD.{4�k�����6⭺r�0��A&J�률�؏ߣ�`�]��ė]��[�`@i��X�/_���|QE޹n��X��������M��"!\�!� @n�P�(U��I�[e��6��ȃUa-��C�FO��H�^ўW2Ô�C韘�����Q��F��S )ao��:Xު�+>�ؓLȍ�/;{t� �7��,z���ȋ��|� ��to4� �!���O�u�m�$���S�	7p��3]=+��[�?3Q-�_���hl�=��&zq�YB�9Ց�Q�~��-��Ab�>D��n苢~%�9�N:Y�� ]?�Ɍr�o���ݚ�*�j���2�~��[�8Z��wS2v�uR ����7�Ay�cnm��"


 Gg3�3-�/1�8��RN��?�O�Y��������}EE8�A)�t����/���k����8��5��Gd3)p�� y��|B�źPٝz�f��"/�5���8����+Cy�7�J���^�~h� "+1I����&o�݀����k��B(�8S�dla�Mk�P\X���(�?�4��"���/�	:ä��j����|.,^lX����{E��b�9)�Y(gm�I�2�N�}�d��kĐ�
)2ZdW�lhs�����N:��>y�/��s댊�U�SXͅ7#��*(����e��,�w$|]l�O/�� �-�O�[|�����b�i����/���H%I��[�9��4�?DM����<i8����6�U�V,6T곲���ҿQ���?�MoY�~��cW�&x�6r
&+���@��/�E��-�/I.f�n�ފR�{��"E�����栺#ֈ1N:M��!��@��L�I&�ʓ�@��Yko�Wd���y��j�pF^�����Q2Y�EfD�F�Л�|v�I�Bf�%������O��F�?&��6-�HS�흈�����J��\��o��Ү�7�yTp)�9ԓ��Ƭ��ۡ�6 s�_�u47����@<{�G�4��z77շ�/�:v�ޜ�@ew*L�iJ���=�<V�4���d��%�p��\�]3�$-�<�y��ha$x��:���!.$ݖL'�� �)m�..S��q���a�ax�d�1���ڎ�Z�p�
:j��ϭ���V��jY�A�:�w؅8��&N�ي��(�E���5V���L�4����,������9�O��1���]�Y�-��vr�x���H������K�H����l?��FI-ZraӵĜ�J�>���8W�sj|���5�7�+B�� <�-{r�\����6�W6M���pM�N~i�cC ��;�̜��^���b�
Y�-����?An`L�����mR$�Ng� W`�~bc�@2��Tp�_K���x��-�����O׽&��:;4,�J���ܿ���[�,�a,�D2�{��4�y�ȡ���Ѐl3��%�E�HLC�[map炁wfI�~h�q[�N��M��~r,G�q����R�|tr��P����m�8����+��2|:�R�P�Z��˦Pz��@�jʝ�.� �LL�'ɯ�	eb��"�cۨ����_�W?`�*,4H���]�c��!������sN�)���O�G_xw����`	<�R�%���	�d�F��^����a�2��;ʟ�k5���1~2�6���<�r*%k0i�s�����u�j@�#�Q����X��?�^�f`ӱ�N�4(���֛��������_�@��{�P��\�ִ̼݇�fV�%ҁ7�/�۱Yv�x�`������->��%?��B7�Ԑc��8[` ��_����^T<�m��OT��:k6 ��/c�ρ;�H�[}�kv���/*휖\��oދ_`�j��:�K�E[<��l[aQx5�ޥ���Q������^�N��<�MC�B�K�s�0�RZ?;):�9�O�5�y�|�S�V~�q���Q!>��H}A�AdH�"b�aU���٩���l ����+L�fu��tDVJh�"�׀���w���q���w��Я�>�NH(r��c�d2M�/iL� ?F}�*�rW�c��lk�C�S�~�$��1g) �{�i�o٧��=�s��F'�|�+����M�	�=��|����v����h�;�A��V��/`�w|f����-�	'�������0��}΋����~a�D� e��}��*�$��<%O2��j0�l�<[�h�Ȼ9o���Z�A�A��I���#�34����8��AE^�q,_aX�r�m:�6�����ļ��>r^�dc~8��:.��P��ll��ip����fI��ZF�/�.«�Z0<z�d��U�} -�	Ōo���!V@��0q>{�d�/v!J��;*��</�Ǟ�~�_ש����#:Ӧ(Z-SA��W$-���Ū�𐧳�a�PǱ���OS���?qR:D;��)6t5�	�#�1{V �1Y;շE�C��`a�����&�L?quYj��J�4�����9/�8mCfuz��a��
T�����u��tڦpʄD6OK��iRTd�;����A-@X�3��^iN�BAy|�r��M��J^1�=��Hh �ƶJ�o=%�G���lو���/�)ʬ�v���[:�d	c֍|h���,�L!]3-3�VQ`Y9iF\�S��C�f�6ISs�5gS��q��&(��r�\�3vctLP,�<���s�y�V좔��؇�e����+����1A�c��G&�L_<x��7Z?,�O��F�#�������j4|է��"�<
����*!���l�'�.�$�]ifWA
έ��Oܺ�@�.���H�����r�\O����/D4�t��VW:���Fp���z�2�6_�1u��x
I���,��Ci����7l\Kz���P���N�I/Z�����NbD��3r���z�Q� Ӿ�r��DG�p��͡��/^��ߥ�!�O�rЬ�!O�x�Y��1�;��x󟇢`c�f�d �)���a�Q�|��*kR���s�p)Y������pY��� ��~�^��s�偵9 ��~r`�E���*��ہ���q%n\�LBǖ�N�$�D9�ʪS61!�OX͝a�?�2����t��b���mr;+������Z�x�똀Z�P���z��Z��"���"�\F�4&������f���`��øF%3.j�+�Z	@�d���bR�z6?
e�~E� ���m�s��#��p���b��J�VvB����?|�����Yx��O{�53��gz�������.V��Y������g��~�_Zݱ��4�FfEω�F*���rU�q��L�ϙ�9�����G���9���1�O�����v��Bɏ�U�@�t �Y������=�o"�
IO���=W1��7�B�!�� @Tfo�\����(�;D����Q΁b��)�k��N9����D\���PC��d��f��2d�7���N'�j��7���N��Y�c���Rd�|�.n��n�@���#�>�k�!��st?�ZPw�gԋ8�8�G<��	)1g�S��}I�)�D|K���R5ɓ��I�!��H����ze��H�:���h,˩N�:!L���gkV8
5k�RP�B�ȍ�C���攆���y��C�*����+���$�yg�8^
�"yjL��V��IO�u�S,�$�WI�����	��؇���4�f�,��؟f_K�,D�b"^a�$0�M%$����Wi<S���7� ��y��k��/}n=�SG&���S����\�;;��@^t�*O]&
`��u^��n�r�ý�@U�D�����?V��^1��g�7D���p��^H�O����|�C�k�?̵'��������珒Q*͒�����䅳��S�*�4{�z7wfR�������N��ـ�θkRP�H�9��ν�f��t�a��(Z|�΃8�"��4Ur���z5�T �Nss̖����ܻ���T�����{.ne\���,�v��7�~l�P�y�Y������v�I���Eu^=Pt4�(���� ��U9j��F���]j`x9���=�@2/�M��|������� Y������?�C��l�$� ��d������6	)=��maf�������Wݹr�wEX��s$�,�5�y��ض뙽Kw�����&qcD���n5�l��]h3�i�-n0]��M=��e(��-�]����;^���֎C�b�1dH���a��Wz�F]G:2غ������0aVϴ�
d�r��t��1��66��\�j�7Gr=���R�M����-ջ�
OS'ہ"�m6��|��>���uFM`d���A�`��a�e"��N��G�<Q3������M�Ȣvl7jU`�y،���]c�̸$���)/In�e(N��˼�7	� ���	�	�CU��T7�8wSB�Ա]8s��T��,����?��:)[�}�4�� �R�]	SNm�_��t0�.	SRa|�~_��I���Ի_;\�i�����T�>Kk���Ҭ��ݙ���C�)�׊X��~�ΌlPڔpGfY\^	e&�������7�c(��,/WCm9���r�K��r�E�8TVN���y���B�
%BL=[зP�J��Sݗ�� ��5C���yO���E��!��=ٽJU�W1�䲚��O�^\�=t+G���[��Z�mz��3�Lq-~m���s�`gyֹ����r<+���
�Wb@����׾�6�S:���#X�q�ۥ?��� z�ʓ���N�}�j�k@�������[����8���'f�Ϋ�l�rz��L�i�����EO�E����< 6Rf,z�� M�g�[EMA6��|��Ved��o�_�����`q[���ް�����x�C��j�b��1"�P[���487m��ͷ_] d@{V���WxC��-0񾳾��*��k�H�|��yS-Fp��*S<���C	����U�gI�z�㼪Ķd5l&�k).�@B%>�
�6Gĩ�^�g_�Q~ҨD-��S���Ȋ�ŏ���k#՜�@�s:x�a�t�X����-�԰ڢXKOf����TͶƤ�1�̃V	4�eܘO�{�|B귷�j)ܰ0�i���@%E�P5��5�[?��7l��E��4��x42�)X����Q����������&�@��F�4��0I���@��('�Ѐ׈l�)|MP�`�=#%}��0�3Xp��[}���T�@_"H��V��J��O�J��t-U 
Ij�#��y��L������u��l��T�7�N^�m���f���W�4�l�>�?�bW�=oʰx.��w�Ӽ��0z�]����!��~qf��3Q�7��>]��lv�{��*��Zk�Q1@�� *q��;=+^���
r���k�:��ܼ�9U�-��^�Iv&*��:�aS{��Q���7�.vP��E�o ��6:Hu��L�)ۦr /ώ���p;�8/eT6�V��Ϻ��cW��KNu���d���*�g/Aʤ�F*���_��ƒ�҄��O�v�e����'J��c13�ko�/j��ݸ�UR��Z�&U���|�B�< ��%�
����O�Q�e{��d���	KI>lپ�|���@�tL?��ƛF��o�J�S�7���}IQ��