��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��S0zz���״O�����w��듼=�yV�)�9��^���L��Bd@R�.rl�6 �B@�ßt�0tI�%[)d�/E �v���d_����A���1�*vpB���HZ�g���f���MR�����L���/F�W�v-;ƥ3�n�K�QR"�㖡�s�I�Hu�,
���)�+e��<j�J���� fa�x)\M��OR����d7�Vp0 [�N�t&\P@\�̈�(�~�(;N'E/2�ٗR}	����4�(Xl>�)���!��vSl��L��kҞ��o�a�ǁP��?&���=S��(�}�������N�ĦM�i=��'Hy�+[gp���.�?NH��E�g"�I���:�Kx�Y�2����R��t���yG?��br���w2�� _��4�ϰmOߵ2wР&dۂ��(j��P(?T�Ө�%��-�x��f�I��x�(�?2#!�k����� {����D
G3q;n���?_R#���*$7�������A�஥����g �)����%�1Lt��$�����onYU��Xt�+A���l/�]+���D���Eȁ����k$GNޒ*��?F�j��t���՝�ADHǐ*�+���'r�\%�ϴ�L�g��V/��o�����|�34,���"T�m���,��V�,]*�`�.������uJ�^p.~�MR����d f������| �)�o�Q]��M0��`1pz��ڦ_����us��C���}/1��{�~�mL�ܟ=)2�����==�d����&{�$M��X&��,���?�G����,�${-�L�Ӧ]_�S�X�ěf=�������ً��w�I��ɸ/�b,����/�H���mv1R��M��B�~7�8��;[Ħ�2�y����(xuz譏d@q��*u����������z��3%��c��:EN����U�=���u}	��I��� +� ����kt����Ȭ(�#Q��
v��
^���F���_����>b�a�����?��r;�'=)���z h�*p����{�Ư�>�N���G�6xk�tB��>��!_Oę�|(�ڸOc�_-h�B,��1�N/U��q���;EjS��Ʋ��V�U�:��T*�K3-^@�1�LV��=ͫr�J���� �V�Yœ�[�c�����Ϫ����J�D~�r�@������2��I���C����`���Cw��6��,tOT����]|����?_����R>[+��uD̬[�.ɖ	t�ɳ���~&I�	���=*9�z:aj�{l���F��&�7�V&�!��f��Hh�ȏ�C���P����A����9 �|j��٭h�fȟ�W ��竀62�0�K�c�C�kI�?j�����q�V��)Te�u�o�Ј��¹W�cu{��/�%e��^ɟ�V5��/�_'㎔�p�)����#O�At�C�ɓ����D�0���zC|�W��� al6������EBG�i�m���d�FIv��M^�V
��S���s��ڲ`�>�vB�c7\���r\ˤ��� æ4j�S�'�HD��ĭ~S�ٰ��rB��7E<Ѐ�I�	������bf�&O�K�8�����>�O�Ȁ$]�kg{]�wm�ۇc�C��B���6h�G�'�+��v�DiNf��%w�����T�xt
	�R9�aO�ǛM��`�,��<�B�#G��L�lٟ&*���n4���,k���y��7�٨�_4&Fk�M"�X�GwפWlV@�����C�|,g�gf���Vsq���aF�m[�q� ���7jm}n4�Z�W7�q8������=������0��ʌ���DI�)�Y3s�C�a`	XA�ν1�dW���R�q����t�L��B
�{8��X%siq$��M�@�o�-�a?��m}jRwL�ן $����V���p<߆�%&V�@��$K B��4��0���"yi�/�R���d�ㅭ��8"�v�k7���,x��V�&6ܳ�<u��� t�6?�&�9?��<Df�<V�1O;2�9U�-�V9T��a�O�/����+�K�[:�����%�((*pn�x<�ɖֳ�:3��Mp�Yg\9�����xR��
m�O2�x�B�t�
��s�#9�bO��ڟ��X0Φs�.q�k�o&�?va�6���0�z����wVsz6=H�:�S��s�G�;y?ny�M�:�0i��m��eu�h��E�]����|M���ܮ�ݽ�5Ty�ǲ�&��d8���)��Ȇ*���@�5fp%����M��jkl���w$�]�h�w �AVQx�~���S��z�K�[`z�9p�7�Y.n�'ZH���y8E�;���@t���F��fǹ�rA��{��<TE��v&/a>_��8M@«�m48���X{	�&�M���2?4�Ϣ���aش�8|�u�-�U
������H���+J�u� �x�<�I�����z{$�E�"@�J%����QE�mj��#k��p���y��+�
�]
{������	��R�F�t�[�s��<�G?%�QƝ��~}��<>)�у/�T�I����:�Cϲ�����rD&���5El"��,����,!&����)Cn��.n"x��������)�P��)z[�U��]��pl�[��*~5�����?�M�ht��8�N�.�;z��oSg�����՛����J=�b3	v&�7X�&�|�����X�Rl8�
@X`A?�<�Rh^�����BXV�|:(������旲���m~�k1a��끂���s=6�PFk�ع��?��e�B�{s碦��;�2Z�jr>
C��^�IFsɅ�� �Ϥ|��H��}�ݐ=hP��%������S�!K��.��=q^�@���U{#�v�!~�t���J��F��8�;��<�2�Ŗ,�o[
fIx�)b�BFTG��ɺR�v�X�>%������U�z`�8NNX7p9o{s_��27��$�YQ��He����
�����z��!Ə^ԩ~�֎� ���r�� `<�@Y@��5�<!��?q�h�z�/֏�_$������ރ{���^e�q��;Od��9�vڪ��sVK;{�^y%2�$ա�H�ǲ��)����ߊBq/d?X���r�]Ls�z��R��2�F��͎C����$*6��	�I�Z�OƖ�Q'�I!���Z�����%�K^�nÓ �`ԉ�X����ƣ�@���}��z>pY+_�Zv���Q/��z���>6Ϊ�#:�{�s���;�������6�A�N���	Z|�ʋ����%�j��H^�D�r��L�<�~�U����� �+G��Q��_��|qO�`���җ�Q��,P+GЅK��裲���?7�&J�M�I?�ѬM��}>9��f-�1���H���l��c�ޘ�ȋ>(C)P$�ԸPb�Je0N�Ʉ�������?�r4�-Uj��ڇ B2���Z�(B��mے^D���N=�*�P�n��>��Y�����l?)u��qs���晴.��x�|V�/ȑ���h�NK�89�����g(���<R��C�?���`Oߣ��(��%� V5�)߄�ۍ� �{`\��q1��h%b�h�f�eqIϦ�,A_G˶��V�y��4�� �����
�Ig�l��=Q{���B`�������BB�Ԕ��W���֭�@h�[d K�E�MG��es�؏4���8;5(���v�'èѧ�.)��3��Z7��ʃ��8F�|o�r��ڝ`&5'1�Ö�-jSe,��6�@3���А�P��a뭍�_�����p6t@(���7���jA�Ud@^����P(>,2����tVD�KX���h����rZ�/A1P����X��{<@ׅe���T ���|'��=3���Ѧ��OFe�W�V(��jłG���=	���9eu���ɐ��Q�?�x��7_;w&c{y�1| ��sR�sqMP���BD۴��so+�H�v���DRh5YM�S�Y�5)
�{���ΝɈ�td�'�'	�A��C���-\"����R�2�Ü�ͳ,�p
�l8Y�kRt#���e�O��0̕�M�>&��o ��,:+I��$��!ST��k�c�_2���3�sOO9��1r�~~R˚���f���!PCւ ��e:@"!X{���:m0���֚�g�`�v�OK�����F)F��!�yG�{Й[F�7�eDD��6x�z�F�?��ޏ�������O��� ���v����*�U���.�����|�䆕�[֐�w�ze����N�,��<�VTm�ep@K��೘a	���g��!���{2��b�p��u�ǉd�z�*v��5*��W\��|�b8�9g�,7Ħ-#�X��$F�i9�}�j�ׅ�3�}�%/��i�����v�B#H+H�[s�������e���3��s��V������I	��eJj�i=����n�\~�	.�U���l�����p34-׈��zB
�^Q6�ƫЋs��`�~�1�����B�!<N�i�b���/��o��$da6��G��sXMXP��T1��sa;�Ι�0�ϼf�\{=f�_T��1��W��n�<�aWw<�|a�`UW6vr���LP�!C����*Q ���h�g�����$Gް�0��ŰYG<�8�XbA�]��^�nY85[(9"��� <�/���=h5g�E�M 1��!�+Nn�'JJ�]�Fr*���hA���xb�A���3fD� y�݆Cl{�k��ަ��wztΤ ��z���S0������ހ�}�냆K�.�u`��۟p�06���1I�@�.��#�u�*Ꙇ���٦��\v.-j���.���X:�%�g���YE}�_��8J��y�����
�R	[D�S_�/'���vSn�l��-�fN�E'>��(�jt"�f��|n�hjJ��g�gJ|�s��<'��]����h��A�������+�nm�s�E�;��58�f"��Q�������M9{�j(���p�zo÷.(b��=�׶�K����C2��N�,��ZX�>1���7�}��~�MNk�ܫ�p	�8	A�!�r��Hi&�BHsfq��J����0��)�:d�)�`!�b%R������v��b�c~��R(�=�8x{���ﳢ��]�P-���~'�G_훍�������@E�y�����`��Cߎz���Kz 
�������nM|�����g����Af��(�?����,��!��H�� �_Wo�2qNp�.�n�=tGV�*��!��_
�q��p�FƟC�O��j�M�H��7����@,���4�I��O��&�&IN;����4+4�\�rd�����X=���`$!,���ϲ�`�?��X;�\���WR��R��xa��{��;~������}~��ox���i�m���bMf��!��[m�'��D���x�U��H�d��n�AU�1�����)���c�S^�l���N.!�:l�7S�ǧ� �]uC�)��o�o<�5z2!1g�/[��CʙV�{!��RńDA���J�|�~w3A�!�kY�*dk8��[�J�Ep5DþV�i��Xj��ei�>t��X��i$����w~�X����!�p���� ��ȓ�����h�)f�W����I�ale��q=�	:����Є�j~f*)y�Ӡ�s������&����o�@<(��]�"��o+)��9��sQ��:�V�s�` f����x-4T�J��&8�w�?�M)dI���\��3��A�A�9�o��u�$����du�^}}Njg������6A�-�8TVjXͮ�.�.=��#����w��]���ኢH����S|Ny�����Έ��q3KL5����R�����B��rk�{r�<o�����UMib+�|����f��@�B;x�R�s�"{?lח\��LPOᤸu�����i�h`�(��Ȍ�lm��ى��=u[�	�\G9^cv���,�>ƫ^:V_i�/��K�u�\5������e��ȩL�r7�I~�� �1����M�#���Ju�ƀ��";n0Kk��0����50�q�����R�������"��O-"P:�n1���9�U�[�J�
�X!�)U=_F�H6�csR�z;~���=�9!Ta`�cw)�\�}��JW�qg}���Q?��:���]�+`�6dI��N���Yc$?�ḻ��U%��5~�;�e�V�w�{MB��Zlz]���)�32�X���`�図�w���$�R��R:A��i��a�X1Jpӕ"M�@�c>���i��Z�b����KD�'l��婒��������a0k�:�;<CZj�����P����l���.�����9�@gW�t�B�RQ���%�����_v6�ԍ�I�[����K ^p9*g�c��1��~��ɂ���*|]�PMɑ1��X�������p�r�v��n)����Ҙߔ��F,�@[�����&%�Z������M�|C_��=-����/��cQEp/�� ���԰W�����w&�쒷�X{�C���D��Ɲ��Q��M�}~"QMg���Rك-ۗ����nKۛs��y0
ip��#˛PZ]��I�ڪR��8R�΅<&>�)��E���%2�5�W����R2\����2?<�Mբ�Wi��[��1�w&(_����n�/bZO'X��s`��з���sI�����r�@~t�X�l�W�	��yV������2��_�z8����=U��i`���9����:Fp�mU��j]�&ެ��0���h����z�� ;2���_�,.$����3 ���L������PoW�Ĉ=F�@9�����K<��	B��v?_��T�\pH� !?�b���b�J@���9}k/����O=c꾰�%��X���8�~Ec�J/�q�a��*��p��ܸ���m
e���eP�0����GK�T�x���U����h�XpQx��YZ���!ntt�^��я������í��8��0�1�>g��͘�*Z�`i��y�}�1��[�L�������kGQJ�X�����)r�u)K�G0K�ҙ�e?j�d���A�<,-�yc{��!F���	���Eu��������nI|�|i� U!E�\W�'�G�Ӑ\���k܌�!��"����嚖xɗ̌piLk�i�$�v�����d�dҟ�}-�AdQ˥���mM�c��x2�@X�� �DӌNQ:Eȯ�Pc?A��W M�k���*E��5�q�
��ÿA�"�������a�L�}ͧh�	Ng9	5��qX;�:gC3@��1diu8*���X@�].߷�y���V�oy��P��_�0�IΑ���а���%�dq���%�a�{�g�*�3N�ùy��}�H�ʻ>qe�Rb�1>�:%�(�=`I��l_DBlBG�0&�?��Tⓗ@y�up�H_Θ�]�e�yT"����\�/�� �-n����iZF�������r/
�s��4?5��~�v�u��
6M�-��� �T��c��D��Q�{��OeJ�c���6���zO�(���~A[��BHo�S�+�>v����3�8�U��/��>P%^4��qF)������Z���-��_��C0s��mR�pX�,k����/�+A��٣3=c轃�K���-+�$�� X�����]c�ۣ�P�B!��B��m"��(�U�0GEV	���W��n��'}��cd��Οכ`����v.�`5I;�#Ts���ï�[�#%o+U��7�1:(WF�M�����;s�J=P;!�w��v�������g���]�z������v��L��*r�$t�[� �<H��3w)H*���V� ܤ2|��H�E�xV:� ���@����"�3�}�V!��gr���H���U������,Zr��'m�T�G�J��	LX̠#�CD㈧�Sg��UD�<�d$2\�T�
��!5c.�U�ڈu��Q����\%�mǝU��@s-�y��I+����s^��LX���U�aգ�S�-�t�Z>�w0�d�|0�����,~����_	x���q�<9����CE�i/��H΀���֐�kd�lz<��4�b�E�9��{:�{���աGbB�����gCm�l���`�[�J�;��\t�Nv4�U4@�xlu���U׀]o���N.d~�󻟆"�d���َ_��SE��\�ԡ\R-��<"'#tlw6 Q���.mL�&��� ��؏V�n��t�΃S�y���W\�
г��:| �H{2�	�L�|��U�Η��Lg�y|VsB֮���+����)t|�U��5�L��A"X_4Qx�˫�k�Ђ�(�W���Z��a9y�Ӂ�L�[�T�7ڬZ||�+	��h�iXD��a@
k�x��㼕}E5GTU)9�z�f��Q���İ8m˸W6�⾨�X�ur��b���=LxkQ�E�Y�~�Ɖ5)���;��o���b�a��ة	���Ō�B�b>����s3�
�ըk�O+�� 7fW	��66�w���Zu��3$��}`u�^k�i;q1�q�BhԈ���g\�TK�����@	�r�y8�_ 8�����hCw�4T��o�2�2�-nD6=	Pu8Cqx6��������t�>��<|t�W���v�Z�#e�J�-�V��ֿ}쥕a�2;�*'B9tl�A,;�TX�	��׬�����r7.KT����
��ǌo�t��ʻ&��_Wo���/d@M�{�^A6�)l03� s�PuN����}Ǥ���V�Őe�l�=+(sl��9ϰ�U�\�H���<�!j���m�wPπf�o�,��	��?�pH��;�w������l�e�:���z�2�Rh�V�$�<�'ceY��=��YY2��8Aj��k�1��fgWY~icm�e*��;��VG���xW��X�[˖�IL����ð�ۤ!�qR��c2�p���A���*�&ՂIH��j� c#��2��Iu��b����NI!}0�J��� ������/c�+�"ڥ7jt�7���4���Q�j֏=���`������=��"�8U[T����*��A��M�ncX1�Z�J7v�΄�8̂)�QSۜ	�(v�����M��,匲Ǚý]��#�>����a�F@��4| �}�������ﬕ��'�^�<zڜC��16�TD񸙭�p������XĈ��S���X��]�xJ�">��/�8x�'k뙕o[�AI�:vU-�x�<�!ؓL}�W2�3�^t�%���F-��0h8���$�q�j�� ��2{	jN~�:((.pSF��{򒠒\'�|�T�Q]2�Mv�1�p5)_��o�G�_V^�� O� Rl��jpxsj��Ն�}��*ub	m+��{������6�)m���a���,�}1ʚ+�P� De�;1T5np%�_(����B�9�H�e�K�q��{�m�~� =�0j����lW���3���Gf�$
���,�Z?�^9|���G�;(�(x�c�PH��tXR�j���+R
j1�����o����--���kMP�k=����~�;�И�i�i��M�eVY2�0m�UG�1�3�j�k�$�ѝ�������)AA�4�
E�RJM�}����/�I8������ۯ?}c'�[v��b�7�9�����s�@�a_�	����,x���QL��o�H�O��Q�S���k�Y���f[�Lb�j�� ɚ�-���H�[L�G�v����N��+l����!V��(�[;Q�}7bI�B����	5P���7Y�"S��T+���<' 2��[�pmm�;X�L��K���HOc���o���0�P��~~͒���µ�y�^�|Ei�V2W��jH��wμP*A��\䷜k���O_�F�|����{h��C��s�p:]也�P���&�����N�xmC04�@���y�=Y)�;Ȗ�^ⷀO����51�d�몾F��ԥvdK�5��$5��G����=v�����Ō'u��d|߹E�2��b8<φl����l]�=�H �"�P�w��@tZ��a+I��"���i.�DX��/u����4~�t��������ir���'��� �'F�����&}�O~�02�j���20b�^����c�P�G�����	H�R�ŬZ���L`.EwQ���a^p/��T�u�H��&�,�8˘�GB�`�/����6(WY��|?�	�) �,�����[L�k�Ò2�Z��h���H��R��)] �C %���Gԇ� /���B�����C�6�<j�܆(�}�g�eAq����`�\�c����X}Y�Ou��~�}���9'3���	�i;�爇۠9��u�F�x���ɪ�CPs0�l����u�1m�