��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ��3͖j�Fgt��N�ZS7>�qg�W̾ñ���� ��Tv������o]|������XQ?�,ݫF��ɦ��C�b� ���3�ù� ��tT=�S���A nN�3�˿���XV�����8k�D�#G�4^\�<!ȁ���QeL]#t��|�s�A�Ū�~eř;��!�N�:2��л��z*��4�}���H�!Nӂ1b�qIm���D�=dq���N�������ޑrָU��ce0+�ݦ��+4���D�'������IG-e�[ò�-jצ�}����������:�����![���G3/�4�P�pj;XQ�,?�bW;�4}�+8�뗭�r�<+�TMjH�D��qg:ǻ�����팊� ����npђ�G��I_C�u��?^�S3�C��C��4~����}�Xo�>�]@�e=�Ѱ<'Ơ�h�O�A��Χ�x��`[\ַL�D�a�C�#��U�ypAj/g�^i `��A)��}�杝�ip�U}ە�_�I&(RM�8��F���X�)��m� ��r���H�>������d�0J��YJ����K8�Oh@��i���a������O�㽏TpË���iˈ����c�-���@�A�?lg�tPc��+WM��].���b���U(���B�lA����c�㏄��Y�N1�1�U/(s�UW��8����X��yW�p
<�ѹ0]�W(^
����� ��r��+_�_9*ɷ��Xm��E[��\$�����������r��˨��i�x�+����Ry��,yz)2��9�W�[�J��#"�/���~�(KF��m�rA6a$J�Xr_�~��fT�ݹ����Z2-_7���n�+tnzD.�7-�r��x!�v���,���|=����RH~����Q��'�w�n��X1�l}��v2:̀�M�E�6h�V/��2�6��0k����(���
���7�%G+�._�ry֛��|����2֔o�p�� �}� �4|�nkM��w0�S����^��/�@���E㶈��>�5D^�Hu��W;S#���3r}��GL�Q���Q6�e9�
M�֨DK�ɮ6�Mʿ0AgJJ�|q4���I�a~��C	��T�Y�d��8��E/�W��~q"�|zSp�t_U5,���#�yK���#�
��n��7����p��������d�g��K�7������p�Y}rq�9Ui`�%ւ��I3�*�_7�oc%푙��*:�ٗ=/��rt��c	�|�[�?���6ә!��l� �赨�D�b3�T*�ޘ�����S�W�-]�(D7'>bG���;]�ЖÛ�zaZ�Do*���m��ui9��w���p��Y�5f�	���4�qPSb�x������g�EET�kp~W���4'j!;�4@`�zB�H��;ͮ�[y9�΋U�բ���P�#��o��֥bL|�*Gp����q]k+ؾL�� �	v����"!��Q�g��%�^3�)�{d'.	Vƌ:*6�<=�b��B�v��$�C<��Rc	� =��Mo����k��*�
����N����r��&gJ�i
�ii�y�[��Q�w�>������q���5Q��d3����T�4�1]C����vjVl����C[��|N��6����H.��@��9T1R[4P�w�b��M��f�B���'�0nR<<������hݹ(�����C��^@w�h��A&���H��9�>�]�;gT��J�.gCyi���K3VB�:Z�fw�b����5��ͲjϿ��g�y�F1UW8�鰦�i�<�T/X��c��o��CGRA�"m�u
�%���7o�9�0"���
��0%T"q�9=�ivĺ�0d��X� �a����I�X��F]��V��r2L�r$��fRyV�uaS�CJę%d���Ꮕ̾��X�J
-�Tk�ql=�]��o�>���ڳ�3�48�skm�=\�!��䝾ݻ��q��9�[b�<ن�@p����o��j_\
2�
����¶�<0_a�{�x?�~�� C-����7��Aei�ه����>�"t ,.��q����`#�J>�gÆA	+6�K�����#�|���+�>��I�va��Kc�T!��`B�Tv'�!�@�_c)�+��W�jDE9T}��?ʛPPS�j���)m�oy���ph��c�ɶ6��i{r�$2m��A�\rË�����$U�J����?Z7�!px�J�L.�F7��^;��
D�k� �ʯy������$�ÿ��}�B2�G���l��T�UX�	V'�R[��/;�80�.3WM����p�6�oY�[61̠���8R-KW�-�;"A��p�w!by��Ĕ���C���R�Z6&O��$��х"�&�d����v6%�K*2���Sl�玡ۂ t�3錿�D�����jb)�����Յ"������!�<&O�E���KC^�!�b��� ��IRr�b�"��Sd�H&�-���u�U����R��Ԙn�����������ɵ������-�A]� t��]�7ڍԌ�Q���9_)�0oǧ�R���u\=�ay$R�$�6v�_JH��-��~8��,-�m��>�tE�
'����n)��I�����m;^�M��v;Fz�/1�eU��,B�Ծ�j����k���!�+�*Cj�$��_��s6�gD.e�	���N>e	�b�r�c�;���1�䷒53v���7����˷�G�9F�O&�_�l�K�5&3������ۙ�3"��h�����\��Ҏ� hY
��	9,�&ԩ�c����D���M�B��]q�3���������e�� >o�DEO{t�l9��*��O-��H&�2�Z%$qO��܃̬c~Qc�(xǂ#O7�#���M<}_͡��o���{������i��[��V���DS�b[��2^	�ҕi0A�����U���l��/(:(���r��D@j��O]1 ��&f6R�o�0uK���F!�"fQ��H�]��$ �X����~`Q�j��=��n<�y@�
b�W6�x%����6�3�# �+�R�hE2�$u�����������p�(��YĖ.&^���r�l����RL�:��{����ї�%tx`Z��.��J�8��Al���N����W͗O��������
�잞i�M�Y^c-�k��FZ��0���m�j/�X�z-J���x��J�>�<�	NdMCnj=�@ވ57�|��ٳZpS_���v៸���d�u��o�9��˖{<2�o^"��n��3�@�Φı�=ש<��J�����%a\z�Ӓ-�#^"T?o�;��1�/�@<�E�A�l�M��{�h3:�u�`&.����_��[�LI��x���>�:h�� s���=������� �׾	�Z=���H�1D�p��b���!C��?�[j���E�Ͷ�j�C'�F�o->h���2��F8PB*���I��@z�� �WIȃ���վDW+����dx��/�e�&ہW^ΓtvpqY�%�E��!�^�m�Vh*Kk%��*�x��<�Yt�?�����R�K2�\��Kj��'�Q򮐇u���%��2'5^\���C==.�A�DA���ɣ4��{ �K�9P�.��T����&�꾑s*��"c}_C��Ԅ�I�.Hmjٷuh�`\�l��7��c��el�g�څS�F�S��k�B��@�)��D��_Aquh�?���7!$q�5o2�6�r59�,r� e��si5���bH�t��A� ��m��S��t��f��9���_Ш��Gz��&�3�r;ۅ�f�e��������	�k�X���Ab�Y�Z���^F��	g��g��W }oZu� /4.���*��\��u(���@���D�2�}�P��x��\��@ȰȊ0�P54$3G�ĻU�N���$�9{�Z\R|�tt����W�Uo�=�����o�/G��{����J�����o+*~�}]E�����nG��he��3d�||3g7��Z��S�Z^�E��K!fV3_?<n�-yI��N8��4�{{�!�}�r�����ǒw<{Z��L�i�:"������zN�s�%�~������Q#=D�6SnMe�9%@�A�7�pS�A�:���?���6[֣��r��t���U�Q��o����S���RE�C!<]e�Iw���"�Nt�/���zIw$'��[�9u��}�Z�t�bE �tm��6��S�-�R���f�<�X�O�<�#ޯGj�P�!3�-%@�q�A�4
��,8��l5�@U�9d�)�:�v1��IV�m��'�%Bi������dϠ-d��4溪B���-d}6;.v��"�����{�jt�Ʉ%T�����(Un<�w�J�
CȒs���j2D�T��s�[FeT���D�:��D!�4;��b�F�,�oE,ʶ��)�����˦ ��#�.W��TO;��f���4꿢C��^�ː����������O��$��[;Λ.�*�H1>��n�8T�ꌈ�'9
*T;B����5�3N̝�K��-QAW�c@���
���:��"G��'Ӝ�ڀq�h�<)�8�����x}�W�����W,%�)�h�^��U̐ЧE�F ��
?����'!�^Z����hq�x:ȼլ�yȨt�|j�m�Y�uB�F����8L�[��)"C8�T�]/��K�TӅ���Q��a�L:�c��#�?�m�	�)�H��a�:����o��n����r˨5�aUܫ��Y�J˟���AC�#S�+��ݯ��=ҷ����X:|�t��W!+�<R&v�q�	���D�Et6�	�>��
۞CN�`D[�o9ɟ���}Y���8[ü���.�$�#�_YbG2�6�hH
a^��o�B�[B]�`�UBZB
��5��ԗ8+n߃�4��+Xj�TT�����mˤ|D7ʰD��a-�,A}yϘ�5���9�[x���c��ɡ�^��h�?�T�$�.4}��Aw�]1��@u�T����i�V��8�]��0px�D<c����{�p�<�7���r]2������ U!���=��n�ҍmMi??`Sp�WE�C�id�9�u��R�7�5aƿ���l-E�@��4��G�a$�2��M�Ō�^�\���:ȶV�D���<�[��m�]�s<��4�0]Pd-��L�LB��k�|�E8�l޷�V}�'�[.�����6���A��-�z$�@� *e62u��7�g�:���Ā��Y�V��~YF���ׂ0�������sU �����y���u��$��M���}��P4<�A����9I�[�kj��,^�v1K�J�$a2���F�R^#��Зx�_f83�	'M��.�|}2#O��p�x>�Ag9

G/������=�:XP�ļ�x�8sa��`0>���+Y�BSW�}A�s��-]�"޾��K{���d�S����	�{�`�"�pN����f��w���UE�4��\�ŧ�[5�[�=��c}���&�����y��XR��Q���,�D�� �t|$��}!��TY~��A�h��h���Ǽt�?��¼���>��'���)N���6vh�����
��AEg�(�B��m۽�=P!v�<��Ƃ�ko=J�z�Z��8fBҏ�";Y*��V	#/V-݆�	�9���E(����<���,���D��ȯ����Zf��3T��p��ƪ���ImR�%���=��嗂2E�U'�
3���x3_��	����1�FD���<���/���t���k*X�9�O�Â|�]jTe<&͹mrMs�9jC����x
Vx#YB��c��԰�������(��$饛FW6��R��|�ُ�BE�A鑛ɹ�	>V��ز���Z����w�m��r5�!b!ZZ+b��Q}]Z<���^�\F�ǁR���ǿ��I!�������gD�۵X�b�	W&&b4Em�Y�tX��W�;��V�a��Y�E��⤶���w8��J���:H͍R��\���|�ѫi����<g|ec_>�Oε���V�Z�a�-G�����f$�2���֔TWkPk(��������Ί�큷��� ;O�:�q���-a�q��6p�<lN�k_��?�I�<T��c��kq[`i�.y�I�] :���Jh�}�a��lg�Γj{6belX��\>�odr��i��5�ʝ}.W�>k)ٓn�D�I��c=�<�3�v�q�z��k;Ip�Ї��c�|;�w�x4�ڜ6��~��u��&��U�� w���L���c,��P~~�ՇP���*�mE$�
�*���9�?Ħ�?����)N��)�(-�~
O�J���Q��۠�5ŹU%Ejݦ�9��SE���J��:���F�g�>�At�x�t�u#dT̑<D�`����2aX�@_��l��'s� Z�O,3�0R�>���1a���S�
���ݸy�T�f���sÙ�]̚���������p��.Hj]���OQ:g(AX�4��� 7�͇<�m�����A}��F��-����P2���p�.a*�ƺy�9<���|�Q�5�����W�'�g��{��w�ttvt"td�L�m<��7�����XiN+\0hό�+-���8.�l�H�M�Cn�c�X%�sa'%����Y�9E5�ML�������w�j�G�_�	��7*vG#�t �怳>fY�UPL���&!��m4
L�ش;D��$��A� �� �7А��\b�c�,��_�y�T�K�6^� �EhU/�����V�k�GC��=���T܂aK���x�,��"$<j1,�K�74yR��[��x�0������, fy�_����Rт���h�6�{��F�~�"���&d^"���g�CڻJ����q�pq�*���Q�O�W�o�{a=|m�fFK�O:{����4�+u\㢛�)��hڕ,����]p�>��9�u�C1�|��@�ag� P�|U�#�g�eVmJ�{Viwn�r�d%� �8�u�/�tB\��,x�(���I0��Χ,wD;&�+�úI�c7.6u������M������;��o!L�M�-�K@{�j�bRvx��)ѭ<��[A�P�Q�%�R���|���M{D�P�g�ʕ�Y�(\�)�<�5X�u�a�Rw��/�ZR&H_�^A�%����r=�r��.���`�Â&�����v����t'<(鵓��c=@�+t��sHs��>���v�5��Y蓜h lF`� ���?&�e*��VV�VNc����h�;uڨ���:M����-��*vA;��Q2�d���g�)�'#d8d�6v���}¶�=>�H��*P-��<ݓ1�1"�І�9�$��0��S�dc�Բ!w�Tc``�����3ا�a`�0Y��)q�s76r8`��_�3�;����^췘��I28���Ь��~TxD�m��y��4c��ۼoɦ��c)��pK��蔒3vy�~��k�-Z������Ӓ�x��+�T���0Q"�d�ݝN���6�{J�<��v=?�t��n	���)�_6kFsK"�l����;���9!\D��	�a�@����h*0����,��֊|<�py1>	J���}��f-~&:���#�����[;�i�l���V��W�$����.f�����v�&�� t��j�e�w(�r8}�����t���:��J�XWX��F�+|��q�3��Zh�!�o�d���CE+#�}�zL�ErbVH�#=�[=�T�N�ld�+�=JC�&�>t+PA�+�Sܺ4�8�厭�0m�o� �x����mK�����%#5�4Ǡ4]ÇL���ȭK���A{/�-a`��������ɮO^��"�vӁ$T@x�7&4�y�p�E�	�'� k��Ε$�IW���:�r��L�%����k8$�t��P<�	<|�!7h��}�S��IvD��da��oW.ت��o{B",ϊ�M�!�F�}�ȁ*��pC�nIૂ����~[��
m�id�9,��C��6��1��)���/E�������2G1����E�sy�b�� &]-r�5i�2���B�jG�eVxG��	#'<"W_J�A:%��#!�a�L��=�P<*��z�w�����X�*�P��%+�7U��|��'@�҃
K���ဝ�����U�� W�7�"c�1��Q��d��(��������BI�X�ԚL��Ҍ�$�ԫ�hi��i���ބ=�6z��)�X���5����[�q�E�=��ݓ�H��3tV�_W�KG 8\1��t�9�� �ږ����K7�fߥ��<df�1��u�1�Q��vk�����C��h�E"{�q�B����T�loSk0�"W��7�6�>F����&}듺Y�9H9 �����`��'�y$�Ă����܀��J����H�A��SM� X�m���i
r�
���Li��:a�6��U���6to�ң��Xv{��<���x��`O�6�W�r��k��oc'ؑ�K���
F�Lڠ�ױ|~�Q����T��:�?�N]�2��u�3�w�̦;f؏�\O��'����. ��1���P1C@yڝ*n6��w|g�eC��ԻԿZ}tjk'��9>���>d�R���Fx>3�{�3�����;%^g=�vR�1���Y���[����)����6�!�f#��u_*����H��[�_�����?
��E-c�M���3��-{������5���y�5 :<���e��s������e�2�;����X�E&i�xךz�6\D���j�x������^6|%���:T\�2_�W~�,TU	qKH�>s:d �\��"���.�9����8*��>���=y��骉GM�3}���L��žW��\� �NN_��yB`u��]/�����sK[�gغ �iE��|�'�yp�X��(� �<,���x�r�ĊH�#�u���35Mq��ߍ`��;�,0A����(�p�V9�x�,Z�`�,�����Z���fo�2q��� ������oR�Fȱ>���~�����*zr�FO�Rp�P�	o2j$�#�ǜ�T����?:�Xa�Ü�~ߤ?������A~M˜��?yQ
c��B�k���NAR�^�BNJ��ÖUƪ:\���&.��Z��HA��z�"���)�+�C��e�8$����o���T�!�jI�;<�����}!J��U��ٕ#A����L� ��ԩ-��=�a���,J*��Lk��`��_]�"`\'�[Ϛ�ڃ<p'v�v�
�^^�^��g��d}��s��0�ݙEzJ�9�AJ��yK�4����%��~�+�	s�Q^'\����3�a
�T��5F�rd�kfJ�~� �.�~�����?�`��845M��l�fa�b-����@�}��B�7B>�:~ɴ�<f�9��2�1���T�o�%�X>G؈���3[�Q�3Oe#*4oN"���,�~�}J�����1oa�9ў���Y\����ނ��9��n_$��t�L9Zb�q�S����"�kܨRVRl��� �v`��1+����6�^&_|���.�����.&��k�]�et_�ݢ�O�g,�d�k�<�!Ի9�|>Ռ.Yv����Gy�#��(��v��^��Ћ��V�;�h��.�u
���y�yv��	��ɨ�Rb��X~�+�����ߠT���>ο ���W��<bI�X��f�2!���G"���2����-�T�����=ZHsltn�R�x��=����rL3[����hn��ӆWs��� ����G/��j�ֿ��q0�S�؄����ΌD�L�t,�ZxN_Dn�l�l���sͫ�
$`�۝gLgpL&9K�P-ŝ�a���<r�# ベ�z��yi�D�[�~
ø��@�'�da1���2����<�.�AS�y�:��8�X�W���%��O��m� 4uH|�{����H�C�/=
y��^Ԃ�d-�Jj4?HC{��Uś>�6��[abyGjW��ض��F,�k��:R_vB8u�B��eyy����g,+��4��U���n�=��uX���JO ��_�QՔ�D?��}G�5���H6��K%�#��RƸ�̅�J�R��+�G�Dx�%�L��B)��Hn����_,�m��ߩ�QF�2����������6*!�����Wa���
$�4+��tm���^��.�(�`�����A���؜�L�#�=�_Pj��n��B�F�-��9ձ���Ũ�Ԁ��r�f��䯎�u��ڮZ��0����8��%L5�pK�0~��p(������}�!�y�2#����|���v�P}���k����G�����9!�S=�8x]fq���q��z���f����ֱ��fh"�uM���:l���'�����������!!CY��^�D�����t��s%�T���T�v�(L�+ޔ㛒�25�u�7�����#Z�4W���@�xB4���xk�	t����Ŵ���"p�?6��j�c�L7�}R��-�<q��
�@�S�o~~�{�Q�z9oe[�umC�S&Uh���nJ�n��J���*(�&o�4j�k�4�}��v�3������9y	aͻ��%mu��9Oi�u�mB��.�çy�^[	Z"n� 0!O�0,Om�#���*��	+�lmޣ������n~Fܦ��^��S�[���$����nȚU:o=��A�"�{����G[�h��DM�?��ԆH<Fr��z[*���D���HϺ��U��9������������୏���$�8�+����Z�;�x�ph�o��T�{�Dy>p}[-�Ib̟�L٠Z
k��):��I�StY���}���l7g��)q�w�ȴC��C�s��m��-�9hR��Kǌރ�2��j4I�8�{����Fs���e x�o������=���W���8>��"k��P�L��p E�q��@/�^����ޥ�N�Sܑ�Oz���X0t�r�j��H%�#'(}�Rfx'�譊PR�=)ԥ��K�r*gsh����am�����E�i���r�$zCP��@�r!��q��MR�7N@��Кs�0�xL>�j���uQ%���3ɏJ]�d����xC9	S7w��w'��!쬚 Z�7Z�MS8�����l�/�آW�U<ᴚV��I�cx�����ο�%N}d�U��̳�� ,_�3%+�X8�V6���tC@�OC@�r��|X|�&��F_W��q��|S|w�U�2!�[^�e2z��Y�&"^�>Q$+�_Ѡ3K��Q�̕W�#P���cYU�E��)\וl��!��ݶ�\ߞh4��=��a�.�c�{���I�c�O������
%���ʜ=ǉ�1fֈq��t��򓋒�����;�W�K��m��ڇ�Z��-���|�9��JjӔp+f,�^<t��b�&�I}l*���O��L�z���9��J�G욼�ʭ���>ţ}��9�w؃ ��c�ᅺ7�0��0����R#�/M+��!L݁��+����^M����zm��5�>��Ҏ���@�#�5<'���Q��;�m���g?pz4-�3++pY��K ��H��f-�F����m!T Q.��F��&N=��Gʓ�B;>B.v��0��u���9Q r��?H�­47����ܪ�jvc�y3�.�IZ�t;�F�M\�p�s�&�lJ\p;dBXR�w��W�p:�ml��*f���˝zpe��0�QbM��GL,�IomKw��2)��^Ć�5���%��ӟ}��?׳m3�q2�<澡[���?��@}^�&��Fԗ]� �9��=X�Ծ �=( �(m;�ż�t,
�x����]���Ǟ�+���-�݆t�bP�CXneɈ��j��[VKF��"�$����N#u�O8����R��C�ƌ7�^����+D�%��҈��B@����o�e1-�oXl�; =}�!(����욈زthA���^�q�:+��*�t^4U����c��k�d�\l���r+GyJ�aT���p��#/���DӪJ�HI�����,�����0�ה\�0kk��'i>�s�)��Κ���(@48���`^���H K�b==�{|J��Lߙ�P����s�h&$g���JNs�!mP���2�$o}���O��oy��v�L�����x�[�M���dB��i5}�H���n�-T��.����j�9�4�[ɪ9p�qU�	��@�4�x���~�*�P�k����w��/DN�e��`�a(P)��Cao)8D�Q�d�էũA�E�?v�X��J�l�W#��_��p>�Ɯ�2Y#�m	[(��}EƮDO��L�C(�«�D�iWV4�"���M�g��S]4*����m�,w��b ��C�]��A.��T��,�Z�G�e#��1ޣk�O �� �Ԏ,��U��~	4 �w�E���ǭ''�J��T���`7�9��7��0;]��0��a5����[Uq�I:8Yܜ��-4�*���I���u���vV=79.�
ܹ�:k���]��&��R��`���=$��b�5����b��X;��.�h��w��
b��!�,]�t�uq3���E0u�^�U���FB��ý�/!� �Jf-^��(j���v�esjp?���vX_�jT��s��߆��dUg��~��i��!Y��o�k��9���%��h���@[F��s���}
\�C�ʅ����4�9�G�:��4Y�1�[U7m�t:	�?(W�5����GƆM!-��\�����0pjj;�/`�iP裧��^M����(��(}؉�ȳ�H�	��j��n��ܔ2�������;��I`&�y��@����W�1���;^66����D��6�6��-y���K������s'(�ۜb&���H��u�w@?��AYZ�H�$���B<o��$4Zfq�CJ���������Ȗ�2!��~���I�-��C�^�������jb���q䶶.){��fx�E����	���/�vqv3NqB��Z��%vV���J��w5\��Ʈ~�O�l$I��`pu��ȡ
�P�m�$U(����ᶯӂ͙��l�{�w�h4����s��'�.u��za4��=7bR�O(�@x�H�,���s�li>LX�h$�z������3�uL��ğ�;���*��Y6@C��O��H΄^�
�5�yU��6������~��!�knޏ�£+K�!�y��=}�U���V|�K��+*w�c`�$2�9�u����|�;�!��X�J�����X�oS}�������ݑ�bx�>����T˻%�閿�Uԥ�Io�S(L�G��ë�t[",X+���/�w���5@}q�,�/`��$��Y��S�f��}�fH]�u���3y֗��@=U��uV�0��y���U�'f6�u�(��Yi�O��Gnkf����@T!��`&�s�_�N��F<o��0��y�[�ߎ(AU'�Po4�`- �ࠒI���%~(7E�����p��,��z��7�6���|Q���r����Ogm����8�N�K���q�\�v/AB���'�iEb&���&�x��gAT܃=�����-
.���(�܃�P
�t\n��
*-��~��ea�{2^ ��ө��#�i�<R'@X���nr��� a��t�G�'�=�P�>�6v, �X��`�γw�@rT����^���窑q"�7(rtK��^e`��>�ב����������R�7UF�_$��Ux�|�6�f�#����rxf��p@�>`�)D����D!f�n�(@�>U)W��N4���-H�;Y��0p(z0�B�텞m�$ݴ�2䎊e(�������2*ұL�Y��3H8�z�G Ӎ���$�g5	�6YJ+:8H{mHx�<,�	�FW�w��9���p?m^����(]�W\��.��h�=��~g"n1r���3�S@�0�U�ɨYީ���V�ʽ=<T�������u?|YGxj�� у5�@58�>.�ά҃�,��XXr�ӭ[4ؗ�\����Aɴ'��>zV_ 
B0 �g͚�<�#琷�m�L���h��[��R���j=.���	������ϝ���[�Ȇ
ST�,Ho�tYڌ��u��3���LL����^^ d�A�=n��ms��z�ߛ�yJlώ�O�7b�"�T��$=:*��@��ݪ�Pb�����>N�b��U�ՓUͦ#8�P����=�0�����;L`{�Y��y�^L��x�#X@R�u0m��a��M.�C�bo�a�[��B�ʈ���0�%�f��
�|q������������wI�s��T!n!��.D���Z�N7�pd{yր��πhR��O³6��Tn��4'���z�:+ 9h#Z$6�!���z�pO��e{����oĊ����fҷР�9/8�>���EÔ_�9$͞K�_)]㶠X�Fc��j]�r)�J;��`45��>�OP`�0�k޴T�Y\��;g=
]���+CC��ʞ����`�G'D�DIk����	׎f��ܻC0u���K���]O��>Oޠ�v�K�>;�g�Ƹ�-;-�Z(��r�+dE��Z�S��}��U:H�<㑣ek�{l�Ŷx-�R@!E���oy�B�V�8�[2�L�zJ�� �	,dl���m9��B�XӺ[J1Lп����p���9�o(��
���y�i�O�KvUN�ͥ^t���+�q��t�d? �,Ah�cr~ "����{�|��zͻ�s��э5݆l�#��%Q�wg�p Nࡄ��K�]�H6�����«�&�����C�1�0`��Ժ]ڇ��yD!8��"�����V���G�rS��X��+lݥ�x�N� �Ӽ��)>�1'�8}���)�׿e�*��,be��b8yO���Oʡ꼢�vv`�3E�t�=��U����5C����cl��޹&#B6��9~(f��t�U�ʃX��@���B�����Y�����Ixԋ�r�� ��N-{]�X���܉�d<k�&��X.�ūY�f�Z��,y5�6<���-����X�%�����C���5bs�Nb���xS=~  �P@[5G���T%uf��,8�2묟
���k�x���ݾ>��ZK�#=�+� ���.p7�6PZ�%E��[6�\ZT�y���_ΣK�P��26o�{�(+M�R���:vA�~`�u�;�m�R�&��1� 8�vho��ŠǢ�+�r�$�\Z�a��}LP33�	y��(c:.��\�c#k�
a�|�} ����	��y����#��I��8�W���<��!K�չt��0}��9��"�d&q!dj:�P�Ä�;W���P�R�����#�8���E)���UE��^��Z���(����64_����!���ᇌ�k�@��w�,��$0��ߑ|W���M�K�+f_�
܇ؑda'3��,Nb��������I�K)˞�DF�F�{�s݀��	�E�2�v��r��UP=��a5���;�W9-z�r�'j����Z�Uk鎡F�%��*vV���S�#Æ��HA�C��d:�����C�f]����j�^F�b�����z�����<{��Z���!����V~�v�E������\U{��7��)�Ż�3�pх��U��<S��/�
Yױ���?O!�I��M9�<<e��|,��X��tE������M���Ӌ
���ڇ������0�3^�A@+�R���o�͹5-l������5N�����@��rf��)��	��`��~r_)�!O�����0��n��u�p��/��c
&�;�\�3�l�,g�eP�a�uKd#���d�1m��c��c���l��8/�����D��D���l�E����1�}��f���Ok���-��;�qVn�T��G�����cEJ2oj/��|�œ����B��օ�ľ���S?)�0��5:�&盱���ϭy 2����5���@����yg����b{S��'fFQ�'�#(�q4�����>6����V2nY<��$��-z�^6}���o���E��_���M*��kgl�ҋ�2,=� u;�N��A�pFq`���a`��[�$H"�:!
/W�d%��8���%�sZ�<X5љ���y��B�0� �$�L��A��	*x��ϗ�c�H)M��d���&�4��ϳ��E7����w>O���i2{V~�h�*�U"	7k��	Q-��Qcm/G]԰8S�kg-�"��HK���ū��g=~���L���w2�0G?��L��vk�BzErI�='e��b�yril�;a��%ڀÛGH8�o ���y9�Fl����^�&���F��=���l���,����b䎔޺��s�a�ND��֏~��n��"[��bv�(0Q�U��%�'�j�i���#�I��O��+8RȀ����R������G�a��[U��X��[�'(��1�?6��
w)g}D�XDU<��m��ۊ�l2��"�lu��Ä,6�E��+��)��$������-H�A{�}������-��D�[^���йv��j���U�[t���E��u�G1�v��R�JR���8���V���®�S�H1��VT�-ж��VI�(�N!L��O������G�������%Ď�ˠZ��E-���_��>���o��+H~���h�K�e�S�?%y�%�n�{��I;�B	����LPpo�BR�.��W���t>^�oG���2]�@��t��3�}�D��i%�&��e�x��;����q�܌٠����.U�w�Pė˼���,�`��G/�rd�i$�s�9�_�G��3�82U>�����	��1�)���t��0�����Y���D�!�!����x 2�E����4vd�,���̀ ����h^CD_� 6���� ShB��I'u������Ŝ�>�y�͛R3?^v�>�^C=�q23�Ӂ��D�p�JX]�Ɖ������Z� +���������[Ԗ��^����F%���$j�|��]?�j�uȸ��<���x������$���ˠ������r�Y�T��P5h����A����c��OacҢ�!�ѭ!�pF�[��	WL��K6[D�4XU�r�?`/d�:ީ�-�Hf���V�����mN�EӃe_x3ņ�d0��Aļ�l�i?l�=B\/�y]�؃��>2��mѸ��m�v� DxL�9�B�m����Y9E[���Q�����o���G�^B=sXW�T�k* fM�kx�\a[��`U�g����ѐg&��W���[ȹIi�sDW6
`�+�o�7�z�t��Ǎ��A�4b�K�P�:))�\��ʪj)���o�e���̪wݓ��h�Z�t��?$}tz�kJ_��(J�l�zV�NO�L���q ��\C� �h�!âGv�1K���Ii3���zB9My�)GցFd�I�J=���y��q�XŦT�3���W-o���d�~��"�%��{�ŏ��q�҄M⏶���a|X�����HI���/-L+p_�J##6Gs�8�|��ӿ�l�F&cki��@�':i�4J�'��=aJ瀴ۂaX��$�B��%U�� �~�;�~����5�g⏢���-M�U��g�-����ϼ�|m�r���#Fk�.Ζ�N�-&�*o��\gFmwU���N:7"/)��I�����v�R bP�G��H�$�����[�ϸ|�Y}(��kk�s&tM��X�0�,>u��p�&���ꡋ��J�1���!�[2P�[>�1~;�4A�F[�.�"%2�0-1n�3�i�lKNRen���!�%=�����c�t���.{y�Ky����S���3�-)Z�g�$t�bw�r�l��٥��'X�%�h���oG�łghmߊ4����k�5D_UY#n�8�"SP��ϯ��=]�`�����og�>�n��)�����y��/2�_g���k�Y�C[b��� �\�*~+ l�"��M�F0x���>�íL�5�6$�Z%���T$\�q�*c�j���\�Q��zJ���u����ɫLڶ<KW�$55{�3ց����%�J�I�м����$�J=s� f'�I��}�G�ͭ�۠�gv�[�{�b�-W1r���^̞���t�����v�f�a(���$TH��b[��Q13�u�F7��Cy��PK%4�N�3�0�D��,�׮�������02]�aR3�����QD��-Gچ��u��j�|{��k-�e�b��̛0H�Eu��[�$�]��ޜj%MC�� \מb��|3�Mחb䙄I�~h�'���ϸ����l`�-8�Aa8���⮧S���	���;���њ���ޠViP���W�xF��Q�qp0-��R�U8�K�������\�%aNqĚ'xG�|�J���ץ!���cs��ԡ���4g��E�h�~��u���S=kی��J�9֡`���k���U��>l_����u즱�l�PE�����LF��z�з�&�+$�c��-��f���r򰄪��n!$V�+P#�L�U�f�,1ZY�	��٪1ĬLks)s:��i�,�FE�x�4)hzS�RҸE��&}:�N��w&f��L��cԐ_RgR�U&��'ٛ�t��Y/�Z�%N�C��"PG(������3�^�M�N��`�;$gp��	#�����)��h�.���%�����?rj�	z<�bg	�l\�֩Y��6�*S���4e��8���4�;<�1�Nѭ��U���*���S��e�ʂ#E*6��J�ｍR�t#j;bԁf61-���u�4������]\d x���l]Q���ª�
˝��fC��ji���Z0��ܘB
�}O9�`o2>C_hX8nG�B�+��U?����X� h�;�|���| ~5a��BYp������FAU47֟�QN�M�^2}Y�%������x�_�זu�o\�w�?>>��ul՛����_�O��?�2��L�o��ӎ����ME��P�gj��)�8�A2�=��=4�zc̥}��:��w��߈��+M�3�9`-�F]�|�m��)�����ʡ6B����@�W���dR�a齀)݉ፙ�H��Ջx{g������8�^{���J�RJ��^8ͫAFu|;�[7��,�|�IP���
W���7��o	I��8��=Hym�J� � ���1����T6���IY,ϒ@�YCrC������Yܓ��І��i�L��ڵ8�`�A7h�ڥT�-�O#}�	�8S�Ft��Dgݶ�+��믎d>���H���t��ez�B4m�8�wɆ˖j�A�am�_�`����R.�˵�囅��m����"c�"�����0V+�)+鄚�F{ ��V������K�܆����A�&.\M�ǿj�16L��-i(\өx�Vsg�G��¡ې��G��3�����d���u����eFldDH����W��������(���~C�_��F�m�I����g�켫=�I|�
(�d��z���z����v�:I�' !+/�����n�U�P��}f����E���g��_���
�8�d�# k���K:h|���L<)�${�VN<�{���wl�p�=	(�f�.l%Ƣ��}�� ���z��M�Q�϶� �:
��:�\�ᜬ�\4�]Ч���z~���8p�ϵ���-$ɰ_뉎�l�Hֆ(J�,>l S6=-��$]>���][B�'`�d�E(��5��H��*"X���Ը�u�ٻ�S�
��oj��;��8��j�@��3x�Hm0�U�?)ޟ�*�9mi��p妊����W����lrMo�Q(����X����
����V�S�f�1�f�PTA�e��"3�~%��_p�"�a��Z�ĺl�O���p��čX\bM'S�S��(7Ĥ��C��Y��M��¢���.�XM�[�;�U�`�	}-���N�!{��j�r-�Wk��ɑ���Hz_ҫ�Y�"[�B�0��Y�Ҫ+��K?<���`�|z�I(�aW�Iݪ��PՑ`;g-����/�/^ć@���Ek#EG���2�%W4Nіb]!�s��"�j?iD����C��y�A�R ڌ14��Nz�z��$
�Xʱ�3*�Z�i�6P�	V����Hm�׋wJ[�z���"�=�-�)�{�}�a��7��ݮ0'o�R�RH��kj]܎wMퟌ�-�?Dmٳ{su\o��wN�͓��%,���s�����!h������NJL;�pz��ƥ m����i�r�]I����WB�j1QD|��~���p(�<k��
N4�U���; ���j꥜rc��HQ=�ㄋov��T��5i�J;N
��J�i�����nzG�:xLn��>U�ޭ���q^
h9�%ę���3؎GW��49r��ofL�K;���nw�n�HV��m�9��kK���;�	*7h�n͐S5��y�l�?��j0���J�T�.��|���y�ɭ����z2��c�&�i�
yRt]F�)���F�?���:�~@�b�h����S�����b�HΓ�vf"T��x����a�z{
Fn��4k�����a�Ќ��v b�UD₤�P��ܗxpձ1��[�rV�9�Ɇf(�����o*����*�F�i����yǌ����
���Bu��Q��OϬ"�Z��2`����ZVQ�m_�� N�@�x������Kʽw_�x����:��6m·�O}��.�hX�H<��YPj'�b"�>}��LZ�v���e�T�˄I�B����5Q�����\p[!����[ے�����;8��ʜ�(�Se��13 ��0�$�G�	��Y��f�f�qR���Ip�eHi`��/M�ś�Z3vAa����쪐=*C��
sڗ�c���D��u���q$u�aޗ���쩩�>����9/x�H�ee���;.�ٲkS�	c������f封�r�/�Z)�z��;q�wiwF/Z&h��v�1p=�Z#?8mg��=.����ME�����j�ʫ�}� `��{Xq]>�,hI��:JQ+@�9�@yش'��D��C
g��75��ED;��n�:Jن�@�;6��4.A����Hl~rz\B�|��f ��Xl8	�k�Cu�uS����bQ�?��"�d-��(WY:��	F���"����i��^IB�nh8����.��dMQ���;� ��Z�]��^��}b/��a3��.-�p�m��������u��U�x^@�R�L�G��U_0�X�͢4H�\�n���W�Âۛ��]iE�9�_�!Y��o_�0Vޢݫedwߑǈfr�����֋}�h����'(�=+��"g�k&:2ɐnh�pL�S}��,��gP�i���׺_p�Cw���]��<!H��r�������z:�}��̐�!M��?��h8�`��##rV�''�@�3<��v��>�W|-�2*�K��S�uqI&)o�+�ߖT����:��{f�A6#�j"Ƨ����e��]�3,!�QlD�����%�1�m��D�[�+��^l��� ��כ���4�gU�c�؏�A�Nc�F���͉�>�Ye�੒��o����>��`1��A_s�Rݔ[*��S��X�V�Ŕ���"v �b@���tD��-CX������%�]D����
�dul���٦e������%T*�vv]HkW,s����غ�a�@Q㕹���B���z~�P����������[F|?����M`�*��_6ސ��8�%Cr�BR��ţ/}��,�\>�hk)�o�%?g�O팇;��LM�O@ș�D�h�$��h]�ށ_ʪF����\4H��a+�=�ͧ��R�*gm�:3��V���[�������_E�m(	_+A�5ԅ(-��wj��������NA��k����b���eﭸ/w3��d�s]���Q�u�g����K{+ ?��S����9z�U���sg�q�b~��5�Ƣ^�(�9��S+��-�A�����PJ�-dI�%T�r�B�N_\�Yd�T�{����s>�8_����tt����M�	V�}}:!��X���Z�jE���0na�ǓC�#:��ɪ��K����q(K0PGiW���`}�wvEAtF�˦�H&���ڄZރ��~h�:Q������~h��"#�݌s�ܦPf������e��>n',�ێ$<٩mo�H�9�A��o��JG�BƖ����v���-�yLT����w��.%�G%_��,s��]VЌ[5R��g�H�J�QK�>�Z�h�hk�`0؀� ��&��.�dt5��]n��bJ����"�SM�Ӯ9�+��tY1\�f��7�����ٶe�H�/d5tb��chU;�*��*����1��4H�E%��B*y<J��G<hl-�![�dǳ6��(V���
��j��i���,@�� Y�j���Z��-�`�7t����$��v����ZM:2N �]I=��!l���m6T?�
��0��VDM�I)A��/�pC��?B�U.Ţu@�9���I�s©Pj�<�sh�
���� �ݓ�YP�5S�y���|q���D�}�ޝ��Rų�C�u���ӈϠ��1�p��?�+�זBqə9'y�����ا��]��7�#/J&>���H�h]q}��Z�q��c'w`e��W��k1M���Aw����R(H�h_:8�5��pƉU@���og��1����Ŧ�A��2�lg�M�d�6�/�p*����0��Z�Ekv5ރ&�ԜK�#�u����������l|J���r�0����KQyK���d��,Pp���/����4kQh� ��K>���e�s�x�m�L꒮F���6�������w��ĳN+į�N�v��]����2���5�~d���y5��\��Q6��������s@W�9.��1%X�����n~�b�̙{��p��l���
L�8�R���=V�0�;�n-x�Tx4��,�#���A��!곙Q`�$Ց�(U4$}��R�f"��l�\������G�/�a��Z0���Xq����6҇k�m-n��ڍt�����k$pL�|!sF��DPBg�CU����>�ȾMc��񎵫B��֔���A��L;�,/�_]Gx�k�h8:_ND�a�����x�~�w���Pӊg:oG*Vr1DP9�%թLU$��P�_^Po> 	���{r\��V
ܟ32�j���}}��@�XA�{�~;w�R�Πu;E�˪̽^��#�.�����:I��a�@А��M���}q��8�h�v�@�$ȰUő�,7e����W LP������|�ƫ�8�XH���*pNV����%�o���;�I=Sd	;{�[�%[,o����Gs��Ğ��~���X��l9���W]tj�S݃�e�1a[E[�v�2�H�����p�؋=��?ͪ�Aex���j����SO�
f�����������_Rܫ��["�S&&�r��[_ț�Q"�H���d�aܣډ����Y�� ��1�RX/ �`��)��o�|Q*�1a��m��Js���a����z��*4n�������䅋��s�BF���'�ξ���z�`�}�!%��
^Ho3�~���M�p�+�8�����˖e.�]�,m�`��@���.޳O:�DX�H���r|.#}���S8�{��`$�� �Fo�oD,�F6G{��+���HO��{�j[����{*RC�����п�~��PT�^O!ηf֗��Z�.���A�V	�L�}��?V����1�K)��c�{�A���9JSv��[N�sdg�45�T&t3D�$���ne��t�����ks9V�pm(�UӜ�I��]�t@�(n���w��(D�z�0�A��ЙA��v�RxDi1�*����ho������i?[���A��9��W�hЖV��i��s�ws�TO�(�iS �'�����i�p\�bi�^d�P���*��P��x���H���bL}:#�Ƚ��9xWnǢ��2'�z��������ADDH��@%d�=��	R�40�	����b�/��0�;�9�W�Tmo�� ������Ǡ2|��;�<aG�����g�`٪%�e�N70�KW��}�ʬ4$,A�H)��<�p��=晲X�y�P�|��Y�ڂL��y�*tѬ�|�fp�/P�1B�����x~vs���d��0ܝsp��NMr�����U ����X=���k���gb��L�Y��dsB`������J�4e���6'��&Te�܂�+��2�
_�a(S�
b�e�!��R�t(SӤ�:��Z�0"�ts����cB�Wș�`�u7F1�(U�z�4�7�q6+Pr�e`E����w1u��"K(���ԝ��ـO����o�%��ۣ��z�3�_Kh�=�8��qk+$����������o����lc
�~��:�e2�&�B$����4�Q����Ƒ�H?�*S��-�̼QPr�sr5瑵�9@	�g���,}!g���w���ZX����ӄ�=qΣ�����E����\|)���o���H�G�����_a�C CSwH�R>��苒�E������h_�G��A�^e?"j��y�P�k�v�:��Z%� �T.�8i|ά{�TO}+�1K�C��J�'�*�PT߰��{�YҘ�Eo9�cά�Z��E���@��c;iU��u�� ��:pb��=+���R~[y�k��鉶�Ȱ㚀����UF�"qs]��o��Z���ms�����ǔ�Dk��i���ȇ���O[��%���ʳO]M�����r���u$oF�,�ޒ����p�� �RV�r#����/� ���B��M��CYm���eލ��Fk08�yZ�A�.��o+�x�9[�C �C�x/>gi$_���k��C�/���[���F����&3�q����S`'�/d�w�o`��΄���F���	�E�U��#t�i����[!~��)!	�������) {ؐ�]�Q��z榯�|4�l,�F��]��X>�8��!�����¾�����&Ro�̦'w��\a�����l�]�u٬V�5�|ȫI1ז�%�²3ts6ȁ?k����0�ŗ�Ȑ�p�\ю���1|��'�6C�_,���H
@�S@2��Ka`��e� *��|�6=1^Ly��J�8���{�dn?v�duY��z��o�V��c䰃�D��W!���W��i��d�À%��CM���4�j1~�0պ�/Q$�{�0l.��j5�*�������dK�}���d�&H�nǸ�-#Ob�fF��?��ז����-�\c�H<�}�Y{%{�Cי� ���x�.8��N�JUpE���0U���l4��ۊ���h���=����d�C��Ws/�i�Uw�"�e�$��/+��R@h�U�A���Wd�^)��l�RP��m�?Z���$$1#u���B��[lXH��3{Z��((OꑾU��	y�q]���v�lJ���n1�8a��݀�����bQ�8�
�G�V�)L$�A��λ\
�y1�ߞE��'+��P�ZM���έzo��}�x�Ӟ�X�f�q@��r���$��Y^��'���l��(~":����S�R1�$�����v�0��dT�Éq�`Y�T���L���m����G)���q5���+RzVL�n+q�M�K+��ф�YӢ*,
/'�g��D�y��I��lC6�z7���5~#�5����Z�e�
U��I�L��gd<�1��
;�����mr�S��������.$�����i��
3�������=�"+�*��5͇�#$��4��$�l�b�]�'�T�&b-�NS�34�� B�X���P�>iwf
����VM������	"$��[C�d�k]8[6^��:&O��'��h�w�M�y>�u������D�/9����*����TƂ ���d(hz!�[�8��ip*m�?�.Ɗ8�e;?�t!�&�fD��KWH@l!E��y�*���{��-(�"��q�HϹ�e���%-�t}�`��jF�`� �95��O�z�)�2�ǎ؆��q.)�9�25H^u� DF0��?�7��,��N؁��޳$���[3�f�ւ�R�6�.ɎUP,y�����e�/@X������y&�e�FIcirb�nn}�g�x��^���W��=�/&����/���>�v)ͫ�-�c~�^Ɓ�nq}�qQ���8Јp
�۱�O�o ����бfEp�E�Kh��#��	���W�̒~�i���r�a1&��������4��뵱���w���舩� ���ӆ@��4Q���uɴ�V����l���&�� �:�Q_��ԡ5��{�7>_%2��hF)R�%bO�x�Vn����EG����9�V����T��`�Z�d�h�����ѥ��.�1q�n�w�K�j��TG&GN��]? բ���6�6B�5���� _7���r�����p�ҽ<ɍ���_��Y>e�A7�O$9P�{FT�E�P*<.�o�R��O�b����;�����T¾�pz�.�f1ri�,�Xq�>�� ���i^E>z{�"Gj���B�Iۗ�fL�W|Ϣ(�>8����u8yH�ӭ������d�bzW�|nՊ��o#wi�Ȱ�mEgq	�i�8O6���2��$���x*,�e��PW�A�Yb�/���fo�� F8�/)���>��� qk�n�R8G���ԛ�S���]u檸V�Tu|��S����R3P�/)�'8������Dv�wڱ��0��.��.�	D���bY*
c�����<0�k���چQ�(~����X��^�{ͧ�s��Z �2V������"t֡��m9�+jM?o�a�}:TO��`Ji�k�����'�u:9�s�?>'�5����Ċ��������x�l�J���7�K���ÓKc�o�(K���w�%��^z$��9�Ϯ,�p>3<d����>Оɭ0e�u�	:a%-��#S@�<i�&�PÛR��J�-�$ZP�E46����H��%�E =�}��F�G��d��(�9t����rް���浰��3l�F|��^Ch�D��{�~kU0�6H���� j�!{4�)ؠ��$��n�
W0����?��f�PZ���,Y�ao�|��#FS~|^"��ZN�'�l����ԊT��}���;��hIx���X�U�@��$�3ʡ�[J���pSiz;��t�p3��H7��G�.�cs��\C�*��\����,u�w�B$<��r�\	����>��L^V�ۣϡ5�����*��+<�X��kg�K����hb��/�ѓ�M�P�/����$��AV�4b�G[�}���;hF�0��ۡ�tj1��ۓ<��>��2u��"�eg��\\���� �CP�-�m���k��z�<��q�I��u=`yؾ�/�B�FaӪm�0�Qɕ�]ӗ�!/�d����b0��K�E�a��30�������tӊ�K'��K�"ĥ�$l)U�����vC�J������8bf��1ʖ]v{�_ϞA|�w�&0�����p�,ՈB��~l]M	b���'8�{��[J���a��V/�M�z6!	��;]�o$H.1��S�s���dI�b��&�<��wJ��b��Uō��E<�ζ����_ZQ�p"�T%$"�Nߗ)��Le�<ڢ�h@Bئ��� <ht��!ƭ��<[��L<�K޼����d�����j�Zf�_�,C۳��(�me�E���ڃ�ӳG�{�c�(Qu^�����y�t�R�v%�c%"�{�f�A�B �dvV��ϲ��ΊFt�dO�x+�S O�U%3�5䔯���'+i+�Ul:���7�k��/�<~[��^l�����ֵ�:�Oq.U�0��EI��el��L�&��Əř��ceO0��X�Qz���{<4�&*3�x�9�e�Z�?��+3�xLU�o��h��Ġ��_S��l�>�[ ��2��$P���i1�c޵E2.c�^WV�1�	��5�yN��2��}�����"����?���v�Kdܕ*����Ę.B��I�d�#_/lW	0�:
s��f
cA��k�mD���˂�w�( Tk�#�Ou����,�m͔m�O�z}�Pl�;qs
)_�\�E��3���E��=S�VY��E���Ril�������F��2w���e�\���Ɩ���x�?/�����W�S3��x�oH��o#���h�s	�p@5�u���]ԗz�W��j�� �c�����<�E�X7�� t���t�!ƌ����@tDGN��@-|�~���z6���F��[R���xb`����t��<xp����ޫ�����[S:�G���^I,�PoC�)ťl魙3%�WO��o�n����¹�aF�	Evi�m�Nr��ⷔ�U��4:N�����|<L܄k
���9��>��^?�#eC�T�}��Ud'���an�6y�~|К�Ɠ7����]��$��}�c/�0z5�S,��Z(!��#�+ߝS��r�!G���"Ofw.P}h=�
�����O�_��J��#��0��v���0@���$���0.w��_�"�%S�9�#E2�H�͵�s?�YT��a|�P�R��{��a2�^��%�G����?Xo�6�����7}Y�o�巄�r	�A�V�^���ɖOp�������Oݐs?b���e�O+~reɻ������X/�T��A|j`��8P׮����J�3� >$��qMꄛ�p�̒�
�#��M;���(�O죛֠��mS����5tq�j,P��W�yIש�(�%[����9.�7@q(rdI�``�+K���|�����1.����tL������Q�]B����+Ԙ�s��ܔ�4����p��
�K�!2{��~����^a��(�޴n��Q�֧���������� d�Vtк�
H�>��Y�;����w��-�ʔ�r�b��:��;v�)W?R&��*�4x9�R�r(�8�����l!�r-r�����Qv�Ѣ��;�l��E�
m'�)� >�����~�S�DC��ư|�:�����	�}��M�ϋ	��^���*ɝ�FaL�8�鿠G�ؤ�%؏�Lom�*�}� psl�G	k*<>w���!�$aɔc�X�SZ�F��<V_�F��ƾ���7ǉ�N���m�>s~�ۉ�Z"/Y�P_+����]�FK{�����n?��_3�-�e�� 'T*:{t�ͩ�ְ1$Zz��7�Qj�ū��-��+�=y�m�쏆BD6��V��fK�.)�F�2"��)SK���JR9���T�炎�XҌ-����z^fD2����x�Hn�2���e9� �.�����P��ֈ��rǢ,�����VU��BPLg��9�K�T������� ��΢�OE���Ol���T��o�uS,�xU_b�2xA��r�cj��P�4��c��~�d+
��O�\4�����ݫt�"����R�u'�K>� �G�@�����fG�f̎i��,������j/]Q�r|M(�sːQ���,&�qkJ��m���F���	3²�6�-2�q��rՋ;z�a���6�f"�6�]���^Ԩ*��� �7�`"2?�h�T���6u���?��WB ���}�@I����S��R��8�s�-�U����V��]��G���"�V׿rSN��q��g�_p)-E���wt[��)+h��4p��ր^WQ�^j�rLXc����Vޝ]lG��������c���H黛����M7�igR=���T��9���V1F;ms����~���؃;�3�Բ�zj�*��FѰ��iRq^��hs����=���%�U�C�T���|�:e����9�N����R/8�"�p���wś٤t�����*�2�\�O՚[��"��ϊW��N�ݬ�9Z��jw��#�$jK�s��H�ol	g="|<�=���Ȇ��Ӫa�-��eG>��V��'��yϫ/���@c^S1tR滛�)�/m�B������7x�YF�c�AU��p�f[���8.������c�?�i�MxpL@�
\����׆�m�t_��n_��	mj�$���aӠ��hi����}@ֹ��=6���pU<kq��_8�����1z��D������!���5�[����.=��R�2�ͧ	Kl���a��8P	��/xml�f��>���OP�x��1"�T�ĥ��,���)ϲ{2�2iA�D ��;���r����W����6͞��x��1�q"�=�Aw����iu�juI�!�y<�=Fx��lǥZ���Z�tIN��v�Rf����.S,dj�Hq|,�S��_r�Tbm�.t�G��	�Q��x}B�˖�8�x1�r�iJJ{}h���6��6
��ׅb X@�(��A��m��֍J�����:�.�2�{TL���d={)��=����S`Ș��X!�<�᧽y=�Q�G�9��*�d�8�����E�7�j�ׇ��˰��Ut�b�O������N�i��/Y����*`���k��1��PF��L~�ve�I[�Fa��������	{�&T�[�lx�YL�4F���o���lJ��[mL�&��:������5��������6֛Rݣ	A��(�ڟ
&��Y�x��oKI�FXlZ�K��2�q�P�Ai����b��vZ�l$G���:�]!>���1��/$JN��:rB�ḟ��/$�6J�F���>|mM��/�xi��[��*Wҍ�M��˂.>4���8��kA��e$!!��Ô�SG+���r�_M� ���K�B��K��y���&Ac�M.U'zO�����B��>,��5��P�����g��bj"I.�霈J����F�w�����I�r����A�AO �"`ï�,����|eL���k��Ÿ�o��3���
!A <�ąx�� �ɳ#�.!%f0>dj-3[o��'�I�=(3 �@�U�P��n�q�����o��50Rٕn�����l_<�,և�O��cX� k�-�!AŬ�:=���$oܹ$��7u�\�U�b�Z#����w9���<}���K�/L�����o������"
1�MhF2z|d�xg��bk�b»�~��i��T��
�kI���ɷ����=�A��^s[�su��)1�)	�1�l�Q"z���t/��`k�qP��:6�����D��w�A2�v �d��z����pw���P>?P6��ic�Hj&������S?'6~j�b�ñ0�� ƿ����:7&�Ω*g�W��H�)Y+�T���YP�!#� ucpMx���I��E����"L�=����]��G�?�?w�Ѧb�ō�/S�J?��\�u6i5E��Y���U*��.4�AZr�Rڌ��l��W&��E�ҚD}yiT���a��2&�Ǖe�VvG:[u#en`��ߴ�D:StJiS���o*p0����g)B"_Z��wN��f�ڣ�0vҗ��H��M����|0GHb�8e�@�`��e��'�Lh�NrT�$���)I�5�B��U�ɩd���0t��zq b=;�8��?��h�����mbu:v��DC�@Z?%�Z}���m^��Q!�g>�:�`��h��0�Ƃ��MH��ʐ�O`!�`�V��g/A��ؚ��]��i���"4�j�y������>:���&<v���&�r�t��'�Z~� \�eY����>�Q&?,�����H *�ڑX~��5���*�$��	�@Dbbx�(����۝����%LկJ�qΞs>"��H6�F(�E���7K��}k���]0c^'��1�� tY��ի��
a���2!���LL��"5Ntؽ)��� s��+5�4.g�[�Ѽ`��W�~��E�z�R��ѡ�?�l��$���c�af��~n��I\y)G����ڙ��\<:��yzs6V�o�ôIx�6�J����w!�f}�H��h�����z�R�2���`���.�'��/����U�I�D[����G�L�n��ֺ����L]z�؞�W1�%�t�o�I�j'k4�nt�c���J�D�j��An't}2�tmӼ���^�n�2Z�@�h�����b�� )B��0Ƙ� s�ٰA�og������F%:.ta����U�`T�����Zn��rwR����ޜ[j�K��r<��:_MVL�J�,|���7�|�~HC#�S��*w\=i�'e?�(d7�����41����1�
v>�z~��>S=QY��3���>�u��nȱ�5��
y%t}(����@�#����P��(�}\�y( ��M��P��U��a�sҗ"�.���n�5�b|�(�֍NkD���N�̊|����Jҍ������Ū>~����@8�b-�����0X�/���ho{��;q��fT�W%��ͼ� קQ�����M�'��!"�c�h�����P,�8�^��DH_ �N��)1��Ƭ���o��������I4 Q��A�� �q��u���J���ޠ^}���3Ib�H]i�����T\J�W�!�pD����bm��Mv"\�YĜH<6��[OIҍQ���Sn�~�%�_�)}��!B���P�a���䱸Н�Q�7����F��Re/n�D�_�mL^�f6��Z�D����f��>�;JH��]�N3��(`z��|��I~���B��)r�$aM�@����`�ʾ���ȦEY2�6l�#��Ɓ�F��X	��������2ҥE�������
��R���p��P��u��u���FM�!#�&b<k�2���Tn�y����-S��F�4��B\օ�Q��.��):~S���ko��4T'�,^�{?��NW�����k�>��6��#��30M��#Jx�u�i�
y�SUΏ.\g�H+�@3���>��U��t�"TR2D�\����k;=}w Xr��¢qab���/o&W*�4a��'���y�(��jq�l�Y�D�q�0��Z�Q9�3_��[i��Lf�����3U�m�_VL�,
o��A)��Ie�3�"VL�X�O��d�y?�"ɫ_xkj�</Fw�F��U���^o|��K�z���Q�d��oi��QP!*�c�T2�+T�&+�������� ������K���KEM���Y�m�+�8/��+��t�UQ)|���T��)ԫ�c'y������8+�k��1K�"��=��dO�<�od7:�F�d�*�{��'�D�4=\�!*y��իtN1S��x}Af��37���2B�8���\Oۅ��E���J [(�eF�W7G�ή&�m�5)	���({>t�1���	0�ݜl&(���d���B���J�|.J���=��X�H�^�X�L�b:�xOı 1UE葋Z���s�
S��N]wyx�\w:3��۹�r}ޝR�ePn�CN���E	^�*X���*ح��2lm$�$y�y����B�N,1�ǹ'XqX���HPv�uI���ƼK�U��6H��5�2@ a	��CG����[�P��{�%�;�S���|����|�1��:>���ׯn_ТſH�;�td;��prh\i%��
��s�ሴ��ቺ�B�1>��∌�S��V3L}zc�k�ʒ@���7�yC3�Y����T6���_p����Гm�

���k��ͫ�v�bR�틝��;$�y%�|L����b����b������_4����Ǭ����x(|\���6�T'�	ynM'w�&��J��L;��{h�w�W��C/P�ؙ�/�ty|�`�E3i�ݚ%З�B��M�>r�Y��<�xQ�z��I�o�ã�����֡��s���;l�Y�ߗ�RQ��D�������;�CR��Ya���W�l�v��M�D������d�J���SR�{��M���
���"g�w�nk��!d�Fwmŝ�Y\�: ��֮w.�a��	�*SV���/�(��������_�h� �U
p�,�;`1�l3GG��*	C��kn�b �6�L,�eψ��2���h�l rh짫8� cOӴ����W�>CTZa�����\��eV�%�I��%��cNA��~܊�m�������z�hBHFϟ^qAB�F%F�z�'G�ܒ����?O*�ٖ� �c�|�'�aX�8Y��)/τ⯹�CF/�4Qe�f[ ���-��(���W��B�U��k��(�M��pk2cM��([3�����K��?Б��]����`8}P�e�Aq�m@��D��p�v�Tk��{�&��Ƨ�m���M������l��k$Y��Z}^>�R���H��w!S`$�	�d�dƹ������O�(���e.��r����I���.9��Q�ӍJzJ���u?��7����h&�������gI���
�M�1!>TM � (�]h�.`��Z���ه�o@�X���~u�8����[R�6.X�!�ji�������KDe�O�0���)悐y����� =4������c�di�bDaGAd�h�r��_�l�+rs�����M�Z��������_��(2��Y��<o�{;����!�9.��9��/�Y��D�=�0�h�z�_����z��h�2_U��0�I�z�m�>��G��jkK��)�2S`_l�ZN]W�>�O93M��*1�4ͭf�DY��O�Ym��J�NJ�%��fMo�J���)�E]P@���^99`�9O�����4?C��հ��'3�U��(1͘����=��Dt ���l���1�'Z�|C>_*�Dm�{�.+`��`��Y���iU ��f8�d���{W�u��H�ZO�A��:��e�8�ƾ,��J�_
���f��W`��{d��(��4gg� ���a��,�G��
����S��d
T,���i|%�tv����T}�fk2]^�X(<����qTs����	N�|Զ�����
�f_;�T�B���i#t�G�&d�?��M_-�02&S_��_.��8����K�Qk�/,����GF�]l[�3����,���g�&�}���h,�(���;	�ٿ��ӿ������z_?֊�����`e��τZ�$�ѮDIi,�.�N�[��ϭ�
�D�.�酪;�\Q��C�Z��E�'�e[(�`<G�)��03i��ScX���qoR3g�Vݘ?]����`i��_C�;#֪�+�*���u��X�����"S=�ڞahX*r�Y-�^��9� n��P��-R	����L�W`���{0~�f?��A�s?��-�C��'0�G9�{e���ځ���=^�)4܃�B�n�ӯr�*�����M�j�v��k����l��/���h�'��cE0v���,�l:E�͢�]6u�eįq�d��p�������Z�'�o�pxF�$�����c�s�n��:ex�o0�*^,�� -,l��7��݊�:rE	�ޥ�Z�0�z}���G���-\fC��j��`M�p����C��( �1D�z�����l�L����$�ƨꩆcph���Y:�ZO�����W;��J��O��a�L@n���1_�T�Օ��&?s4ӳV��t�g��\s׊�4B1�>r5!溄���=[�^0jڸ�%��/iȚ�F6dD���_��ùh`��呐� Y�MK�Ây]S7������Sc��5��n�H��2��Pn��ߤ���k�>�8����<n�'c�;�}��6'�|רQ$�)�bT���xk�F\��������S��69��ٶ�z�w���� ������/�
G�zT%;~���x��n=�#�������8q(���N����$��E�?V����? 1�<��~�F�3���E��[�/~��w�V]�M�B �x[Ga|���~��kz�1N�X�A�Ii���_߈H�
�w�Z�~�tQ��&�n�(Pe�i&��h�U~NNG�2��}���Q��Rĩ�hZ:�2V��?){��e�������pu��X3�l�f�m!^��]���M��2Ɇ�݋p����`)K9�4�:4�
��zD&U�E�i������wW���u�#�y>����G�������o�K��^xF]'�l'-�j�|s8ފ��vF��%��C�EYܖ�E��x�y�C�7��	h�M6-S!Q��6S�@�5��3�:��k8GT�M�'�"�L0��;h4���@�%����[��G���,���X�jYbl3ZI�wP�!-EH�I+��>��gP��w0�o[ϬvK��1Of�$%=Y�~=��a���9� F}TT`�Fa�`ħ��T�bm5��|���6�����gP��i ��:�m�d�"�z9��d0�נ�+���"rNT4�B��`6:�M3�,�X�L�&u���ag��c���@a�˯n�yZ����U*r7���~���I����.���cG;����P�+���p�p�e����9�S��@Mi��c���B���}����̅ve˱f���ۂ����E��j��l7*7���Z�洁A���w��&���xxK���\6B���[S����I;��3��OQQ/�:��%@��{��BJDߘm���ٙ$���#T���%�#
 ���A�ЩE��u��E�_(8�#����#��k�]8���gPM��r$X㙟rf�s�y����M��E��؂�T�9�hql[{��a�ÕR���xA��k�b9�[�Ǿ¸j��=�����,{|abM���M��iy���QQ����J��&	aE#8�t�:��J��9�(��X�Js��٣M{�<#%R��Rd��@�"/�B>�[OS�*;LUT�Hr�	8���[=E)��P���"�Vn�˰�6�-H^�	���__l`V��Q��j��x�b�.yVl|��@�O�۞�sP���r���%~_�9�=���ht;��w�Rr�p5��g]w�M�`���[��
�yV{7;�[�<c,Qɓ9�3�Cl�d,�P\��-�И�Oo�)��;�lFc,�յ=o�y����ļEy~�<�c��B܈O��q�/�K�R��_��[�q��a��Y����!�y����c���x0��[�:��b�R���t)���SS�3Ec�є-Kݛ����v�'q�M�j)��!��2|
B��,2���ɺ��Ds6�͜��yi��.x&'�p�f��k�c�,�-Ѽ�_v�����{)���L��F+v��xx����\N�i�U�JIYO�E�G���ᬪ�����t�겨�}D��Ӡp��k�/��zhkYtkO�x���]o2�b��3O�̜&Y_�ec�?y̠u���p�MJ��Q"��1�3XyΥ�:XS�ǭGȜ�\�Z>��f�ϧ�ί��-n�b Z�޿#<  {�t�A3a���'5��� ���=���\SY��0n��*���`if���������f�V��&�եZxw���r�eڈ�;�llwz:ҒR�k�3�"5��q��[u���������he^�CRU��w�#pε���b0t}Ur:K��!r�����/���E'Aq�lfkY�ve�P�˽2���Z��
�j�4i�p�;6C��>�O/��A�����_�k�Ѕ_p��&=�ҳV-yZ�)�k*U+ߗw-
*�����఑cȞә�v�a��-m���?�it���	l��|V��`,rB���ʇu��N��%+2�a�TJ�+����\~�|V@�%dt� �x��!F�
9+r��߰�y������`=�����x�����H=.��c/�0��gڏ�HU���A"&^��z�/U��~j�������^�����L�P_/&:����������{B�Hr�v�C���� ���sK���"/x�\O��k�F���5τ4	BM��WN�����"8.���BE���/o;ڕ09\|:�y5��>�t�2�M���.~�>�E ��h�]{���4E1E�쌒�������w��Z(�8����~Z�g
��[�5��`����{
���C��+����N)�-b�ń���]~c��:MM�C32�"^�4�#)��_{��c����L����W�D�����?����DD���0n����F}���$�o}cI����ia�x)H6��6�^�������Y"��m�tU@<nJU`P����3V�="#⚲���̾�3E��l�:M�nb����	w�>��P�
��"�p�d���S^�ak��$D���"���P{׼|��61*��J����LXk�ĭ��UR��%�_�Y\����|y��m�Mξ������k?$���Ep�#wk����1����836Q�I�&գEh���u��t�8R~��R�^�)�o)V�')�֓����l�MLyDB�$"cl38vJ�Q�ɾ��E���ye�.�Z�Li��1���OL[�%(��C(Xtm�����%͓��T����~8b��R3-{�B�Z�7h�~��eڕ��$}Y��z�TF�������x�ކ!��>	c�}���clR@J«(�r�ܯ��K�k:`(��=�Z�:&�/������y���L��C=o�u��'/c� �U�w3�H��6>6э�yl�mKh���bBP���Q��+2ѫ�2�?��ÏFZ���ϝ���	�_�Կ�iMsz�'�k}���ȓO;�""������'E	���8��S]�6Y�0����<�M�p<���nG�;����S��ۖ,�̓��d�3;tW�z�xʽ�FB���f%nCf<a� ]�DI*�.)�G�+Y���[oB�G-f ���.W�X��lQ-ECt��$ԭx�w��Y���-`������CĢ܎d ��.w�!��������C���a-�>��8��6����+�.>�H�
kt�'�OX?3_��{S
&=5�8T�;�������#ЌhD�9�v��o�J��
���.$��s0>9���(��^�h��.	�`�3!SR1�{3^Ԅ��밺=*�1�Qb&����$��l\͒��o��9�􄯛�,��ҹ�s����4Z��T�Wl~���ŝ��Y�� ���J��5)M�T�2��&5�#I�4ZÚ���ۄ1�jJQĸV�u�wMJ�lY7h�⾐n2Q}Hg'ӵ��/ �[���X�*a#`#i<�k������$;�1J<v�5CEEP���5��s:�0��qq�I}%�������^�_�T�hHE�ǘ�9�`��F�K�ȓ���\7k([���ȟq2���Tg*]WW����>���,����Ø��.�p���C'���w����lS_�7�n�Ud�r��N�j;�ٻl�m` ��e�3�-q6<��3b�H-��>��[��xu�٬����U��`|��)������2F�$6e���x���NhB�>*�bXO�!f��<S!:�Zrl3�Z������Q�d�VMnv����H��@1t+?���s>n$��>sh�*�N���p@Q���{)/vL�LGhv�-<G���ͳ<�Y��)��$�v�^D�J���x��x��A��K�/��<�(�����l6����7�@��*{�Җ�;�rш�lC5���=8!��������w�0F����n�cnV�tG����W�(S�\cL]��b�� o�?G�`P���G>����w�<Z�˔M�x��{�_M�䳏��J�,�3~�?�k]:�N
��Y��j���w��d=�4����h_������/� -c�-<q#eonH��
4ov��ua��A�F����=���O�	vcG�Zɹ_�gn�ķ�n���X����V�6JQ��V��,g6\��B����X@�)�7f���k��+MԿx�)[ox�F�+w�inC�����-m���	�o��7�w��v�qez�~L��Nk[+�5�ٝx������JȘ��V(\'��XOucEbV���|����Ϡm#_�hf�a��~��LQ,�g�K V2׽n���f��)E�v�	u �al~-��aǺ���i����a��j<���Y9ɧ� ��m���.�^�l�w�e�_�f��
��&���8NX�`�����i"�"Wр�%j�_Ⱦ�]�=؇Ĺ#�Go��}�8ܞ��[��g$e鈞5�G�������bW�%o�r�(rp+ێ�[��L
�E ��F���6��#�����h��ױx��f��Y�T�Z�~C?�j�r|�J؆���~�@}P�d���EgV?��$fFe�n��]�#���И�P�Q:������m�yI뮕,��s�Ԫ�oQ�R�����y7�J�v�����h��E�"�Y�6>x�}�I5P�L�ڟF�q�&�=�I���7��bJ� NoF�4��ljΊ.2M�*z�aIiSu�nSB�
��}�Is}��z��������ZB�y|���Ն���A�~�e��|�B���P54��� �1��&��V�_#������I 6���h�oT���޻�	cO�mcG�~�A��BE���9.u�UrX�$����1!��$cSm.��?'|��K�<���he�������Ճ^F��{��r�?xO��|�<򸤟O[��2��W&r�!%sd���zo֭�U�[�o��[P��c���n���%�Y�P���P@��<7N��1P��k��M΍��!�
{��@23*���X�3Җ�!����c|�X5fS��F�����=�(��)I��,8��.H����p��IQ���.��-�IY��|�ψb���,��A�1�E>?���E�+	����Uoܹ����bb�?Q�2-e<D'����ù�3a��R���y"���Pp�	�Mo��M�8l?�0�
���qBk�))�dY�MB�;>�6�����2z𱚤�� �3-P@0�	肂4�Ƽ��T�M*�O~�����������!?є ;aQdW���=�yDģ!Ѿ����>���8�/q/I(�/h���)�l���dgR�`�Ys�4�d:9W�]oAO|:Pk�5pYy]�ag&����f�v�~��tn�ʝTf]Dվ*Ǭv2�
�����2���`T�Z9��^�+��^��7hHށG��ש_��&��#�T��:{�Z�]]��X��l[T`-���&�E�h7����:�b��;Qh�~`7���mf,Y�1�T@K$w�9��@���"PS��kN�r��Y��)�]��%���[+Rg� &'N�x�'������T�`t)�0k��;c�]M��k:fE�t��0�^��ʥ������ABB�ĺ�|N�|�=a�A~ms}a�S��f���h&VZ��k-�a��8�:Y��s3��i(���d���L�o�������x+ � �W��Q*��1fĻ���~�~t��=q
�V*���ҿ���fCh⮱Z����u����e�2Y���jWa���@�'�_)M%�ҘO��V��;��E�g�W(�0�����mM��ji���$�aH̏x���+h'ŋ�"��l����t9��._V��^����0TB�)d���qY�P����ѹ�Ӯu;-*����
}zZ��l��f�h
�~�>-B�	����35K��ê�Xw�����΋�G����ԓ:�jǶ��L�p���܋�L�I���e�O���Po�<�TI�Hg�;�Ò�R�bۖdk�*
���-e���0-1�g�k#�r��L=�,>'?�/t�Z{�+i�j����r���S>��!D���]�ҙ���]�8�^'�˞Dh�m��������u����ؗ���㐔��_��\U��3�뫕o�1�ڿ��-����T
8������x*1�a/=�B$�Ҭ�L�b�w4����Q)ő*G
P;R���G��aD�=��(�!��Э�P�]M���w>Mi;�g�&�E!���4t�G�
�[rIܴ�L*ORӟK^vX�s!�n?���4��g��HD�/w|U�N�P~�����}\d8�*��p�����~�|����ٱ�r�
k���C�n�U�$��5��+��d���Xv�������E
��r��WZs�0�'���1NL���H�Vtl)sy�dh٤��%���  y�1�(���W�q�[$���Pg�������hB)	�J��o��O+�cF����Eu�.4\ʨX�Ը!w>������������O�J�Ⱦ�	�?X��4Ԭ��6�Q�$��H��� GX��&R&'��7��2�+ږʳ�_���[uu_A��ط����k|�lD��}�zڝ%N��#)���/:.x����$������N~Ŗ��2?�(�Qv�e1��5�%��|2~bdz3wU0d){�bi.���6��9hg�qs�R�&[���FJ�9�"��w�ǆE�{݈e��v@����Z�'dEC ���o�����P�-�߈`�?�a�=#�+�B�&_A���� :.�|Կ-Ͷ��S��t�h�'/���8$��ك������TK=yҧ*���;]�jm�����Z������Aw�W����D���2K'�N�9���l6#��T��_���A�8��ռ9ovNa��}�F u�9i�A�H��,����I�C�ƾ��o;�h^o���)����=�֤�Q�*-�;=��q��Z��8�YY#9IS��aH���y5'a+y�;�w��qj;s��&~-��^���n�U?���.߯�m :a<p����u=�9�7�a�� .����<�6r(UZ-����>U�yJ@�#tM�E��]]���Pu�y-�/˂J�׋��8��:���e��T�36��i�G��C��
c	��U�b����k����2P������T��IgN��ܶW�)�\���\P��Dת7��iЕM�t�0<V�Zg����穬e�������_(��'.��N���8�~@�54����Eg�;P�~$�mD�NoQ<�m�떟�t��è���i��@��m��0jp���ͦHd�6�XlĲ��Z���G�?.؅�S�w����n`WA����GŢk���H��Q5"$�#�@ >J\�����42	�Z�����FgF����fC�:�iPo�q2"^�ޖ�$��L��Hmb��#/~���v�	�Y�{�lʗ���Ϟ ��%E]@D��H)=����(���`S����
xmm�!`��7�׆HH�3��l=��,�1P�U�ģE�(p$�6�ntQz+V�C���~���q!Px%���P��մ��?���D�z^��O�L
�-����JM���X9E쌉���}�d��%V�dym.f-�/rAĵ�}�,��"僾
9}V��|�~/��8=����f+����:�mL��f�]��)]�o��?ybn���l����@J�����.3I'm�F�aR�m�R�ۻ�yG��3�*v!���]P&�u����w�X�3���g��-���y�þ��p@�ԟ;�C�_z�rH��&�|�@���\f���1Pϙ�V�ɽ$%vԵ�(�}�F����k���b�m놿Y���ݣ�s�J�j���bv�1!HIS(|�k�|�ޥ"�V^3�8O~U��+<�;���P��.�٘fi��觿�8�� �]��d:��i������������<,��
ۖ��9u�"5 �!F��}��mE�|������C'8��8c�fk��L�%���n�5�.aX��'�E��bfnʫ���]^�Fn=���{᭬,�<�׍Ǹ�Nǅ'�<~��B���.������6^l��{�Ų����BL�|�Sb���zu���^�8T�G&0a4N�8�\D>��+`�.��pWm�8�!�ϐ{1����c1˭��<	;ꉡ 䖜�G���Jt/�`���o�6�0�/ű���S7y�h�h�)ӣ�Dp�k/&��Y^��
��%H��8�d��߸f��������5*�r�k���ɨ�X�xa�T����F��U�T�z���� ��[h�务�~;3�i���?vH�m�/6��k�&��ְ�v|�4=T���^�� j"vW����~WpInTlj���#:2	��{�r�n:�ȃQJ��ȣ����3^!��`	�e*�Cۄ��lS�dK v�"}�}����ϾJE6&��i٪haW���V&1�����l�oX=�Ln{�z��hԃ6dD[�0��}�:K{��o�'	I���H�9��wV���5aϖq��/�҆��z����b�.�0[������NO��F�s�~���m�݂"�YTrJ�$���^�'�p�]_�G>B������P���d ä=Y�A��!,q:rX�����l-[�qYQ��2X��0p�RM���p�+i?;[�S&/��޼��r@0͘�ϫ���v��:i~%F�`
e�����s��qo��o9e���.���3$ʶߜ�
����� �^m�����`��k�č.	{=�
`��j��Ǯ}�V�ԙ�
e���*hcQ�����eІѹ5f ���;sST���..�5�0���7�<rl	f�)����t��y����
*�$u��5�t��w���5�n��	�+�k"�s�$U����h�����љ.%T�{�*��}����7o�l1���T,8��2�)\_ ����yR��[ҢF�E�7�abꕓ����i�[�Sׄ,�;\Ǎ��w+�r+�ۿН��N����4lJU�4���n��3����}���5KA�z�X���
��aCSw�#-y����:��~�1�t���+ͥ�tJ�5�����:u�*
�������v4��S�\���7.0	�ڪ���#���n�*��s�&F#F|{�l�2�/Z:�ͥ)���2�,��c �а�s"��OέJ&�چ;3��$��n�������᰻�*O%�l��rl{kڹ1�&�H�0��Y���K�[���\>�~�9f��}�)p�A]|f�tq�� ��!h��&y�Ft2����q�)k�]ҿ�{9�6�O�g�ʪ�[�I0�,�d����2��O���k �l�w1�_��C`OW�|����V�.�9��l�3Bc���0K ��g`w���&��xaT��!%�c� H���P�������7���0�q�( yS)rVI'jzmt�n�nE����~�b�"��¨�	
%�
wK���A�^v�����<KUL��ep�Mƴ��*&#v1�)�EJ���Q���Eq?��SL�D�=��1	�?��¶�z�#�Fȧ��[E��a�<q@4��{����v1����jM�7�c"rV�u���͠xC�E���jD�)���錏�[���Ƅ*QW�}P��R>�j޺~!vv��H 4�BѠg��+L�	���(�S����p $�nO�&*(�|�_y�n!��J$<��A�/H�2��>�xB�S��z�~-�1ӷ�i�hic ����Gp?O�^".��MMX��%�L��	mWd��K��Lݍ��k	�D�>�NZ"WP}�@�$yҴ��,ΐ��%��9��)�ylV��D�T
p����|M<�U��($��6T:\8i����)B���%�1>��^7#$=��: ������}�x�1�P@�@��@�K�v��o �g[��S��~Ow��]e)K�~�(R���7(+P-e{���'~�J����Rh��Q5y��/K↔ǬT�|�
�b����g�B�9J�y�$~(r�6��[�nt8�� +&·Aqֲ ������2
���<[r�*��t&t�2ǹq��b�W�0�ؕ�P$6�8� �V{O2v��K�@�-4�,�i �hk��/L��=�3���v���I����r|�|4>wb5^�G��y�;m*�; X��� �?^N���!�yv�)i�ѳ/����ڥvBi3D�A����=�̄�
����$��M�O-$9��BŞ?�˟|ߦB4G�߫r�`6:�d�',�����;/�w:-ȩp��i�[XR(&���4���W�G��=p�U�Bz|�M��|F�u�*V�z*��.bQHk���;��!�������P�@��Y?a����׆�b=
����\=���M
X7�l]����6>⨏lU�h�cn	Hv�;d��q�j���!�������)�ݘ�_�hT_0����*fH���[�� I_���%,{�M#>��I.����+dg�=��ec~O�V7��Ip����3�i,n�1��fk+�v�8F���b�8��D�5���)���@*���7Qj�Frx�<ێ��a��@561�0	��?��?���Ab���J�(y�H��a=(_�ȭ�����;�V0s�hy��kM {��g���$���7�@� �+!°:{� ���Ũc�+�I*��&��S�s$�;ځ�1S��DTD�(�����
/�m�8��)�
�s��J5���<�b�z�]?"�����$
J�Gk4�]HJ�>�+��U�)ǣ]��M�6��.''=�^�_�m:��KbxT��3��� ���<_!��*�y�q�.�l0��y�c�h�KݪJ*$��㝉o�w�ݻsG����lJE^���O��wj-�d�ːB_�����zOFY	 �3=���Q�)ַ
�Л8f����]��ON8��li�ױ����-�A1�<��[!��b�ʛxnm�)cc#�^Źc5t����Y�^�lja�������4�Fo)�-JY����� p��[��[���x=��DZ&�����V�-��	g���������������t�^hn@���g����gV���O�!!̄b�#�>�X�}:݂�Ε'�����n���tIU�X���_Ȕ����|�h��(&���Q~ߔJ��Qbon��јk�BH��n���}n��h@k�s��* ]}�ǅ�������s��n �Փ⟬r��.$��5ע��qS�� ]�߀�����_�ᷫ��B%�mPh�`��	~����j����O�J�hk��q�)<� �n���@Q\|D�wŖ�����2���#���+P;��2�`1�Y�|Z�|����=|�kZ��݈J�c5�a@Զ_�C����6��lʢ{ԗH���T������j�WN47T�g�Pw�?N�Y@�$9������J��m�-{ͻo ��w`���v;Uf��?�%��T>�p�D9�ωS>�~��uo�D\�9�G?-�7Y� f!�29�����@�ڥ� ��h�薯!������Y��7R+���?�q~7������j�K�"$,�~P�QS�~�C�5i߻.(� �G4F��6�f���7_@q�du�p�"̊��}�����_阿j�?3>ܻ�S}aYfDc=�ݑ��żf��6i�@������ǗQ��k"3[��X>=���	����GϯT4 C�,w��Φ�y���l3���m�*t�[iЩqW�����T=$Y�٬�߮c��P�'H(�N�e#�E'N�[�`u��vm�J�ƯO;G%)�BD]��Y���E�m�f.��h�Q��1/f�n�R�3�d�i�j��s��op��@�D������~K���F:	��f�b����z=��	�F�Dȧ���pj$C���[�~����(�i}o���QZ����0Tw��及'���C*����e\}��R��r�6kꡜ�g�x��8�C�$��xjg�RP���v��d��R"�,
$����-f.W�?I��$hr܃*�Z
i[Z@��:l릯#1�D݉c�i �E���%�;��5�E&�T��`{2V�w[IG.�f���;�n9���a0��a� �CB��e��hn"1�������ժ)n�im�b�BG���Ҳ^��m�H�PET��J�w���BPs�����#�Էm�Q�2
!�eA�xBXM�ݞL&��E��Z�}t5v����Mm�F��֛.��/�֙�s�cK�*R�K��hH'K,� a���Bw����Iv�l�u�6E�q�K�@ˇ�,~E�q�L�����9���훈��������OP���B��Ƶ>z�F�2&�����)� �P������X<VF�(�Ya��ԋL�:ޔ_3�Kq�]Ǽ��u��Tu�k�콙�Ż�:�N���q�sg��V����Y�����sUӐp�lry�ڋ�D�&��&J�¬�C�xg�n8�#S'�
���S�W�;�N>
�k�M�WI+RV �m�/r����G��=��-_}�|�0��=�'3�\fk�.��Xy$�������#�V��X71�uCT(ȍ���G`9P�M
��oo� �Gd�����ɤ���5�d�j�/�.��/�Y��6Ӷ�b�/����:��g���\�A��_�6�6���l:�3��?]�*y�x�X_!'/Kt9��w�;��\�<f�ֵ�yW�R�s���� �E�CY�紗�?�C^�����$3X�)f� VV8
>�:�*�֏Z��^���j ����T���d�T�D�
o+�Hi�U�� �Afዤ��V"G�$v{�͔g�Vi/a3F\(�uǂ���زz-0�iu�6���� ����K�݄��2eN�E8 �V�ԶO�9�'��V�EB�1�*49�L3k�kt~
� o˔!BsE��צ�5����^)U�����d��(�5�'Չ���4��͛�p}��"+��Z?}��j�'0��j<?߹B� F3!:z�&}1� �h�c��y(i m�L]��y�`�-`^�K臅��
x��a{�Ӽ�ip�ߣIɰD��>������{�кܧ�ē\Pz�������s^�t^+�`���CUX�6ri��Gˇ�f�E��(EG٭�����LSNMy�g7���NkE�C��߂R�6��v:�>�*�4C���WT��dV�9�r	.?�t���$�gՎ��v��ãɷ���c�M-�f�B�ױh�#�SQ�t/3Cth�@y��.��U�Ъ�bx��9��Au��h�:�Ϩ��̳*�e������p]���i*�Vq8��l�Uۢ>E8���6��<GP"F8%GX���U�@������#�V:�x�y(��\����u��aP@<Tt�N���j���X��5υ���ȩ��n�q������@�9H���+�@7.{BER;�Sfg-����j袪�^��-�R�S&��G����*������I)C��<n�� �fӱ�+ڎ5�[4GXj>��"��Yݰ�s�|]�e�+/�fr��>�l�1��˚�^��;��xΚe?����:���s[y ��QBiB;3�?���E�)��u�{lQ�wf��I��DoaM.����α7�����V�sj>�0�J�Q#�	�KZ�@.)6�;%�;S�}�Hl;Dg��Z�����N���,6Ҷ��"	�ƣl�|�s��;w]*�w<�ǌH����2l�.�l�b&�JfjR���!��Gl�i��MΫpST���֪��}E�����q�-����n�-��?�dBC�����5v_|P��Ӡ+���ue���9	n��*!�=۪��F������T4�Y6bxy-ׂ}���_�oE��C��T�G&׶B��Sq&���)�^D!��v G.����a�0�X��x�嵷�9�jMrH��/����c�h�҉�? j/U�V	�F]WS{��p�(���1�tTaқ��P(�{dyA]0��HZ�Yhv{�H�7��t^�W��0�~�L��
g�=��N6�_v&���qX��	�aY�)�S�kW��"�b�T�fW)�!�^R/#m,��ז5>LQŰ�Tr'v���6૫�#o�|f�h9��Yu��iN֠�C�����ڡ��M�Ń���^�-�|N���D'�k{�1�H�����dG-��c��C~|[C�� �l_eI`[�m�͂�k�eڙ+�%�q�G[�����q�; T��\��62͞k�f���*�lf�b��ZQ#�s��U
�8�b�^<!~��8���:,�V��=�{��]���.�K�t'�H�Cpb��ˠq��ҌV�	$y�R�Ţ,��m�Cq��]&?�"C����Wd$�r&�pV�ө�_S{[��J4Ŷr �>p��V[��
� �3��
y&H���3{�`�_�&>�*h�s�r�QĐ�)�e6�%a�n�������6dAʶw�[��F�d�ǜ����b�}��/�_���pJt���׺��)��pĖ��� .

�b���ѓ����{F1�2�2�q���e�?���c@X*��R��[N]�o�I�*���iuG�G���
6��{��J�ͥ���������VZ)M"2��JR�{w���\cG�F��Wx�P��ݛs��B5ɫ��͔]h{.+�ԡ&��%�:Q��6�0k"���#6H+`c���Fk&����x����+�:����S����4�	Q��4;�7ӚbVj��%����֮î�a�����HG���3ճ$��m��D�/M�������DDP"��x�~��W��"=q.m���g`�ቸd���g3,X�80���\&t�,�K��F���yV�	g�-�)W����P���奜�@��٪c�p�]W��_���r�h��U�!� -�^2����G�;��G��SI�@+�lm���Z2=�鷠�a��8��q~�G
BBuI����@V�ʰ"��� ����F�Yz���n�n9tˀ!�W��.�u�W<�hq�W��,0��
����"e+�'�_��� �d�|!p���:6WF���]oω��B�l���R�q�:P��u�ۉ�Qƿ�Rq�ݔxP�a�c�gv��u�6nRb���3���6�t{t oo�`Kې��@yR�8���[�r��=�yP��S��Q�f��M#݋�˩��C䐙�t>������@?�'���>6����m���K8����1ZfO#��C�i���`unK��i��:N�)��x���6p3kSʸ��+�/� �l�-�[��i�����f-���L��3u����A���:U�����n'�9��1
��z>O4��ƈ�4Ie��#�-f���K(3��K��& ��t
oaA�,��(���I`���iV�3x��i������	O)�_����F?���[<�'����]�_��M#|�>z�ɠ�y�W�����8��M�+L��&YΩfG�p1t�>� ����Vn.6Σ�\���u��+S��GD'7`1}	��w>cq�?�RZV�e�4��O�j6ӗ*H"
���(�\�ˈ�3O�&�(C� ˖��sE?_b*�� ��{Q\j8K��C�l��d;?sb�^Ԓ���?c�s���UM�.����H�"Vf�1�r�5�/�D������VaB�[�EI�V��H�E�1�O��5��Q�)��'
\�^9;��<nN��u���1�ð@��z��Zl��Ll͇���B��M�b)k4�
��F�C�ރp��](`�Қ�ֈRo�����}�E���;��%���hfi������K!�3�N���c�ҍ�?�6 =n���U�ef��ARS�H�!��[��� �W�~���*(y�a�g���:ݴ��Y���ܰ�v��3q�@W� ﾷƓ�,`D���B�GqI)I�F:�.�)�	�V�+Y�'�nsT�8;RT@�Q��p�o�T1�Zj �l��^fS�1���xyL���o]#�it�ԳͰ�?�v���X���y!J,�Z7�0��gz��U�nJI��*��;���=,��DD�uM�%����Ex�':
��a\scٜ=`�.��\������S�t���"���=݄�p5��2��MeS��?)~{�D��S6�����WR81�,�x^fwT�`�?�����G�O��@C�� A;�N�x9�%OzuL�fRO��L����/�Z�ox��]�����!d�_�KA2��2�\�T	/�_��C��r�tM�H]�&�j��2lh�._RZz��ƀ�:����ӈsv��[�Q��g$��������6�XA��!8���,����灙�`��nRM�$
��,Tg�>Z ��/��iV �G#�ɀqn�=,�8���@\y%M��ǚ���3��y
��z�z�1�/�l,LϹ�8VU OK7w>��J}mQ�~�
�r_��C$�-g�~� �u�"�+���Ra�|bP	�Ty鄮��Ӎ��/�|I�X���_:���q�Ԭ�ȉ��\y�a�r[̗I����Vy�G�
S�V��O"��Qo=m�F:]"������^��,#޵G�t���{���db ��D�9:$>�|.@s��8���om���	�7}�'�u���!g��<�CӧR�4�I��dJ�Z���s��>��b�q��m�r�HMo�������~Ru|B��J���+�$B�H��h<�21y���Q�>��<B�X��!u������ʅa;^���y����W�%�����%'��gQ��y.�ŢA; ���L~QŉK��j0���c�K��{����b,� ]��,N�f���w�D;w�a^��3����c�(p�P�hl��K^(d�V�F�
��:�X�V:�鏞L���i�-9Q?��	�/3��:�W�{����GK��`ȕ��_�K|�󤭨0��|KJJ}�%���n[�ξ�`�1�["TM8�w���C^&-"#?ݪ�_o�:�S����7���T7fI��~��<�a����ŗ9��l�	)����q�t��F9���޹Etș���t��)��gev�òa����Yhϳ��C��B4��¾���c,�Z�|h�P�%e1�tmR�e=C�=���(��y��j�i�]��_g���t )8�6��@O0Hxz�:(�p0��aL����kQ�h��RĜ�k2����N���Te]Q�g�H�
����숣j?����Q�'�v�9�K�%�����*B̀���$ ��S���',U��md�̠
���Σ��GB�3{ܝ�jt���w�@���!�t�'(��$֑��lb�r���U}ݎ)�*�xL@�����
�Cm$e0���l�� ^�=Q?�GoHv�:Kܸ"o.����s{,��<T1{�෧��g�/�_1r �����_��4q(z�<L�I�ۚ��*�?��p�YX@�����V�����Ӽp!O��r�I%�X���x6�r�0���4#f�hv�&�:���u�*b�[c��d���_�0��'`��� ~������<�I~d��>�CK�x���'PD��u�TM��2����͎Eg��M�zUo���L��_�%�- 'F��Ӝ^�Gl�Է���<��U�~2�ɷa\i;w���z
��a���d_�,3�,n��q�!T�㢤����HvÉ(�9 �;��ȕ�Z�e��r�m%���i>١=���S�8q�џ����@蓢���˽p�\��FlM�DE�u��	Dz!&����B�ޏ-i]z-�}eK�v�/��&}O��;1q]�/IʲG�T�Δ��!����";�_�0=�|7L����#=,��=������%|zU��+'h�\�$g�-���*�%�; 6��F_�Ӧ�hy��Y��p��d`7��D�b��*�S�-3á)���Q��`��s'��7$a~�\����25>��R����YQ= i�ݍ���s ��-�gL?��r�j�v�g�"Z�^��E�%�$*~o貍H�6�����@��m��;U��NPq��U+*]|YrM~�Xj��4K<��e�m��b�\u�����z4s��UX��O���6�g[d`Fp<���O׵<�F)�k��zѡ
���L�?;����G�Z�����P���p���
H*(i�UI'�k.V��|���-�T�x���� �������5nNC���#����.�2����
cw2}�o(P��H�tF�� o]/� i^����:��v�
��x%�u�#�SQ^���5_��nK�����޹��i�_��ǚMq8DG!Oo$�+8f��'R�B��/�����6�+��~i�2B�lͷX�=�G1���󬂻�W"ə��������ƃ?�+P[Bdj��oQ�	םφ@Wˣ��ո_�n�ʒS6#�I�y��-�0���腝�M�I0R��"�j׽\3��7Ҕ*�g�A��#Ā�$u�ӑL�üR��V�ý8c� G�:.l!�$��zuh� �}l����;K�AVaK�R[m,����!=�j1Y�~N�J{Z���9�����=n��k��� P(C���1t�?��t�	p]7���P�:&�%��6rG�*0�m٘ ڻH�Ձ���v�a�(E�,Q6��OT�G)���1g%��uX����q@Z#є����?SS�Ȫ�JW��AH���3pِ�{�c��;o�Z��_nc#�;�v{�eե<�3���2-"B�*��Kc�W������+Xj*D��9ȋ���3m��ђ'����޶�̒Mrj��F������aF�HM�Q�@q�P�㪈<�xL2�z	e��J8���Q��/A�3oɄ��S�E��DB9P�H�)>*i0�/��x)�����We��#ƽnu#�a��cd:�d����@��7�G}H��SCn�S��ba���WЪxзru���Q�?�α��}�:� �����(�d�������K�����y��B+���sz��vq?.��Kj�}��H�,�掱U�7�@�F��P횏<=|�ylM\dkϟ�3�,�#���F����=��a�v�����$�h=+�����{[�p��՜�m��1�p�����m7�e
.p�?U��Ώޘ�t?�����C�i:�$o"��������,�z&�K��u�i��Z����A���r\��G����h�$�~��*ɶ�pݯ��j�3$�ťO�V;��iOMSA'
j��B�D��''9�X������:�y���d�Ⱦ�J�:6�NT�����LT�=5�2d�����6�Ak��뗒�����쁹M�C_���k�*�ar�����>�e�,h!��&��f�|��YM�N	D1o���o 'Ga�[2ePqg�]5ŦAw��ꋾŤ���Ve��=:�J�w��Ì;���;M��Es�E��R{{?��_3 >8��.�#�u�A*��=������˩���3ZR������L���;R�f�q�)bco�5c�Ҍ�{
m�����С�w�v�Qs�΄�I����Ʃ���<�xbQ�
�1K��ո�Џ&HO�����'X��8{��|ݓ�J��l=�Eo�s(�դ?,i�be��HR�g(����C�3b��� xyP�ϓt���S���sh��Лh;'\T��)��焛 ���o�W�:�q���9i�4���T��a�pJMق�W.H�j�iA0~GÛjM��V����G�� ��S��đ����4_WN����Y��i�t8�"Fء4aR�J1.�o/�0�4�S_o!�����-�EޗJ�Z���P�W����Xǜ&�^���]�$k�����>*C �@[&mR�?>9B!]�e�瘟�EGE���<7�_�4Im�"�P ���C˻��3���!�Va�5ޝ�t�y�1oO���y��(	Ύk������Re�@�Zf yW����Ƒ,�`��Uo�:���P܃��On*-Z�N�Z��^��[ʏ:}/�u:�e<G��ncA|tˇ��l��S	B��ry�]�4��%�5�yI��k�Q��X֋G�UA�;MtM#�w]��'T�¨Q���܅:�F�J�5�`��"���,�|���O� Sy���[�<�����l�#$g�/�@�.tf����+�ˤ��םO�R,�b�̟`���P�a+�+(2���[���������0�2��}�|ي�6h�l�O����b���^�%�����hh�p�6UeI'FwZ�'�+ABy���U���myѸ��ɚ�$�+,��WrO*j�w*��k�S���+�;�I�$�L��K�|��S��`�s�6�m��ڬI��5���a b�%v���+�]�t��h�ŸvQ�D�	�僊��Ms��kr.��>Q�\PH�*����BD{�r5;(f�L.l�^}�y��|�����d-��.9s#
>��Q��#�rl}�w���3��N���4kp-�פ[68F�Q�c�K��їE^�����_th���@j�v&�ѭ�E���@������u�q�϶BȔ�}�V�_ԧI4�8��� `z<���儜�g~< �{�Pz��q8Bn�b����#�)e�̛���e[V��Co�D��)�f���ش��4���u�
r!5"��٫N'��c�z�nQr��W�$v��--f�Ψ ��V��f��w�i��ڛ����x�A�$�zy@s\C���"����S5��7��Dxn����C�R�]�7@Nj�Iτ��z�E�%d�� ��d�ĨW��<�-�垡�'n�-���o��{�����ARdp��jf��'H�k\�wDYF�}��x�أ���Be>�(��%�$kI%���Q<hJ�'��ko��+e��_�S�)�Ef�dZE;X4�m}�!�&��d ����6��K���t���p?�EJ\l%wj\����
UV��S����
+%QB 2�Q�;�5��_���%����:���~�j�Ց�7�և�N�Hw{��b(9��Ap��)�:i�	����:�-����ִ���z=�e�pH*}C�]-_r6�p"'=w[�C�kb���	�O���xhw�1p��8&�M�k��>��hpJ�4ص!��*�Fm~H#�}d�h��l��U��g����.;`� �C�����r��)���+e�-���l�˹v�J"�yՖ����C ���G]����0�7���dv�Au�r�{�"��-�"�6M
�������$�B��Am��_��L�nb�4��{�Pp��]�K��Z˻�_���\��pA�O����vJ�;5.�`���S��M��tj���Q��j��,vWj��,��v�I��w��sp�f��Kz���r�L��c���?�).�:�ok�`��DU�Gr�m1��cz��TڕP���ݑ����a�w��&S�x��kk�{��ǽBg����ͤ�I������d�dA ��f�@Ȳ�Z�\�h���0�(-�8������W�5��@����n�y������V���G ��Q0T˘����4�@�H����P�%m� n�?B�(�H������ܙo+v� �/I{]!Ws�W7��9�*�#Z}�:u"*i6Z��A҉o���iJ��g=q�4�.��u��|�7-ꉧT�E�C��ڍ m�`��Xx7��3�MS��A��'��F�0%��� �Wǎ�?|G�I��.��=~���7Ժk ]���z���/'ʗ���>ԟ�K�D�컉��J	�h,�}�������,�RU��:sx����2I�Ba�[��8$��-�p����\� [�$�xd�(����@i�X>`��P����$��}��n>rxl̜���܄�m}!>�wŘ�Ќd�L�Lx0hЍ|�Ǔ�Fs��s��%��ꔐ��y��w�����l���R��?h�q�ڸY2`v��Эmi5�_,����I2E�W�Ak���5S@N=)���3eu����}p��U ���61�G����y��vl��}�N�Ģ㜥4�ut�	��d[��٫}����ẉs�LR���d����$�h�M�b6[��SV��z��*�MZ��x�"���3u��Y�zn���?��e��4�Mr�?Т<�,7�y�O�)v��K�I��v)�J�,+��^`}��t�/_�^3�5j�r�R���QB�z���yx��3B�l���3L�{��Ag>ˎ�/]�w���?'���ظ�_ī��Ub&��ϱ���os�ஔ�ꐪ�։�ؔt��0\���Q9F*b���l�\�>� "�ײ��*1��Wje<���9��.��*B�=�)UF�]�_���^D~:)�29��\��T�I����V�����95��L�#+�'r��J���4�]}��� ����`�k��!\؟���²�d�_�8,n���i�T���Vh�j��^<�G�nkcFއyҗ��A���pj7%#�ih>�B̨��m_�v�)��+Wޜ4h,�'��H&�W�˸��4���O_h�3
�In��pƚe�;H
|$��j�W?s^�N8l�@�}v�!M�MH*��y��������^4r�����D`35��*���;_���d��g��Y��c��2�%Q�o�w��HC\[a#��Rɉ}ݺU��M�?�g���r���X���S�+9�@�QA�`}z�^5�W`��+q^�"���S��
�H�Q�IJ���A/%�	q�f����I�^�3�<7���S(��ި6L���P���[O�!B�KR�} ��~�B#��Ji3���w��%�{̑#��q���fG}�A�{��6Ny9���B�۩�.%�o��A���H�r8*	2������fU�:��@�fb|��s�&n9*Xe+���QWA������m�e���xZ'���CԊuF�E|�}�{�B����[_�������#�v2���
��?�EW]�}��<�#3�}Zx�i<ܣ�uԽ/6��((d*�+����D�Ρ�|����
6K����g<�ɋ!y���x3 �T����5��JI0��?/FF�%�Ee�8����Xʂh0��J�W���U_m� a���.��A��W"�#��O������C���������TͲ�B�68:l�Kh�bv�xSp���8G�㌴�R%�@5N��$e\|�,�7c`�7Z��7@�8���f���vP�С~!8>��.����7�ckEb�U��d5�\>mdG��
ݶT<h,�1���׾��B�|�%���OЖb��hf���?��_�ϭp���+^�1�k3�߉Y�R�6+�f��F�-X�R%�PJ����;v69���v����ϱt�ha��c��j���[��a��[�(0�'���L�ݎ�֦E&5B���J"�*���}���;�d�M28⍸~�hN�u�9#�wP���,�_���!���]j�s�0?��ꁳ��-��_��	�8����Xu��;�#�f��3%�v��*�&L�Dv��~I��+�p� �&Ɩw~j�ID�h������+:�h4aҮ���V�(?j�H�JΙ#P����	������W���Yk9Մt�4?
��x|�痺�0���,�� � 0���י���i[��L�:�I�9KDZ׈(+P&�~'eduk�f��nk��~4M���� �N�W�Ȍ�D���w�62���� ^�d�����b� �r1"��F0�`�]�E�1. .ᛶ�mI��Γ�DDQ.%89�Q�g�Q̏1�?�zH����+�ZV��ck=pc���s!j�r�֪}F�5yOU����U~�o�<S���9ȭc���B�������֧�|���t�^��R7��2�_7��)�o8Ô/|#-f����.|�=��=�n�̕F�^��&3CZD��"[�N� #�X��G}ҭ���'i�[�ȯ0��8�.�|�;���i�[zW׋v�V��p�X�i��'�G¡S۝6`�F߂'�񢖃v�}o<�_fv��V,+���Fb�5�L�K	����;���������m� o^
���	��%��D�&I�\��Bg �[�L�` ���<VȾ�Zq���N;W�S#�щ����x|�%�4W6Z{�w�]�\l���H���N�xT���+���]؄V8~�o�pi�W��`���]�Fd~W�&H��]�࣭�xx�3 �Bu��-՟��d���ʳR���d9u٢�"a��]F/0m��5Ι��|��3Ô���q
 \W���qd��
�wk\��çޅC���c��L���
G����-�!f�]w�]���@���,�Ե#�@�9maO	p�߹+T��I�b�7���P�20F3��j���"J�ӽ�I��
��*���;�����C]��PX��t���)��O7�jg����V���z���ز������r��SѮ�C�S���;<�S����C�Z
7��h�s �o���&�/�Lz�l��*�y����$]���%�����zD�$,�Qq���Ӛ;>P�E�����R��`Q���]�|%?�&��6�lXa����x�h�<k����
�L4`DXPZ:JC����O��b����K��$ �s@�i�`�R���q޳���}�4��#u�0�I�=[��V�0 �ʜ�3BO���-�!��w;�r�6\�m�;����;�Yf����@�ki��LI!S���o"N16�g���Ͱ�W�[�g�e���2_�����Cm@� ڡ`�g��� g)R&���NՏ�L�����.kK�EYj���y��z�'sס�n��nb��v�̀�5䱕�=�{��<��G�"�6��@�����S��M�C�*�rm�'+�����D<v}]�oyL�j'w�xf�qh�h�E×�
b�Ǡ��K�g�B�9h%�P$�xz2���wߴf����*����>;T;[�?֥��� 0�!1�Ft��(H��8[����g��pT���f����p�C�CY�9�e�ȼ�|u��+N3�XR�)����ܹ�s��K��R���'��3�J��1�I������n�nJ��SE	J-I,��3{��g�+�A�/�6U����英Ŭ�o���xYޢ�%����
�DN.юdƃ;ٕ>fBR��]�B��~�H�h��*���j��A'DXln�*N���A���#�wa��x9$!Ih��	ۃ��X�fāg��u���C3Y�(�jQ��$���y��}��p!gݦ�l��2m.'�ҸA�y|��T$��?�)|�W$"���J�OЉP���m�_U��>�g��Zf�U�t�p2��L��0wۧe50[J���:�k�خF�� �R�|rAj�Y�Lo��oLszy ���=�\��i�MT���i�X�{���8��'�Y�	�O�ë��G@��)�4d��ig����h��wtGE]H4?q�)Q��rX &,5�K���w�'<�'B����à*��ʃ��E<��O�_sr�F����ac^���
�>6�?A�B�%]��QݤUAs�i��BX��ų�����o����!6M���V.��~��%�A�\ŲFf���`����#غ�P��tfvbB����X�%�q
�+?!Bem�iG<A�p�%�|_�5 Um�	E�3�/�!@d6��/g�}�~���%�_�����&�*��-���RQ��A�: [ZO�X��� Ed6C��{�3��W��H��a-��N�	�3�0�G17+�h���E �'��U���T�虦"��Y����3�����f��C#�Y/X����=Σ�Yp����r�wG���tArI�q�w �S�����K�Nh�$_S�wM�s0lƢ�!�T��V��L#�m< y���\W��d�����x`1��C�f��,}#b�=��Ek�F�� �u/6r��ff8����>�5�.����Q���΃]��wC�wΧ�&� J�D��j"&�o�QU��V���HDF|�L?<p�cjjn�����f�#l�l��B��E�k�N��F�N��hXJG9�J@5�[���oW�OX8����t��'�� M�ڷ~�^��t�?�J)whx�J��l�����IC�Fu�9���\=�uRV������sf}��_#�<��)'W���IAP�[t[K>Yh��?������[�K��p��e�
������&�B��M�X��|;�S.�Y��X
S�+_�<�p�`�V�f�F�.�ި��r��ω���r�o*^?)���g��m�ba�
u��IC��h����g�?4r��2j����$�b��
���c�:o5g��t�|]�_1Ⱦ���T址ǕWө�������'�f��~"/#A��W:u�B�+A
>����;��Fz�7����A���q@��a�L�;L&�T�N�Y���x$����G�u}jb�_�/��)���n��Ǝ��!0����n��!z��������M�2�WΝ�"�9{lYz/��o�3;jo����V��ѽ��5aaW��W0'�\@�'����X�w��}��ȳ��A��$8x�Lm&�{�
�u� XN�e3��R�h�y�c+0��m]����n�s�B}O��Q��0���h��tj���ǽ�����tcU��])!�b��;2�(ȫ�"��	�	E���n���x���
��f��2`=������~�q�)>��#�V����L���y�D���
�:�g�� 9Z��^�Dki�ҹ@�י{��,y ���؉�'��N��Ȇ���rb�0��ɄC��p&!7�@g�X�+%�#Q�C�&�a&Q�_�a4ȯn�Ш'�t�~���'l�6���}D'KI�N�� k�RnS�h��P5l����h6��fS=�ߒOex2㎉�gH�Z����^Z�llZ<�r	lP[7Jzt���8, ;�S�"�C��b�'��"�bH�@�C7�v� ͩs��������a��)��t�<���U�/�s����7c��#J�Jg��.�0�떭ɫ�=��"�j�$QӉA��P�`��-K�����(���U����:�-�Р0Ka��r�P�mv��3]ߖ���Mp�!>X���P�.�k�����%�S)7��%'�S��V|,g��_jt��m�깃ܷ�,F,Xh�Xs���S�@h�/��A;
�M����-�/i�V����ߒ|ln)h��%}�X_&�,L��k[�r��J�.�E����];8s/$��!���.�"�aK������!����E�6�?<��6���A�#����&����uRt�h�X�"�>���ߜ���L\l	*/1��z��P�F��ݷ=�O����U�1�p��-���F�=��-d�͙�ѓv1D0P���h�Ixҽ���
� [�pXKa�*E�J���i���Z�^g����N,����|q���B$�<���/kLx���}a��6=����,��M�\�g�,ݥ�L�\�\�8�/��H'h�1ƄiS�~^���|�%�l�	���-"_<��	�?��/Q�9�<5B��6�Rp��7��D*fP��#JQ2��,YU^S�u�kns����[^J1a<����d��v�:U��>�,5����bҥ� ��g�)ev�P�N����$��b �z׀6GҦ�)FQm��s(�c���(�q9�3�|h���/1�;�y�d�;8e�o���Xo>����v�9Y��P��R8
č��J���MD��@��u7:��ؚ���Z���K����Qz�\����q:]F�ˌs��q���{M��%�ɸ�g��>쾅
�$�7�ú�H�8 \K�� �)T�U*>�F���f ��9�籾{Xo�o���$���>�~���(�#���@o�!N��OϜ�!
1�9�zKK��j�ƫ���Mkl�ͅ[�>�y��m9�����-5�'M�����'	���4������{�t�kp"9�9��?٦^���|�t�#'`�7���L/ƹ�ԬPm��l )�@՟D��/2�#S�_��Ǿ�V/6��=7D��nv��uZ��F������*�������f9�OE�~��<W�������}��%T��h��(��o���6vN#w������2U��L��xC�˙���q�i�ؖ���XF�@R��!�*A����~�iб��x���O��Q�ߖ�bS�KDe���~�/U�t*6S�{�=%�i� �����Ͱ�Gu��MȲI��}�q�\up��������M���3x��g��	�&\Jg�� Wz�	�ݿ2"i� B���	�K�l�����3ʢ5Tҧ2�]���8�}����N1��&��[y����򹋺��Z�2��E-͐Ԁ+�%-_�	z~�>˗�����b�0EL���M�	0<q��)�׋S���l�T����b��,���_<�W���K��mG��[�{�V�츊r0Kױ	A������������	*��x٘�8�*몆�{�5�<La�Qk�;��{�Q9�����'���{��b�)�`�/W0����^��"9�9��s�ŕ2ӑ�'\�t��B�����~﫳��I1�	4~��1&y�<$>��dP��3D`u]��UnfB\8�y0
@Kg��y��}�מ�'�-��ێ����f���������糡�:�s*��	��5�E�a����j����%��O"M���MGg�4x��:���1�VRl�bV`_��s���R�7,�|6eK�F֩�s���n8jߥQo��r���n|t13@������C�E�Sv*���y� �}�����l�"�G��$��������\�D�%�S��y�hM�Ӻqd,T�r~7�u�'����J�'^g��������r�n�*"cbQ��0c����>���9,�MC��w�\���#rs�^T#�p�	1����b��' ����C vL��V���==��X���]ʫjtNz��<���=�b�~��j�b�4����ۃ'��"�qH��y`���u���4]|�-vOX����Ȫ}R�Y4>�:!a��!��x.H��u��/^����V�%]��V�O))�+��=`O���ł�bti��w�i�'R��)��W!0�'���K6j,�Ne�B�z�ߺ�$�h#�]=��#v��Nà�����dB��3\=��`���[9Zɋ��Ss�$�^Ͻ�e	�ɣ�����W�y�H�Fv���+ N���j�%�&2������Ώ�ԟF��

 ��`�a��uc�7(��޻�^}ȵ���;��@�T;^�o��q� �;�"�*��m�E�8o4�`dȕ�V���u�V3xx�Nsw��`E�I�_
�o���<���3���N�(�<����۴|z���� 7���A�˜H��b�M�}�ti��`
Nc2�]�D�|��Ell����c�o�t��pڛ��Q!���o�l�s{l��uۚ�-�*���c�ئ-�0�v�8�OI��E&wOcs�d��J=���
.GK`Su{��ɦD|�'���e� DW�g�ن߮�(M+K��w3
Н;UC?��yw�!�‣���w`��h;�9��Dr���rf�U����ٗX*_��0?j�hI��j~@#�qA,Ϊ+OX�Ց�gh�i��yr��ةf���钕qb�M�{���F�;�M��4^g͕�F�F���&��I5�*�FF����gi�w��u�^W*΅�p{�n3,_���Q~�
��P��1�J��!�^qu���4aTQ��c�7��
�B��Cι��ha	M�?u"���k_b�e5��1!�g��!_���v2*��l~u��Ll�.��{�U���mD.5�ʝ��&c��Xaա���4a�p#�grT3h��4���b|p�.�8�l��Mز����71��a�ć���P|�v6l��K;ҹ���c&[$&)��S�[UC:���z�^!nX���o���W:�N�������I������$E����ǽ��
ȃ7 yg��u)B�;��V����h��⑮��_b �GW����������]u�ʔ�bN]���+y�њ�Z��FHW�ǜ���?4H���Dg.�3o���� �I�"GT�ز�GF�|���PJqy>�+��#�ְ�[EJ6�3_��	%!��`;��1�-_8�G^bIm���bofu]���DJsJ���n �&�jo }L���`�7|���[+��Tj��S�[���O�c�-�RQ���8D9J$�OW{����R���.�i��'G>��DEQ?VB�$	�T�<���\z��R�غ8��2�m�Z����kr@��~;���
 {���L� C�.u��eB�G����`怊�?Ð��f=fڛ-��W
'�{>�n��t��7 "׳gBd�r�Pk�!Cz��c�S}8�|���`#�Y��V�T�1�`5��VHU���E���g��ֆ�8/�W	����4�iژ�`>Nu`�i)��9�;?�I��n�����L��;�*K�8�$ꓳL�ő��X���ǐL��REL(�q�_0��[{��y����~��x"�I�^Kz0�7��-U��4�דb�ٙ~�%M@+h��XX�݈2�y�$�!��i�Ng��ZP�m�U�;.��C}q�~0D�f,�7E����7?��!�IV|n�~=�I�'<8��c�fv��3��8W��;�M��$v��5jȘ�C��ƺ��҄!�Ɨ�R�������M@��8���G7ZE0f�"�`��"��m>ɟѰgꓡ}��<��5�)���ZZ��;�W�̗ݤ�FS��o�\���v�(ڜ��ad������	)5�)�kpem������_bD Z3r�Z�#�YV�芛��O�� �\Ɍ�`�ZR�������$��KeI��NR����m���]�oƢG;[��ģt��,U{X��-c����_�!u_�	��v��-�>��oM;�Cjs�7-��v����u�Ǟp���듡a���%�g�ުǏJ��R [��GH�J�xL���1w���C̺n��q�#V�E��;bG[����<V��2�J
W�
gd1��D�T�~ɩ�������xt$����/�cKN������g��A~�r�Q��&t��gƛC{y����/�M�Z2�=b��%��2��Z��f���q�g��{�R�)�[&fR�(�]8��j� ��e�[o?A�q֒dN�&9̽>�l��$�LUb]|�	�:�Y�rpvǕ"(���ZD��GZ�A��D�H.�V"Q8����\�מB9��f
�l���@Cy=-9�of�`="�X�q�������_ي0j�9���A�>f�a̓�=�kSk�h`��n�U���֑��S�!��g%��b��E`tB��������fM���p��0�^�̾�4d��鼙wM�fd�A�Z[��/��B=��vC��=������ ��Mo���k�N=��4 �̮"�n����;�BͶ�3Q(�Jn�B�n)\���A�~�B�#���a�fuZ@[�����2�
fdO�8���Z�����W�mo q�vP��%Ȱ����o��D��~��%Y�\����{I�k�f܃�c�:�CK�fJ�m�M��������K��������$(7$%
Q�u��j�x��R]BN���cM��N	{�o�3E��b��)�^f��=Wr@\��j�g�Ew���`�mK�е1p�'�]ْ�C����ވ��&+_�0��"N��䥑���U0�$7��0�id�f�'Rk��=|�n��1�V�^��ӝTY�^(�d�@������;(�j$���]>uu��H$\��H�GI�������E"�o���iDN*��jM���̺���K���so���#N�* �p��$z�Y�훣q�c�$$� B��T3���3��Su�S8n����y���D����h�޶G�槛����Ԇ���3��j e��"��;�xp����߇LD7IV�&��K�Y�^"&7	�ӬpK�-u����Q{�'(�=j�l�Z>�	(�����=[Z?9�	GO�\QO�zi&΂�����ȅ8�a ���2V�����_�s?>�X�G�UP+�Ԯ�ţDͱg��
m¨(Ƞgi�����6!`���V���w����/-��4-`����y����qj�A��譼��꫸M��q�=ϰҧQ��N]ŎK-��Pf#,g���3@��٤�D�i�v���hV��`YV�6����P��k\�`0u�O�}-5�p�mS������$�iPf'�����i�u�bziMuh��W8#is#�3�o�R���_�g*�x��"�c
4��q�r̯��e��D�$$|ѣL$J�r�	A�o,�ܕ~�p�z��n �3�E�s`����!yr4]�����C���})�����J�ڬ�A��^E���~�W?�̣�ap�K�L	T���k᜹�&�P$ng����1��*�1�_�p��ﮊ_���qB���~��� ꜑s�����n*�2�m��l��J��V�t��8(�s��ڝ3wRo���:����c�L�F�a��1�?�n���L	Y(��(�j��Q: Ht6>
G��u��̛�zB���&��9�C�^sH��8�mX�ۖ�"�kH�K����|j�Lot�:5rOig�</��s��w����5bo�Q��:O�(h��I
*��,��.�� \x��e�U�ԏJ )1���l	����f�~J�陝Z��96���)u.�,T�	g׫mZ�0�@	�mx)�3\}K�Bw7��w͒i��M����^���yE� �a9l�XF�hkj���=+.��M�.TwRn�8�k�4�)`�w[��}���\��ɇ��S�>ϓ��vWG�	�'fzƖ�����b�y�v.�wU2me��PZȠ�+X(�y��Y.2�,�c([6;W�=VJ�>�>dQn��ǋ� t	c�µ��8��m�E�����w��&�Id��j�o?�:5���˚�2�4^�S�̏�B�g"����0���.�`G�r҂:��%(���C
Z(h�/궈nhv!�����L����1o�V���T�p%����v��ܤ�� l@J�ď��Ɵ&�mX
��9�����(k- lS�|!����y���~j"���<�gk��j:u���k�i�|��]_�^�hw���'���y}퇱�	��4���$uY��rC��D�Yɾvv�8�>9q2]�X��°[�;q�P�4�����?���^�X�F[!��*[���:�� #��2���{���l�R�ЁW������v�t��q��IC�C�~u\Pס3��̓P��ݹ
O|�/��$�)�<&��1�p��^�� �hw��G2�n}�F�t���X�����+��bN,�Tc�K��wN����L�1C�¢�����f��R�r�i4�no��j��/V����y��m����ưtA`Ԋ�W�b�#�a'��ž���i�Y]i.Nxܾ/1��R� ���ßz���^��?&H���Z���2?���(��us�/F����}�V�Q8��PJ߷l�M�l�H��s����O+�\�)�Bǔ0��Dl�L���@0���Av`%��0Ͽ����a��DO��E�����T��[B���ث#���"*D|�b�)���ߓ����foɤ�0��bX��ț3H߽k.ga����Wwu'����t�\3�V�k�Ś��i�Ԏ$}+�K)�G�8��R���n�n�`��xoW�&��8q"�Iɠ���P=��{ɇ߄qc��?�!C��ql��Tğ���Co�d�����m�%Ƨ � �W����բ��i�j]w9q�yRm\���]z���w��<̉e<6Wʚ��ϋ�j�4We�MS�D髦3�q+b�.�C؃ � �'��Yk_���!W��b\��֓��4�h��aB�{�<BZ|�4������SH�+55�� LI���1�n`����%w�f&�IĽ����ݐ϶+�����ƲU���1�<%���~��F⁪����K?�rX�=�.�q���@x	N?�.����ݞ�;l��&�?��S�Do��뤮Z�Qes� ę�6�&���t�F�o�	����|�i@�����[G�`�^"k�h�n�t3,S����3������!!���i�o%du�(B�TŗJ�����0��.4���uړ���c�����2n�C�Cո�Y����Ue����9Y\@� q�����f]�y�+�m^�508���^!qSڨk�E�����Ӿm����G sl�d��f��K関�O��U��Ő��a��r;��D��.qC5q�i��h˱���ʩ�Ha*�mŖ%f%��g"�,��yo�VQ���h��O���zd�H���yiN�ls3�_%ſ�H�T��X����,�����f©��:Ǜ %J�����j��A�Ӎz�Q��~%Xɋ�rzǐwcۄh�Z��.��̩��*�,�D}��5 �J��;=��}���3��;z�K�ݹ�mB��F1�9��`�uYkVX�/e�ٍ��r��3�����u8L��	�����}���̈8����AM>�yq�`@t�y*������v3����Z_z�R�R�|����	�[��R�{`b�C��߰/'h�������������}4?��	�QCw.��sN�y4ᬸ�p_�O�	����'FX)����1� ��:�h�3S����3?=����Φ/�z�xM���_��{�XtS����r�v3ki��~8�8JL�j瘂p���jo�����V��2�D`�X/����c䰔6���B����S�C��H8%i��:g�dA���u�f1����ܡ�sP�5Q��8�0�m౓N��r��~anA�~Q�4��,�=.P�YL�kz
�B�u��h�~\���n(�+�����Oq��b���1A�!�r��q����!b��h�����4g��A�i��sz��u�i���f�����Z|z� ����'f"=�.��,P�ȇ�:>4�؎2R�ac�>�鴲d�7H�NEH[�ix�S��\#�����[����X	E�>[����!A�C���8kyʫ'����(%B�����CΒE���:�����x�X��b!!�� jJ�T�}�wg��g��K�d���9?YG�Nϝ�� �(�{���~xT�I�?fvn�&<R��Gn߄� /D�h��ΐ�I��@����:��s�Q�zXV���
�t�T�請�\��<`E�	EÁ��9��IE�0����m�~ڗ�	 �_-B��~+}Čcv�`�8�@���c<�,0�����º'T�y���~�H+�9!XDy#G�t@A�z�=q]SaB��~���ۮĝ���܅�0P�J�RO�k��}��C��)��Ԓp�ɫV7fH1S<s�h�S'Qo��D$�!^�.��Q��Z^q*���hg��pQ��M�e��4!�����3l&�[�	��@�<F���L��&�����`�7�\������iѝ�A�����|�L�
�2K�
�d�v[����|����=D��ᄠ�b,�PU�xO�zz>�`���a�:hd D���|���󸤖�#�I�:4]>�哶��4��t��xa�C@�;�'*W�0���!���\�s������s��1�~Y��c�x,P�t�7�u��R�z����������  bcr�0�^��ؓR 4�|O�7��<2���!$�~�	�il�ZzI*���x���
�ԯ���%�(�ފ��*S��bކ���_ڮzk��]�[[����:�TXr�1d��8�t��'��HXK����?�/�uUח�y@ށz��B��ף�E��z&��ݜG��b�M7�>)������9#�WKC��T*9>ڦ��r(�xt@�c�|Kɤ��F'���=TT�
��� Y��}�؍jp(teN1��_޺x��
�����&��#` _��q$/c��Nv�����:ͱ�Mȹ\Jߑ�"�z�]S�`�r�PP�;����W:'6��0�U�������# k��Q5�D][c�#V�DJLu|4�S0ԋL	C��	�_	OB���%>jfar�ELڍ�6:ǖ���d�P���I�(}����3W�H����ӊ�����ڥsG1aQ��G�$�0o���'�����&�=��iJ��f��ar%�x�W�y�c�<��Ս\]j�\M}�=�J��!����s���T��T���i���(���n_L�R���������E\=
����Xi5�Ye ��D@Kb9�#o7 ��a� Y;�3[��=�s$�>����V��S�P�����Z��R�����=Y/�zl�;�60�,��<�����pm}6Q���if**�_����CF���w�X��\Z��(f.l�Uz �!|~r�Y�������V}4p�~������/Q�����7�d�4Վ;�'�ݷ�}�I���6<�V�����y����Co�;@5v�ֽ��k[���Z!X��HQW P1>%�w4�(I�#�E#R�v��F�v��K�#>/XY^IW	�t��Z�jb�~l5���Ӭnb��)���]��5l�]��k�e��gyd��mN���,�!�<ċ�0[=(ى�����h�{���he&C#͙oט�^?)����yLB���t����ƸB��=5�]��
���1&.-��i�[oU�	�^�c$�v6"w�3������������b[B�fM�DѮ*�ir����4��[~N�a��G��{c���B�&�x����DkU��\*�g���4|]����x�O�`��)�EiK�|�8
���Ǟd[���nH��E��6��~��<(��?��f���f�};���i�DKfh��e�Fw���f�Dg����bysȨ3��>�T ދ�n�*�8ﮓ�'���33(�I3���T�"EW�{(_��Z��׾���n��q��"�_J��t����
�j�1�����ޛ��x�G���w���M��}_E��
˶6�߯��C�J�πy�/ �S�]��ڙ?{�N�<��|8v�	;-VH��C�-�zC�n��B1�����o�i ��x��L�8Ȁ8���+�=�����j%�3��즯���r����F� ���4gu��qS"��LQ���Ҵz�8k 	��e����`�6�˨�w�����|{�^.,�b<vfq��GF�|�Ȭ/�5T��I�<-[�p�w�{�S��xD��t^���Հ����
҄��eZ(�럐�9R��ka�c�?���aQ�-xS �ˍ�f��G�t��� ��E4'&�kH��(+g�t�]ҏ��t/�����<<@W:(�)����y��mmB.�"�&�`-6�V�N�COɍ��z���`�Jo���ɡ�	*���дaZk>DZLA���M�k���盯�]a��#�{�'+�ɴ34��u*��ˋ2U�k�������#�-�aPi�H�Q��>|c2	zL��A��c�0K|<�Hx�A5��jL�����J��l�ٲ�V�V?�H �Y�a����\p�d���%����R��ʤ4��|��{�%���ץ�Y�(e��(t~"�T��#77�TnS�Ћ��g�p������VFt���[����q杽�"<h�� �ku��H7hw�T�S������eH�Atx��45 ��P��$�Ii	e�'ӟW�P)
���:�)1$%��G��� !�.��Vq<S�N����M@��V��إ��&�c]P�����C8Q���ˍ�e�V��O�zV����d�T�b�(��`6m�"y"/���w�ڏ(�ɚr:�Xc�i�c�u@��f���ۙf�}�-�ů���[����R���5:�����Δ5|Jf�,�co~����9��g�n�or�����İ�"eV�ǜ�8��	�9t|�;!nlK�C�Vۑ�%���b-ow������Y�����MBp��d2A;� �I׬E�#'��D�k�x�nh�� -&�M�f{w�Y;���RP�n���١�/��,}6x�B�G��J.� ws�NO]�Y��^�������ǾU^�#B�ݾ]�9��_�\7_h6�;�>Wzޞ�8�F%xLE�V�d=6�WL�m+�b��h�'n}���!Bt��cKi�Z=���R�g6�y9�ضo;jl7��?»�}&:M�)ǅ�jщ�����8�Φ�à+K
���J�7o�&2�vѨ(!V��.����c�/�U�S��[:�y��Э��w}b2�
�/�/�L�(��L��N�v��>^�"���c�\�Y�8�W��&�-��6��m���0r�������.�v��\�XT�6�K;#�os��]�k���Vh'�5��,qk�i�ٹ��(�2�b�
�bQ���'!� (���M�|>ɥ�A���Z��c�g*�z���������1k�#~!S�˧�~8h�
jԒ�ݑ#e�m�w ��+]�V�(�ľ.�WZ�0�$���"P}���ݟ�kt������
C�э\�JE5bsH�XJ��6E���-�z��9	[&Y���N�
��wg���y�;��
�V��׿N��<�.J�t��X��\�9Η�-�|*ͬ�`m+42ֈ��X�N9)C<���u|��PoBo�qʽ0��_N���\�-%R�	��t�ɘ�ߌ��?��x6wAJ	����B_#�K��N�զḄJR�"��`�+.}��<k���v1׈��Uc&�v{���v��)�L-�#��9�:WU�Z����Z��[f��R��6�'�@�z�"KZfE�ګL�W�h.�&b7 �P��!�e���, �:�xp�XcO ���b��R�/b{Y�����r�Y��F�|8��*[��h��8������	�P���(��=Ы��l�g��+>�+.�b��F�-fX�ȵ�OM>�ԕ?ܦ�ډ@Ƿ�e���$�� �:�}0�V*����Ǝ{/9g���<�?���c��a�6�g�%���W�EY�
<,��LK�lB?AkPZE��ˬa#	�
(/=͍cɚAQ!�O�N7꼢��W�(����lydB�pkܿ;P�E��)��~o�:��PxĦd��L7&��b;H�˓��\_�oWCY��H���Ԍ��$�.�GQ����ٗ��?ܞGP7���h�T�@�n�̕�e�vD�t������D9]��3lwA��us��QM%꬘��+�5�jW�1���b�&�FB:����U���{|np�]�e�7��ǜ����|��*�e[�yOD^��X%�J��a^P���F�h3���=/V�f�4"ߏu�^�3e�=t9(�?�<[�5Ba4�<X����|`(�"��;Ju%]�oh�B�kX�Q�(�����[�+��(�.��%���"�����0rp��짩6D�}��KX��;��#�� Cϭ]���D-��$��{�sw���~���y(�vj��x���G�wlDm��'���j���o�Nw�~��>(����b�E]q`��?n�w�]����.p����8zy,z�hN�T�_�br��Z4�
�E�c��
^|[�X|���T��nn�\��M$�x���_*�JlN��רD�y��>���Rys�BTy'g��{?]��j��@���/}�l��F�L��kFv�w$�`_X��
G��M��o0���f��^@��\��E���4Y'Ā�ve�B1z��VIf(}�74�*5G�m#K�$���B9�պoD86v�Z�;ہ(Y�D/��Z��)�����bH]n�}��P����)�_��JF<f�&����Z�]���^���N�d�6(���{���"���=��/!4�ppV���bg�]Ho�ۅ��U��˫r���W�:�n�[�,����y��"�֎�������t+o�GE)��*{���U@]~,Q@@�~F�
�N����gU���Ʒ@j�l���5o9/��Z`�|�m�*şŋ�qL�-�fݥ�?e���]�ԧ��������R>{αbX҄��[1��Ux�'���\��*��\�a�ֿ�£�e�H���a%3p�/?Sh,DrcvL~��毇��^ w�rc٭v
�ZR S�X�-��O�R@B�j�XO��T��8�:�g:U�>��}��ÝϣFB���&v_"�.�yj0w����p���u�^,n��W�w�5��N��j@?)��ϡMڻd���*�J��-��z�S�k��c��߅F�-�j��:�<hY���[�\T{�����&��>s���_'J?�W�bQ1��ȅ(��0��KY�!�K?\��$����xM��nº ¦�@q��3�Vtn�U�x�pō��`�dB�{fx�V{+��JjlؓR:�Ԝ�^� ��k4��#�'p5b.��8�$����C�)���ĊP(?����@_$'���k�5"I�?�҆<��N����Μ�*���#1������� ���E��I�h�h�t5T�3��9%���k5|j��]{8G�ܐg��!��*]�Wy_������×[޷��Z6P��a�q0����5���ip!�s\�6�`��8�v�����w�����ڊ�傸�������,'�t�Y��|m���`�Y��2�]}Q)4���.�n؟Z�z�����N��#<L���M���O�����������]7S-��F�;���,�u�l�<�5u	o�l\
r�ɜv������p�+J�
�g+ze�n���=�H�s"=�n*���:�:�@c,5�R�9���� ֳY��g��J�t_Y�Lc��30?\f����1s�myp��*j�(�%D�w�:^M��0Յ��-���B?4�N��p��e�0���fh���);c��4�[`�Ŝ�8�,Q��7����$a���!@I����swS91 hЕ����D�R ���nb'�f��S7��{��ݾLo�ᛀM���foh�f���dUe�Bx�ߠ�qu��=oy>�D{C�DҤAS��H���y�¸�����2����_E{{F�X4Mi�b����TQ�OP�E�,F�6�+�)G@�����4�3��H���"/n�]��B�;�I�X�����M5���~P�%�P�S��;"�H�����f�(lD��?#y"�c��ğ���F�醹�!T�Q+�lq/���XqP*!���7Ӝ���ơ���T�.|Ϡ�f�aD��iV�R��Sw���ڂ{8(��q>ֵ��~�٦#�deZ�4d���r9U���;{Ԋ8P�N'����5>��`�A5Z� -�돦8��+�Xɧr�u�6:����T�{�S�tLҚL���C�Ƒ@c���L�� +�����&pW	�W���(��se=\S<�`O4�X)?a�~�ƅ��N<�H@��t��I"����m8���r49�Ty�'CB��Eha*��0NZ��Vj��L�����(9ZU)L�aX��P�	��b���aw��ԧ�b��$�>�췚|�C	�Dj�4��; �:E����zt'ޱՎ��zgC���`fl�-L�~}'�����} Y�B
Ag3�_�?�k7b>X���gc�Y�F�;D���s�y_:��by��'�Ȳ�.�P���D��a�~�2+J�&i 	BX�*�T��HJt�2����Io3��h�ڀ�.Y���8�yN�pej�xc%���'��`k����9�%�ZO�1��4o�c��6ޕ���f��呋Df&�� 2��qMo�'�{M��%Tg�ohr���b���NޓI�=��0U.|�S�Z����,D'��s��l_��	k����N�q4Zv��t~ݍ�R�F�����=!�_́�ux� �����!U��;Q��t�H�H�@�S��4io%�E��T�m�)
�xhfɢ��eA�8_ֳ�{�.� 5t�bVG�!��D-�c�9OƴZ2іq�d4�S1~���>0~=����^Q�O̸�.����3��~��״�b��2M�	�؏n��8�I
��¿�g�qyc��$�/�Z�e�8=|��R:��gv�{���;�F�^])BAO9Xfz��DI��}��)1e�o�9~b�M)Y�,����,�_d�?���|[U��Rҋ��ň1RgZ��Hv*�CUGL����ڒ�����He3oLR�NI5�����y����������*�a[�����s7痦OU^4\^:�Vk�sg�{�]v�?��/��Wx�=Om�q���?��*���/~񭟯h��b�j����(��C�T릝ԉQY�*��LL�
��bLh���p�����LN�m�'��$S^ϯ.z�����3̾,#���<,a�F'Z�?�R�$Z��w��٣�Rs�)��� �����Bb[�����<ZO�)-;���V���(�*��b�F
p�M���W�\�%��w�,I_,��lY�+�9-�0�3;�(�p���Fr�C���ϭ]a���2�lkV���gȂ�74�b��twOTi�����ZeL1v�B��KԜ��~V�w��(��H����
4��7��0��Ãa��׆��9�S�֖���2��0)�-�i����Q�B�%QC�c�j��H�%wOt
�N҆�X s��N�,�4fx��>�58g�
VZ�36s��⑨�Y,Ʉy��(�0yp5� �#88Â%��;ƍk�<������E��_\�^w��<�G\��=/z� Ma����}��E[�s�%0L�H7���Z�VY��3�S��C��׶4\�������� ���q�/�2�v���B�:�LV���6��H8>� �,1΅�k�Zܽ=�(pL��Q#��_rÅ����/�̌/�>fӣCVc�|��!Rk�M�FA��Li��<�4�@����_q����h7̨�W ؆n rN� �Gyp���M[�mR�	�M����e� |2�0��D�r��b-�����S��O�w]]�~��cU�C�n;�p�75�����昵��@��%V�o��gu��m��u7s��y.s_�Jy��8��}\FM%E� ��(J&��� ǿ���3�VG��U�l�,��%��C]q�{�BX����+Pk��.8�c·1�U0N�ٚ���o��dl�Փ��㞂�0�xy:�P�=�=˺�E�/�|/�*ڱ��*(��>+&�d�`�-2��}}�e̲F���7��"!��� �fam��38�j �Z#�e>峁����)W1�����a@!�D��-�8�)C&�z�bxҾ'̲��"?�/M�A|h�#h�۲���n��k�!��i��5d�ﯛ���O&c�%}a:���י�n,�>�:��s��Ν$B�۞�2N�����z��Y�_x��
2��("�:W�����K34����w�?���g�#�����7'pJp�ot0�f�|����c!��ڢBdL�׽�m�P�!1��r�Z��_Λ1�ǔF�j6\|����(�,�f������i�#�G��[�ד�70"/|�䭗�d�@�2��-��#�F����
ZF�=p��P��剸l�u�AE�a����%�]AjpkC�EN�̀�i�|p?�q��|�rc.�k���r���2��R��-%"!B;p�=~�D`����Ϝ�<�a?!�#����#*®w���t䳘��I�l�_�0}9�m���,�B�U��N1\�]�`zT ����7�xu�޺�
u�ʪ������:�oP@2��J��`A���3G�_u��(��Mφ69³�f�k�硆F(yo|�Y!��������Ad�2'�V���+-��%R	�a�xǒ�4�e�^6�~ �|~KR�Ci�i@�d��:��B����
FFs'��:�6���,�)6�-%+}�ZH��p�>��;�gc
r<v�j����(�l���{�L)sr>|��=M���{���Cu�<��	�ߣN%��č������<�uD��.�'�Z��w��}-�MT��q�9*e������].P�e�BB{;�P�7n>T}��rc��j�7�O5�
�=�T�!z w���	e�)���D���#��v�^!��L�{���YZ(�O�;XR���%���D�?�u'�I��y�K?�Z$Ji�6ОZZC�\������� R-z�rd��|����>ޔ�&��\U�� -W�T�#j��-�
}8�7��%͓��Hz;���3�PVP�{����1(}��������mfQ\����ðv	��)_�m���cՠY�
���~�PY$n�;�"���0V���]0��0���'�P�&7�ezp�
���A��@����T��;C���9q�6331�]]���q�z�w���q|gF>�CQr��I�I8��2s#'�[�.6&_� K�߁��:;>�Ƣ�o��+���xfz�:�̧�Ѝ^�t�4�h��h�Մf�?5��T!��z��D����Q�*�����C^�4#�q����qrY����,	��A�ˡ�}Ct���-�u�_�� ��!=]��+�m>�� ��=s6�T�uM;p����D5.`�M����l�Q�TR8�L���Z'����f��_۽�l�O����k����'����XӲ���L2���&4�yn���ˇg�ΐbJ7��x��x�B+��:�!�W���;ס��p]�S�_��e
?��<��>�iUs? C?���rM�ڌh��5���]1
M�DY�"��N.�)I��nפ`� %w��~���ָ��l/2�\�L.� ��oƣG������Im=���ӁH�?�^��N�F�y�
��N�-��ڠ�y�m)5=Ԙ�@t�̓L+J$w������\��m�$@��#rЮn���y���~ �G�AN>����,�Fo%_��j9ķ�>�g�ZVY�o�|W7p�ŉ ��ze\s�-��V(��Xk�"�>��`���xTO܊D��S�0�)t���.�9;�*X��nh`�8&O����~1�����;�\nM�NK%X�^�(T���Wy��Y��i��ɪ.@�;���Ec٨�M�l�] �{K�lLa@ ��(�m`:�q�1as�(wQ����ܷ�FV=pX���rS����1hU޲�ɚ�kc������P�=.�1VN��=1U�V���N3���*�_1��\E��c7ci;Q�LI~�l"s��ئ]3�����Z#�{,F �?����RMe����7!ߓ_S������ߚ�r����N�k��DCjp�p���^
��6?�?)g��;/T�T@����$'�Ğ��+��|s��9���8+_L�.1؃k�����/��-�*�F��\fAָ����]��|�G�]n�'�^GGV��m�ץ;� W�	�(�*�A;ŕn���R"~K��	�WEr�p-	O���#A�Ø�������m6��Z+�C�� D�kZaȹ�t�J�^[S@�	��aw*��6H�JZlG������ �K�;��B�pDI� ?�Ms����Y�"[�uZ'��b_�Ipܽl��j�rKV ��������$R�_���ǯ�l�.kF\Y�M�!!��y_��*��T��fu���mQm�̯�?[���6i>�_�FL��<AԄ�NXg}��,�r�,��b@3r�|�L��f ���Q��&LG���
?��h�o
X�nv���f��>�l�$��5��-��I�!ۑr5���1���h�t韠;���6�63�;Q�V	���k-S���pqR-��x�Y>��Y<5�,Ԇ>%��0��Qs�D�؟��k�z�����2z=�%_��Xn��ye�fV]-f�U�e<��nސ�w�.;aH�7��=��by>V��4Q�SR�}��Ŗs[/��7�x���px��!9�#~z�K�e�*J N��{d����H�{�գ؉Aus9g;��ײtZ�P�����7�u�������6��:�V7p��G����7F"��PjIf�=jkX/9�A�Zќ�<�z�����2<fa-Y��#'��_�l��Πn2Ǟ=� T�-��Av��/j�M�vm��XE��.+�k���Lߟ|��,�Ԛ=R|2��Ce�V�l]� ���o�1S1�2�׈#����F6�f"D�͎n>�8o�:��/{4jkm�U�Zo���Y�BI�l��̆KG`����)�y�ɕ��9a��$��^ ��� ����`��?#k�u%R�L��aD�jK�D�A/��~�Yb0kk��n4�S~�><:��`Q�Z�T�1�vF8���T/�D��V�#�6�gW�<��#v���d�V�����)��a[�j_R�E;v:b-�"������4Z�^s��J�_�=�q�ﳦ�M� ��U�!7�h�JN�*������2v�1]b��WD>�ۣV��mrj2�L��	M���
�V#S�U)��i���ni	 ~r.�CcP����NL�U�w��v9�ә)+"�}򦉿�[�OuY�h_!�Y�=�d�����$i�.![R�e�0����P_��{��k�T�OQZ>/r7$�u-�J+���!���X58f���1�~~�� �lV.\�Si"�t���x� ���}�ځٜ̌IK�1H�V(Ⓑ^f�����u�I�zB- ��ŵ�PGoE5����SAmjF�U\�+�A�nJR��5�̡�\f�lO�a�9.����� jaR���c]��0����R�ϑ�LI����#ڽ"1�EX����pe�l����(8�-��Tz�^�� ��1��)�޻�ã�?U�rs2!�W#o�NV�K��!|E�t�=i�ua�2&WJ���8e^	l�d�A��F��x�0�A������k�y�����d������[pBL�3���k�`!3�l{�s��A�Z���?v��0�b�@$9�/�RB���q!����J'[5��"��3E:c��%�A����Ч¦ⷳP������E�7�+o�VKw�t��+3���2vaUL��{w�z�|K��@n�H@T�h�N��a�	��b�;�Ӌ~�a.�|ζ��v/�!�)��R�dv�u'���߭��j�L���ֻah��K�XmH�cRȥ����r����nE�!�IXf�'K���g�H�M������g�*:��Z`�\��ab�'��v��w���Ó�9��鐉Ï��϶�ET�\�@�[�7)`Q~�W�'�O����t�·��w�z͹'�U3$�(fG]�|�L�������$�Ջ���X�y;��|��:)Y���O�f�y��`��ZR�X�f+�$)q��E:�?��
z�\"�\��ۀ3�l+��A4Jc�T�V���6;��p�e��2���9m�jwV��Ā��vثi������$������G�R.,i�^��|9�iUF+`��0%���<�M;��){��	o���8���.!C�/"�l�GK� j�<�)(��{�'�'����x0���E&�o���;���2��E}�s���*�[%�KYjjݖ��`��-�t(Eq��x�L���H����6c����hbݥ������"�c��=�O��L-��K86����hH��G��R��68�G9�-���IJ�"&'������Șڄ���.�4@֒�8���T�W�����>��lߍ���N`ß�ڇY�����:��8��#�o��
���5Q���V�1n��<��h�Zl������J ��Nʎ�8A��������{4�mD��6�Q�a5䆔R�5{��w�w���+D��ƾ�k-	��p����� ~�j+a��{E�?� ��p���!��vL{�w	�O#r=�*�0�����B�ΎWw��ەP��P�0�=-q���$�C�oF��m%���o��%G�*�� ���>���x�����Y���_�Ә=8Wзw�p��0�3D�l��6�}�
�#۲1����B��.�p���W�W�C독�b�J�J�	+^V���q��� ��o��.�e658��zd1�;3�v��1䀸E1����/ϕ�^�P�*9׵ݺ�6��P�E詒S����7���&�i;c�_?��$���X��4!g�j��� �(�VR��H�mUo4�95�7D(��^=^V3{�B2���1RlR�=s�@���R�A����ャ(�nm5��-$C�P�@uJ����q#�=ze�厏n��[��R{j�+�,�O8d�������B��X���O�G%�I9=���Z~ :2��.v��g�s!�禬k�C?��%�:�;� ��Y$�.~��@ycNἠ�qc�������$$5����2��;>��l|nt����o���jr[I9�d��bj6B|t�a��#�A�OLZ�|�0�yٕ-$*ږ&�Q�2���q
o`&"�8�Q��&u�C����,��l<��D��DFD��I/�(4N���?��2�,����P"X�`Pu���G���.�%%v�y�d)X[��.����/�s{�q�I[$=�Un*��(a�F!`zE�{P{Q�����F8wWdR�ge+!킸�+lz8YN��QÀ]��>I����%�D��;�w�i)�`[�/��7�G}J=�l�%sJ ���8�]I%.���bC�d6 }'np@NZrB���f'в��LS���5J�����Nf@-Y�#1r�*"9���/A���@f$i/ؼH���Wl#j�[�0PiY�R$E�6B����\�p��N�A%�8ӭ�|O4ӟ�F)yEO�[D|�S�� ��]Q�M;L��#&IUg0ÓJ��p���`^�02J��}�e 3�߿x,,A��p��V[@�X��9uJ֓-�@3yӎRm��&�(�'Ț�h$3�k�rG��3)��d�i �.��;.C���Π���̘�L��N�?<�ɰ��?�+��1�m��F�f��gڊ �Q�K�����tl�#w3,}=�I�&Z5Ef��v��D���`���O���i� :�i#&�8���'8��Z�������(՜��~�=��@��p�?��V�\�J��ʑAH�j��Z���~��B��$��7$|]��at��,�1�t+�\T���^X�3j7P�aq��9��uC�2����5�-�����myW䲹��s���ʚ�((��ԩEU>yV����F����H��A�Wd�r?!5�J�z�2�=g
�wσ��ܧ�j>CN�
l�(F��3�s"�M��d��t���d�[�N�N}�$��ZZ���Q!�߯O[T[��9�5}��j�)eT]��}nf�������2I�f��:,4���p5W��)��W�x/��8�B�B���#l�xhj��E�"OH˝�oQg�M�D0%V��[��Ľ4Ƽ���,Dz+�a��9xɆ\�51�'2���m��o@o�{�z��4fcko��ЌF���Pϔ����i�B�i�!A)aˏ:�`��7�!�-�+K���ȵuh����+�C檖�IX�If�`)�V��sy P]�&8hý�r5��ma���&H�!"Ř�S��I�o��ꖻ�-կI�o*HGH���m���ԥ��ÚjtK7Q�2�����'�x�7J%u����|�/ֱ ����[�SG�3�%bb�Q� 	�㣈�T�Ôː���^p|�W�
o�IJ�>���pR�y�f�#�q1��3��bh�4�1$�$���($�N�o��[3�$�0hT�{^ɖ�q���:z��|�a���	�
�vL0KPS��,,�~l�f�]��,r�پ�w�f��+���qf�m)��Z|��\�uQu0�M�r�52DL�������y�k4����_�n#_-�	�rPB���=�2��ʂ7���.��T7"v�u�i!�y��gI v����H�/��X�N3iwOm�O1ƼM���5�k�'��?�i`C�|�p�ʯ�?�3�M�/۬)`pl��M�<7M��P�ʠO�?�5o�/on5�n�孩<I@���Ѣo��F��3F���F��4NR?3��h����%'���Aj��+M��8��6�ͯ�7$���f�B�.�A\�1��Nth�[/,g�ѰY�����5@�:R���j����ըB��@hm����a�����O�Z���B����#Gw \m�W����FGpñC��Hpw��/~�PNM�yRX�}�eZM��?p�G˷X��ܡ�頙=�}t7�Wo������ד���x��+�:!�)0i��;fϕn���)Rc�@߱��i�[�e��m.�9&)�w���o����h)\����{�kɉ-͡(�〚�l�������ث��ُ@F�"�[�7��X�"��ʢX9� ���o�NSy��KwQ��V����Z�j��b��`㾃t��m�t�i4�+����w�rY-k���~:��^�w�J��n�Q�>�O�P�@�C�-!Q����[���q�%Kc�k>�5��9��7����v�g�*'H�ק�7z��|�J�-��l,i��KJ���ڮ�������(^|����|��TL�I���G�bf�#QY*�{�a0��E��&%�X�~BMEZl06�;>3{~����H�U�h1}|;���i�0�&څ:�Ǿ_��8�����;�a���K�*����޴ݗ6��Vش�D��q�`�MݗJ��{F�r��#��H���q�
7�t��lT>������+p˰�[��R̖�8�O��'	w����^��׆W���}��s���0�k����E���&-��S(����ʒ�eH���Km'����.�{UuwՉu�$R�����O��X%hv]^ �˗�9pJ1<�N�!?�ޞ��=R����X���H�