��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+~����S����rGq��%qULpz�XU&JF���a �/=��Th��e4��U0���B�4f��zG�`F"p[G�~�z�\�M�)-P= )[�ƶ|�?6���e�9Ue��Dt��E	��P�/ �N\��e��{�2Wm����v�}�r�;k���g���o�*��<Pkb~q�'��[������n��*HǞz�A�2��˿h8�:����'/Rܶ������g��}є���%�D[f9����<����\Q��,ڗxԡ��x�9�ˮ�nvї|��#n��J�}��
5LR���=|�v�=C:����:d�Ŵ���/0�F<�Z���粣� !�MYbH��g��恃i��W<k���a&�qU�3����.���ٙ�,dؼY��lGHزJ�-���M��Q!մ�q���9�w�r�GC��R�A����~�!
���_hՖ����I����6WR���έ�c��� 2��(����U������C�T���CSl�SQVM����}}Z�)������X����l��
�JpG�JT�,V�P2d2��ez��.r�Asu�rsA^᥿��ص> '��5�%���x�ґ�S+�v���0Rj��.}tс6��SH<8�6���.^G老��R���E���͜���{Es�2�PQ<�p+��r����{�����v��Cc�\u~��J�����-��#ܗo��,�`���í3}\��J�Ã;<*���I��k<=M�"�2iH�,���O���埌\�6���P�����o"
���5:�sfV	����ۨ�o�����YI�+��L鐊�y��aj�A���bRxM>w����ӌ8>�`y�I<��N����B��Ǖ����!~�=����Y�u��g��\���j�R� v���磃p%��%	-�+�{��2Y���#Җ��-�2��v���-	,�����
x] ;�h���RlڭI���0�SH˻�od���Ҧ��;�&��1=�4�s������`]�Q���"<�S��;�6�E���T �qJ/o:�yjz�mY�!\���Е)� d#�F�J�zu�O� ����cM���I^"^\��y�p�cD����; |.3�	�.��P}�<�n����!B�O��IJ�W���HA���Y�p�}�H��KKH
��h��"��&�J49!tp7��(Fҁ�gD{�K��7b��?>�<��&�pͻ5�5^��t��TD�q��b��|�җ��`2k8�"�Nf ܛ�&�'{��Q]� nBy�Yֆ�]�i������|�p�}ln�>!+�X/�b�q���jA�,qaW�<?J�]�&F9|xlR�@X9�Ֆp�;�jGЫMo�h���()�m=@"ya�A�˺+�n����M����zI�@� \aʰ08������L�2����Fıx�����_;������;�N���V\vr�+�.~��A�vV�>sk�f��(l�%�5�g(�]1�%G�Ȥ�V�}N�>Yy 5�ڼ+�]��s)-���2|*�/{w����	�QO�xD���c3e�ְ��_�O���[����x�}�$��ʻ��\'_^;LRd���o�C����Ip�r;����EU�K�����Ixy�7ܸ��0��4�����v�T�������˶p��TK��Q��h�������._}�<$�#����f ����4�Vf���ғq&��e ��:���?�����
p��h���JQ����B<ʶ�����x����Ŕm�]f���*�Sac��3HĪ�X&]2[��p��"�'H�xʹ-y�^��IA6�*0'ț��+g[Ѯ!�{IGe�Qiua��[f|�e2�:�zw�n��	 �|>�2s92��=G�R ���P�d�}�%R["��s%21D��Ď�΢��-#�XZ�	l� � ����P��������z�j��#6Q-��;��5ǇS(�k_+FW��{�T�W
5�IxvoAƐ���տ��9X+�	���;Զs�wOG��A��f�s�5����Bѵ�����ӇRhA��q�~^hLr�B=9��^Md [A$�G��)�/�,��bl�je���7O��w �x9�l�[�ȟ�;+?���l���[p|���z�p(�QV�s�f�yE�;D