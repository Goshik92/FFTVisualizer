��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_����m�e"kxu�Uٲ"#oB2�-g�j��h�p� M T�(�P�+M��&�[���+~����S����rGq��%qULpz�XU&JF���a �/=��Th��e4��U0���B�4f��zG�`F"p[G�~�z�\�M�)-P= )[�ƶ|�?6���e�9Ue��Dt��E	��P�/ �N\�$5NB=_i�O�Iוo>b�i+�5�s���o#۩[�?�q������4�t���(��ִ�jb9��8�����O�Rd�*���E�*	�,Z��{�m��m��$��Y��dWB&j.(K�fI��3d�j$h�i�g�����������U���i��jm�5�+v[�(��pȅ����kC�O�yъ�	X�]��g�W׫Gu�a�Fʛj��'��j�^�q?0��y>q^=���kb��`�H����8N�	��G����q��N�L��܏"��Q�㡫��:��ߜ��z}}�p�U¯�C+�?"O��Ed*Ǹ-7 Q�n~��x�M���� 6��!��� 0!2]�-��EU�Y8�����%�u��.c�Pp~]�A����Y�I�ڒ§e��Z��%��4`읥:]�6�N%je�����v���Ǎo �?��ueRC0�3��"��kW.�Q�_f�^2d���ޙ�`��IF���*Q ��|�D4�&��%���Tb�%����͘9�����?��$�!
D�k�H�^�t{Z&D}�E�-��`�$��)6f|��:��
 ��3"��(�����g_��W�����P|����P�L���.
6l�B�r�i꠼�f���k�����ot�Z���CP�b�¼���à��H���Z�w�j^l.M�5AnT��]�B��]��h�,��u}>ٔ�R��ེ3����:�G�o���3��;����!?������):��[Z/�����pOb,���w֢_l%����E���	�v��Vԫl��*ƼEsHEZt�	6� ���(�����8�RS��"ӻ�R?�0Q�������#���J!��<T}�|g
�|`r���	��ۇ�eB�>��&�.]�J½�e��4/�uz���fk8)շ�N�����+�.��r
n"m�?���in�R���,�.c
���:��{S<��K+�$�;��|� H'"��z6&��2�~-?N��03k�fg%�
�6�o����G�,(���;��we}�,#pK��ܩ���[y��f5��c�l����/�s~ۿ�I��\�iL��c�=�X�,�n����=�8�J��ZX/�2��GD�&�VV���x�t+�Xc�0���=m�����<jJ�O;���f���������-eT����抢�}7���FK�������e�8�����h�ݸ+�}�!��:4*�Um�Lz4�p,RA�/w�޲>�Ts�?Kӿ~�-b��i[��Fl+�_��$\��L�f�Mi�8?\�p`�ǀ�� ;-	ܹ�ԣj}ѧ�3���y�_��,mڪ*�_�OC?̘遵O��hL�#Κ�H^��|�7aS[�ۊ�~�h����L�r��_�	 �Ø��l�X"��!Ĺ��覘���w��l���d�p�LvR����6�͚�2��/?�KdJ.�XW:_�F9��U͠�^?��*��w����u2����7B��^-�V]��3M�C4�P�h
<YD�f=h���i1���_6/]C0���x��O���S��!ºF�	�j�`��N|^���L6�d)  �(�����a�Ku�����J& ���C��m��Z��c	=n��w�1,�Q�V���-�n�m���1�X#C���tR��g%��a��iՏR/����ٖ��|���~�)�eMۯ&JN��M<�hT�#،�k�r��i_�{�XF	3� �^�U�*���p��R�E�{QT���Y��Z�x��1x)��x�����/UbɂC�Û�@�t�\�rKH;����2$��g�k�u��W4k+��_7�Ԟ��ׇ60|x�'�WE�z/�>�Xl�m(�;"ʟ��l<��@$�6?��V��uÎ���%��B�ElV�;�@�N�2eFڀ\-:ժ�8�ɅKS��٣`�Yy��1Zhh��Cd4�x|�G6��Ě�E/�B]�e���-���ܓ�����s;�!�2hE�_Ѣs\5�Ԑ�[o$}'���=t.pʏ����(�%�D��	�軣��y��dc-��#��cՠ��� ��@*��LgOю����|�>\0�@�:��(� ��(K�V���ɝ!syr����B���}���U=graVT;���kR'Cg���HF���;��j��#teBKg�{h�>�*�����V�鹟6Y�%0��>��H��|y���"'�+L �丗�4�AX��C����X�8U�����p�g�M��\�_����v�����M��8G.�N�v.,��5�M����/�?5�M�!���[��AU5�^��b%�4��0�'��[�گ`�=|�ib��m���S�4.�#��PU�j��Q��ǔ���l%i���-�<#�7	}ԏR�:5��U�M��:��t���xҨ�a��.��j('']�-v�V&��b�o�Y��̭�)�5e��s�C[���%%o1&��h���;_}G&6��>��W��ˡm��Z�	����������ߧwG���r.L�N� Yk-���Nv���eT�a�R8�6DnLM<�`�iVX�	&���C="�{�9b<!�;ǽU�E�i�Jz"= ��#f��9,J�~�Q Z/·���