��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�c�z���-(qC��c�諀2���RF�!'�AǱf���8)�}Y�J���H[���ժ���^��m�&3��L!��wIm��_�#�k;��� !@yOcwz��^D5�)�Y��fr�C�u�7Ʀ����<�ڇ�k�7W��"	���a�:��9HLo��F����"z��!��h�쵤,��u#?y��`�W��3��N����\x���N�#n��>ޑ{��+�33=*�5����z�7�D<I�(9rG�ﳄL���Fa� (Zү��\ȡ�n�I�����=�vvHh�\7hZ�P������'�v��;�ULJ� �n|�0)�|�H�$ԍ�a����V_$A���9 �C c0��J~���)�#�[Ma�nĴ-W�p	h٭��I?��ڊ�[�������=��bHE�Q��'��D�A��ʤAB��>{'.�
N�3Ǜ:,��+ *���~����nޔ��;�M���V�),|�q����{����P��T� y���pI�������|�Z7=�-�4y,��X�s@�7��/~BL
`��`|� �Y���;O�q�Y5�x՘�[/G��=ؼ��wP\��X�O��p)�N�]�=��+�*`���39r2�����KKX���,ŉG��V�_ �_)e��!	u�����Utu��8[���]��_�l��F���:��]��W�@�C=�%�K[��_^���j��>�vX+L�,�
�����m��?�+}�2R�S�}�{�#��%��8Xş���	u���O���&��@��m�-d���(�"��ԯf����x�ƌ�]/�7q6ut�-�O��V	�b��KcC���f��\�O�?��C�p��cr����0�h�������Y��r�Ho��[U>X�ao8�OY�y��ya�J�P���s���Ⓦ�w��99��)T��z��Oؓ������Ё���,bwN�%�R�I&T��鵺�V�b�#����_�ՋĂy��=K U�խ; z6�~��A�pA��a޶�%<S��Z�ѽN��E�C�rA�ܴ���-�VY�m��k��&8J�ʲq�.�a�mg�O5�W-���Sq�҄��C*Ǟ�D:@��?4t�|��NV�d� �6�ݒ Fz�^�1��P���>H �+`��ݣ�F	T�:�&\i�u�EJQ�d��^�]�H�' 0�ȳ����vN��@���d��vV�#�yR#\���?4�K��պd.�	̬~z��^�ovM�u|�k��V�-HHF����:�c��D4�����b�Jl�IEVy/��ۅ�U����/���k��'���l�m��땝�W6˕cO�tDr!-��>��Qg0���LI��Tիx��]�!�a�L�1���c�j��-�[f����6V�6�=���Y�m�'{��'+p���+n/��&_�eor8%H;u��u�bz�w�u1�~yXA-���.4�� �B��a��s7�Aݿf,�6��z�X�FX˥��-����{�w���z�h��=«0�B��b� ?�Zd�>ܬ�[����N�ů1��Z�t��Ļ(�X�v�(���r~?
�G**���R*��^n��	|T��>}7ҕz��+8�1I�_�J k�ڶ�k�2��)�+*\\?R睪h�<s�nǵ��NY�WNUi��N�����Y��׽�V� �;�A/&3/�C��j쥑�������u��-�k���E�?���]`fn��,�h����L����%w��3���T��z�b�_��O։߾�lZ)@���T�j�ʝ�#��6���~&a�*TG����#?�=�^�y�pe�y~�ތ�lŜw��A���8gܸJR�����g����ōp���~�W�&���b�ͰJ���ΨE��/(���/U����!��2S_�>�v٭�W��K�����H���h���
,�x��!~�/�2�����E���o8.�Uq�of�^<���!���`c��yu����W�2�JJ�����G}QALhQ�{�(R�f̠d�SWW��cy�j��i�b-���������ܟ8I�ԡ�J�Owb�_4SFo*L�|���0S�\غ>7::bW�BЖ:C��1�p�Z�������!�����H(�K�����@�˪dJ���л�Q�f��j���E&����:�.q���3�;@��SQ�(�e r��[`�.R��_	^�$��
�@pNY��&��%�T�1�M�SC3*b�������F���kM�����yL�+>6�� ?L+�AS$���WﭿE�|�;��<Cj'u��TE���_���;�!�}q#
vG�a���w�����E��u��,f~��:S�?�����O��S�\c�!�i嚵n�����B6Y�jx� �p��������#n'�/dLA��T
�����R�rl��GD�(n9$id�c�s;e�~���������oGĩ�F:,߻��oQW:~p�Mb��)˖��y���Tq�(������<S>�i�(��x�(�:���O��b��-�+94�k�NX��~��Q<$�K�˹5<�_�y{��Z�+s�~1)���]u������!<��$<��)#$,�K��VW���C"n��p ���Y^�x��;���J%�U�U��D���ړ��q��D[�xq�Bk;G
���TI���x��`� X�3�)L�4g��XX���0�?62�?S�S���Q-��A�	q'���Ft�4ZoO7rRB��W:��"�)��5��-�؄��]ͬ�����Of��p#ht���;~�b��g�u�*������<���s���=�,e6�a�ٰs���dR�B�:��p7�e�V����)_��Z?��o��+�+�/��XZ~37�v~����c�����=�^ h�n��5O�$^�O��і�����_RߊJ�Y��p����Б�~���u�"}kI$o�5K���Rhi���z��~p6����L����?J�Iy8-H�V�[H�m˦'�.t�}�<�=�豓~-�$�*�F���o��i;e݃'.h;���_Zm+�m%��`^" ��U�IR6��3��n��@)(^:�z�ͭ�.�"3��c4!'�Ü�V9j"