��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�|�� �Ǻ�����K���Z�H�u�Z��SS� d��yL�(�k�&�$�7�{�/j׻8�K�B���%�C3�rI9��:�H�!��k��*�����6"kZ�"�(pK>�(� �PUr�u�Nz֬hg���Y� ��?j�X�8��}z�a��6m*w��'�`��d������N E.N*n������g�sK�.�*.�A���ʐ'@��8w65U�~��!8\ "�Yt�(�֤j��5 �/����8G�C��MhW�x�5�+���bp�
+�'�t�㩭�)��)%�o�k@�湇��&a��W�I�3n�����z�TcT�I�}dE>(R!/i^3����՞�hC�BCfܑ����n��U� �Wp�)b��@�OƩ8��s�r�2����\Y��bfSYjj}J-lW�t�Wf�{�.&����2֔S��mYz��c {�z6�L��|K�]��-�yI���=��q3aiE�n��yԒ�ծ�=�X%��fc1���G9gF���t���r�`�vƞ!
y͖��BX6�عPA������8v��2l��ʦ�~��z������$��0�&��i�+� י�?2���z�u�z���@�;�f��E�����Z�����M�DdW��~����V���Ρ�YG��D32�Ϗ�K��Ҳh���mC�Ů<�ս�����ە�H��=��߉5U�O��m�=�Ak@[�(�9w�.�Z�Zcj���s�l�(��-#̽�U,�C��Ƌ�|8���^1���l]��Z���%�8E̊��[;�%��Z]PE):��sɖB��cʈN�{s��I��G�x���N%�3r���,*f�3��٧	�y��&��$�	^��h_��s9q�=��������[_Œ`rR�>@h���r�T��G'
\>8BUq$"-|���-�_��!W�0ָΘJ��v�m2"Zv�:���3R�.���lR[����eZ�A�9��8�t5!'��1c��ahG�l���}߶�eA)�rZH�,�J��͟�#o�+-}�RN�HH�'֙���,y����-�~�N
��@�G���3a9��k�\R҆GS����%z�xC2"	�&�ykȓv>�R[2�K昁 �Zґ�����}�}�/��4�U�C�D���g&A����.��p�5��N��;��Z��"�3L�!���Z�"5	�����"���{�fn='��<7�j̜	�g�"���%��:(l��u�g-j/F�٘�~�kW���{��
zf��ҭ�n��iޘ��v�=Xl���xvw�D�T*��b������m�r'W�L*�7���M���Af�)���S�i4����D�tɛ�/>�1�׆�Px��h�������AQ�	.7aS�q����q���zKe�l]�T%Q��oG��|69&�+��H��L�FRV�"��
�IPkZ�Sz�M4)��f#�a�h>��x0S9�Vuk��2�S^	C����M�3�Ky����/�ۯ�K$q``a������a9`m��uBk%����#L�1�q����R
�6u��	�l�� ��Õ���>��~%�d�q���ou���7�Y�
�Q@D�O��?�Q9�u
OvͺZ����H�D&�t��lA�BJO~���i�]X�?>�Ѿkr���F��ӒLwKr�I���G[�2���W��-Ud?0h�� �����c��\8�sٿ���l��$>�<�~��iYj�AGL
P�C(����7���.�k�ĕ_����l��A&@�t�&���SxI*N�ng3_��� �۴t��O����P�'_ۢ����^�s�#$��S�dDZ�C2v�g�znK��1yw�����/��|����6��>�zp�j�K��CO.��?45��E�><*D�4	B��<����ld����Tc.�~|p��m��aG�Rus��qD���5T5�I�ϋ/�W��̨I����>�A��t�E�~�:1A���� �טN�k-���n6�9j:m��2Tx9p��@�Wi�J�J�sW�Su4�lɨ�8���Bo�|�S��x�
v�yV`tN�_n�hS i�}��	�i#�f�Ҋ1��1���m��^��/K-����_"*������1C��{-X}����o��^1f��L�i�1���o�b�#`��2n��ʨ��gZ6o�I<���ʷf��\���ZP?P�J��� ����Du1��{^gk�-���v;7,'���w��q!ߜ��\x.Z��+#��B��B,&��HJB����x�	��u}��)7�Wo uт�O`�R��A8p��RƉHc��oI^�ZiU�E3ZJ��R���в�-_���}�}@�4�|[�,��'�����:$eH��tLr�� �#t�
����:,�	��>^���fCXx$�������Н��8�\|rg ��Q�Q��O���Ϟ��}2S�[/��;�m�Y������8ˍ�A�|��=? ��"�&���i�#���-��� ���f��hm���F$���b�/�tQ���T��'���.ߡ��X��;���J0f�ѰN�68%�'T#ϳ���)p�,5h��ޒ5] ��7Ry첱@�]MH(-b�rA2�uHUX�3���9��H��,"�sI�gK,���lH�鑵X���˛��u������(�YZ��w����g��"��|/.�'|j��]��0b��k�L�+)F_V���C�\������,� ���p�V��9���~#��)u8��f:����d�g�#L����U�#�8�ץ��Ǎ�22������1�a��)�B����G�5φ�;9���'��M>!.eI,�Mv����L������˼��쟉��e�ߠEn�&+K.:���/����q֛ȼ�8!m�	�\���a�����=�-��`4`Ѽ�P,���@6��v��uj]-ٌ���S�u��P��JVO.�s`������O@�~��TZ�;�����f?Ow��J��0=��R"_���5��y0���%ɿ�^��)c�:��A���-L�pA%Ȥ�~3]�(g���2����U�"=��\�r��K�D�{�u�؟˵`ܡz�-�����b���!j��#����Fh������q���"b혽�4�az�:'G0�߄!��T����>�~}�kaVLQ�I97������	��%�іo�l�^Rh��I��4�#�C+ߠ�����S��J�٩̓}�k�O��w�����9��֢L�Ğ?��*
Ƃ��.H�(�}h�`⻽]�<�!|���?�@���z��LL�R�r��Z����֒��P�&�kF�d��D�Aj`oo�R{�������K�"���(�m���G����f�?��i�3�Q���1�!��r�Y�@!{�����bc�*�R��Z����QB%�����K�O_!A2�V�J��g������v�����U(d�ab�ڽ�"̹9-	������E?Y&9LK	?�z|���[A-=�Mi#���"���p�a
�IJ�4�m��C��W�KE�2~�x�:��r繱d��?f��T���訯���)Z�>�}P�f}T(������"��O��q���R�7��P;~��e=J��>�B��'o^��ztn@E���xM'zZZ[P����
j�7h�a�2\�SU"�И]Y �Ud�>-�ق0>k{>�J���J®z*��v'�<��D,�Ͱ5��-����]��nA�HbB� L�h֔��;�K������f�]m��ֈ�hKs
�͗ud�>*�
/�~�2{���d�M�^"A��\��3N��Cw����}=0_�p��%��<֒[BYqb�>��̍��1�Q�z��l7����̴�Î@�HCd;�f��]�ؽU��+��w��@�;0a��A�?�\���f�1���U�����v�������(��@d��=�Z�:D����@he{�F��ށb,�pn��7Mv���։�A��O�jVm�h��X��]��IJ�Q�̺l�Ot�X�~��J�O����R���2
�L`�������)C3�)�� E�)v�q�y�N�f���s b�]�8��K��jX�*UJd����}���O`O@�79�r�R��;�I�J���Hi��H��(�	�;L�H��,��f����*����S}�4x�vr���	��MD�{�)%�kO�|��/��=L$��I�B��,xW�H���my��+����0֡�z�X���1%b3AZxG�Rz�D��bl�Y�w��2�.�It�$G���� ���fb�N�(���t �'��;��s�����ׁ��
^Jg��Qu6�	4&���W�i`6A���W��z]���E���3%WDp�`m",+��~aw����xo`o�c��a�`���C`��Y�����Au6Ns�h܎���z��S�(>q����%(+���4}f$�Nq<U�#
L��:�C%>��sZ[�
HTt��j�Wؿ�.�U2�_�K��<Ml���m̸Ei�ŷŲ�ʎb�a��ťz��ڸ
�8e8d�6�0T�Ϳ^Tu���>���F�TFc/Pqv�Beً����/l�zs�,��K4��I׍ �g|��#��+�9�z�G��\痝W����Wi���&yy!C�(c7vr��-?��~@Sc�H�Hv�++kO��J~D��<~��:�\^��/:� I�@,�;H|MAGL��S�L�̊MO�+D�����Ob���K$�i�s�2��R�$A2���a�s��D��H�ff�q��eb��đ�A�|]'�<���7��y�<��e��-�w蚟��������=��zG#͏`/Z�M����X�k+s�&>�ES3^@CO�h� �ƻ����������+��x��Hh����Ia���!��ڹ������1W�ts����+[����1��T�g �=-O���d��9
?��6Ev|�w�itPR�� [�l��un�_��S�m��9[�Ϫ�^WC�Oe����	pgE~���y(Aw�'�z6ot��]k16D��h����9yX�Bѳ:\Z���!{b�(T�]�;ǥr.-V�yjM�@>�c�ю�@Ey�]KSFx��,$�	_�����Z�=n�O\�"W�W���{�`e���[b������uBjw�_��aeX/���z���N^�c����%S�,��<��X]�esn#N�U�����#F!�c!�P�ˎ����s��@�掛�u����á��Jo1��+\&1�,��
�3z�����j��;.��p��[�ב�~L؀��D.bz�T���vm�q��R�e���3?9��/�e�����t�'�fH׋��%�Q�q>�/��G�����������-���ǎG q>̆9�T3o��12��N}3����~�YJ#:�K�!�"�o���ud�~F��P�����dS�<�}��}-�rso� {���0�߇�����VY{��j��홨'��tK�o��}��p����]���bj���MA���4.7o�\6غn�+��i$��3�}�4�]	�EX�\?Κ�ۍ�kxd���$<���H7&AS8�Vf�/7��q��	T��2TE��n!:��o��G��i���y[��ũ�cu�/���������U5̘qxL!�/V�h�(h�D�D|��G�wߎ��<,�c5��s�В�Q���Ӿߤ��,N���(�����B�9�I�La,ڠ��2 `�X׊0('^���f�� 'Q�Hl�N��дÓ���u5x@��7'�IN��c��O�|b�Q��~q˥�����	��+�w ��}���� f����5B��:���c�_��n->A��۵�O���H
�mJ$!5�w�%BѶ��1�7�s�o��Mgr�i&C:��\l��9a4�Iс��{
�/�����:K�����Ĳ+���_�j��Tk�� �VF�Q}�g��\�tN��c�����҃�7@G��ڹÏڍ�o����t"P���^w¼�O=���w�����|?�~ .��"G���X�5����	_gy
�ׯ�w��q�w��hO��CC�퉋�bF�6�����n���~�F���+?4�,U|ߙ�'[�͹�Cggw�'�FN��d�b��w~q�ǸUn�}�U�e_%�-�� (|^.fi�_;d����'NN��xI{�����U'p���_r��L�,�3Y��\�M��ve�^�����`EaE�rD RIC���J�D���x��g���XT��U2��N큞�b�fY�������.6Sx��ҷ�T� C�Y&�ff	_)ٴV�y�?^}�Ąͤ�c�ÿA8����W��<��ڎ���.�"��)e�����ӭ����8���F6��JlN���w�9lB��t/o��>a�*`#�l�O�G��QUYi%ś�qe�`0Ӟm�u>fl�O7� �h�ѷ�@�!+[�H��)��.�3b�RY+޳�����|��ݿ����E�v	��sK����]l�?�ZR�Z�y'*��
O����pJ���Q���~��;�א�q�����ʛ�N���h�#h2q+	�4b��d��*�FYr���&}�Ѯ7DK�̇�v|�C�&��e��r�� ��[��e����s[�AE����s�?zP�?�֚�!(��KZ%R���;���w��_�/�`7�*҂�j<��k�C���k�CK�8�֧� ���/W.����x�cb����j0&�DC`N�wjL�q(eČ �cyK������@�Nْ3�@��6����c�m^�!*P�ʁ��(��HJ�nϣ����@�v_�C����jƄᇊ�B��]y@U`g��8�5��Q��B�,�rg{H�[�z�r>尉d�`,ԥo@��ei[����2��D�4�@mT�1�I�	/D<O�9��.���k�%�*bЙ?R%GO���H����0������V�V��3w�ս?������*�{zg��>��=�hO��	�Ͽ�Ч.n8�yOҬ�D��J��Jt]@^��-�P����Jg�fZ� U=82�K��RmgG�h7ңa��b9��,ЉW�E���3zGY~���lR7�[�Ӱ!�
+mTO�.lPgR�J��m#��ˆ!�r�p���z=]���K]+V!���L�7�ZuN���޼�0��V�9���9
z�NF8}�Z<�8E���s���Q�^�x��g��+W�jku_�̼p���O�Ac�x�
�ɂq��Qyub6"ˏW~/��@�Sg�g~������b����f�?�7襷j>��+2il6�U����!z�KwOW���K�*ӭ�N��)���<�ÃHe�:�n� ���rBw|''��J	�A���M���A��������|v({_���m�Ҧ����E���*�}�7�p�c4	JH:]:
yx{2��LF6O��V"%�j����@Zw4�����F�����(�Wڶ�zx��Ow=W+1z���u�W5�Gv��Α�#��VtR\c��Hg�(jq��Jl��7�nZ��5�a;�Y��j~���e��*���^G.�� l���1=Kn_����̏p�gW�-��ȯ�u����R�:֙$�s۾���np'������MwQ\���`-����׈1K�%C��n{�B|��R�M/�*�,���\oL(�T~�N
�������`��.��n����y��n�R���p�+ͧ��"�������+9�ً �4$��<t*��z���P�-	S���&��b���̛B�_s���u��fp�c)��C�aC�f�W�gD\,:A �ed�~w��L���{@x#��ȇ�­D5�lmN!��Ԗ�h�P|S���!'j�����IB�ϻ$C��DL9�S�V��W�����"9���E\̸4}�q���s��Eq�r�ʯC�/Q!�D��i��������0��^a�����PG+
����9Ƃ`x��;?�fc\���oB�5/T�Rp��)��Z&ϸ��:�c�/ߨLy�6l+���m��2]ZC5_'� �ß���R��� �j!Hh��]j��=!ρ����o�M���b�+�%5�)�'�Ԝ%���6>_Uo7ǧ���}�����3\��]gj5�t����c�@~�	-j�y��4�v?f�C�D�'!K�:���=�ф�<�c*�?�\�@���F�|[�d(vN���CaW�^��Y>+��1m�] #��r��3�zc����y� af3�=1�����{��o%Q#�����_N��$��ˆ��"2��J�pL��L@E��ƭ����O��LBg�����?
���������ɻ���VEx�-~W
SE�Њ1�Exl�?�j�P?�8�Q���zޓ;`�]�jͼC>&����5@��nRC��U��e��k��CpY*�
c��n�7��iЂqvt*42��i3���g{T��å)��E�%p_�H��0�����f��b�=��Q�qJy`�V|��W��B�_A�}a�(?c@b9��Q�u��t2��ޤ�{@��z<����pM�ߨit���=O[�,$��~�������V]���t|�:y�->�� �	mAztl¥B�����ؐ�����w�H���|���;�(誓v�J�cW���w��
��En��po��'c�բ;���L�(F��К*�𛎞/Р��/NqX@�Cmˎ=��6�_1s�b�V*���L��d�~72=��]��lbz��ۄ'1�6m;>��r��hj���PV�%�r���pO�J �W�U9��w���􁷄�X V�'H��u9��p�i�m���@�Y���ra�[bq���]F7��n���<P����B��������-d�T�;�e�a^�SW�Hl~��h�,`�ߞnQ���x�)�k{3��v�k�"�ɶX�o20^��G�8߃�q,G�s��6��;V�(F"$%zס"�~�t�|�r��Po�a�ü{(<��ɓ��9�������,�Re��~FOad�4_�3{�+� j�VG,
Y�e,\de�Rl�G����K�<�8�ϰ����!����ۗ��d�.s�6L����A=�t6�Qh����6���t3�WҲ����uo	&��Y8}�'Jr��wc�x�Jݨ91̣9� �H��G��@j��"][�ʡ�AEQc��~+lo6�	��9��"l
%�P�R�sJyit�z��P�rv+:�?�K��������KK����95�9N�q\�$=�-(���+  �=^*�7DEm��5�^�v'����W7غ>�5���Y��/��I��i@Zbi���B��l鏩D]����q4��.��`I���)�2�j��� ��W�9E�S,[�V�W�n�	iŌ��6~hD���D�Jt��tyUVQ��@�M��#���v�Fd��+�����
��#%��	�凲L�[V������l��Z]N��s�L�g�TK?Ϟߵ�,�M���IH1*J�Hi�Q�_��Ytɻ��
d�fo�]hn$��KʖN#�y��y��3(��fb�W��{��ov��o���+�݅�Mrr�x���D�����	E����9�3z@_swW�S8
�����+�=l㲇n��:8�l�|F�ڪ����]*a_���!��ǟ8��_���BOC�ѐ���H�E��X, ɭ�&,�]�P�M��sw����@�>���<��g����t����u�p���^:�[6.� SB��c��I�RC}ukEތ��:y�'�9sh�ն5#�F���I�6����0A.lL����>؁6��w$5��H��q�}����G���J�¿�����(n��~m$�0��LL�{�`[��[�$w��
���.�Zn�hB�#� +��"�>�^gK�X=:�gW�0�����J�	�<������!�A�@�k*U�\�����c���|K�$-ߝ>t��=t�ճ0n0	��=�O����\�K��Q����E�V���d~�&;�xI��a���mr�8 ��^P�2H%$x�[�+�L4�>ƍ�d���ځ�3]1,�n�԰��	 2���@-��͟�=}{hK�*����� Υ߃l��ɝ�A�5>;%���B��I�x��e3ȟ6�}��A�`��㳠$ǥ�%�t߸�u�x��|HqL�Pcͩ:D��7kr>�(�n�bS
m
��?Po���I�+��`�{�3�����p<����3L����p���d��R_��H�*X��j��r��Z�6֬�(L��S-K[���#�<kKW8Lb�.+�i�kO����$^�xx�}������5j���/eJ�XE�8(%޾Ir��Hx���4~=�⩥F��e�go�}��8�T�b�ƆPְ����6���XGd�Yj�A��jT���9Pl�bsi~��$(��!��*�A?��DP�q�Rn ��W.�G�����h	\���$ʅ�?�e�'p	p���t����9j�m�d&�|Tu�oY�s%(���OO����W����t��m��A�d�ҡ�]i�x�-.<�����&�~g��,DW���z�H��y@̀Qޱ�=U��
�;����&����+Y$wF����|�g0��
���¿��A���m��Te��!M���Y.A�4r��O���3Y�<?/�hG�ͶG���2�ϩų&�u2�[��#1��<c�*��t�n=3�0�ZI��$a-����J���L��c2Uj#B�A�� &�G.;7�i_dR��"��U0�/؝���Ҡ���	�ͫj� YD���;�G�P�xR����,��4�%��0�C�HBO��[[��,8�,��)n��Ti�=/�o�����]8~� +>�վz;f�vg�X|�0,RV����_�yg��r��Z�4@�I����?3pG؍�;�����Y�Ų�#��
��:� s�W���H�V|��[�=��u��J��+�e"R����R��@��*1t{�d4���?�-�}����8*�4vq�gT=�
L;��>�:�Ց��N��o4���q����[w	�
����w�[�[L!��,�IrpD| l�6��i�^��c	�Q�X�V� ^��ƃ��*�I�O|����=I>�|���[?ˑ;@�zKq��(ϧts 0Fɠ��%2��/�R��������~�荷��o�{i��̆�֩{Z��H�ӌ�O�	���Cu���aL7/��@��m�&F\��'n]�|�5�7̽��m�Ֆ���X^IQ~���$&�[~J�)~�N�g,$���ȳ�� vz�U+��"�
.Յ5ߓ �d ���򲟽D�{���b$�u�N:���=�W[߽~R��)�� 78�W��o�FhG���@X��=�g͌�%��޲��I*g_D�E�Ҏ� åɼ^k�.�<C��D}��8��Ȏ�ws��N��!Y�-̛���*�����Y2�5��t�c`�2�I.��=�*�~�/�\Byw��i���N���$a��r�{�=��!FO��UvIz�-� �}��t����o��m�-B����T���B[Z�U��}���s<j��9b��_Q-~�f2$�� U�4��َ>~�r��� � �=�~��}�p���`5��OaO��/W׼b��cѶjL���� Z^�@ݳ����WL@_�z�-6?(ȧi�X���o��Y��/��9��y���0V�7�$��:���`��G�˷`��&��23��j��������1�Ʀ�p��\;�^�ԸQ' W�N���V�q�KƮ@�"!�oś��T�����	 
����h�:����,-�RT�OlFO����`��Z��dO�	/�ǧ��"	��,�)kN`�jŻ�a��;N��D����!�ïj���R�n�����\��yY�P����סMǢ�B��k�<|9Y�%m��,[ ��[�HH��JA*��5^T�`HQU�&~&������r�4s1����q/����g{N��<�v$m�5��Dঋ�vp����ߐf�ѵ�+s_��+�C�xCݦ��N��	�֗�j%rA��}dLL��v�lo���hI���p:Q(|�&����+Y��q��.Ǝ.�w�"�WQ���_��Nc�T��W�b�I�r��ڳ7d�Zo�zz�\p�mHܣ�t�
����XE��M�2W���q4<�<Ew3�5���s0��1�|�I�<�F���.���}�/X�?WݸA�%����B0���;4��Q�=]՞B���5{q�������;d���ӑ���̭��T�E��e��=8�k��Yg�.��L�%+=��`%O��3۵<��������\���9����x_��g�"g����}������=���h�"���LDD_��i5ì6 ���1�Q]5�(*hʠ&�W�kڔ���5�q�T �uV�1�yI�voCX�ϱ���-�,��5�&�,$z��w��G�4q�D챬9���]�����h@?��N�᫶�c�0�@��P�\ǇK�`b]@p=@������r��;�wO�/԰g,�� �Ml��נ��ݐ��1G��%<�*VV9җ~����B�VW��C�D)���X����+.����u�w��	��P�=����xd�C\G��S����9���!�DO'91�w �~<�!�e�X+�h�Y�K�a�[����D�lcɀ�	F���Ǭ̡�m!�C���'�mD�db�h�MVǨL4��6��ㆈ�V���[h�{�ܨ�>	���!�X
7�߸�E�lG!����GWG�]*wL�Sfq�K��^Q��{�n̮v$ �h�k�Y<�uj������^{����?
�9��QAW��l֟d8�i����U? �5�
Rqп�*a.��]��XC+����!�=ױ�T4$�P��i�Q0$9�䤎堠E��B�����G����$�R�r��4���j�Fcp��AU a���jV���_,NTHN�QB�O<wl���F�S$I��δx�G�Y�{LIdڅYg�������S����,��R�+�.[�M)��3�waϪ"�+ ��ewS�NC:�}�e���S�or|�=���U�@�c��ڹh�Yǵ'�{1���Y�Nlx��RLU��BlJ��>��lta����Ā�c�yW���`{��9�oͿ &JSZ��l^dy7�U����*%�Hι;"\�^+�� �{8����e�|��~�?4�������`ݗ��/l��ܝ9I�c��b��w�����үP�A,�#�E�}��D����8��a}u]�	W�r�Nౠ�ލeT�$���<���}��� �8%���ݘ-ڮzh����huF�p+N��~�̮$��I���<�X%b����R�.�3G��tH���S&�=Rؘ<�h�=׿�"���s��U���eyvU}E�84��(���$��el�G�BЕb�TN�u��y�t�"ݞ��h����������:�O�O��sԹk��-��r����`�S�n4�#_
�E��1���bW#��B�=yϊ
��"n�o��t��xC���nM�`�}�gw�:���<���P�.D6&����"���F�>��^�YpX��^�]��A}
����_���f&v�7��8�&���@5V�?:mpF�zd1�,v)�_aϜY��L�����q�sޮYJ��q�XX]�������Up�HT-�ҌFX�Ǹ��	UWH�9g�x�mc���Td�J_�Q��J%������)��iժ_�
1O��.�Q�����gL�;�����=�KZ]��<q��(�.��ƶ��ԍU�Wp��EYx�ZG4��rP�4�?f
L�P�l� o�jU�m�h�oLd�n�4S�B� 7ɹ���v��ߟ��Sv~��U�9��ʇ�G{9�:Z�5y�C%�vG�x�!�/?.����_i9M�y���/���w��m��q�D�x�ͯ�� ^�g�独��B����o�Y�
�X�6�>jJo�1#�!��ڻ7^�<�V�wx�j#F���s�n����0AG�?�	v{^e"���-JZC"|R7�Y-r#�Dxc+�{�m4�ؙȦ�ˬ&T�W�}��ip�g\IŬb�~�+�A	z#m��[hiӊ��e� �a��D�y�ԛ	�E�!�Z��[5�\��� �3��k0 �D�;���S����vdg	�������b�l��]��Z�3���)&��I�Ƨ6�Z�7@�0W�X�Q�o�īڇ��s]�����b�4����� �X�6v�FH/R)��xs���
ԑ�xN<u@��n�;��&�;��]gCQ?��������;(H*�ȅ��Pw�N��� ��Ɨ$������#�~�������M�������I�5�$�2� �x+�6MAF�V Y�~JB@D"��M��xTi�3������f�����rTA+(��`��cѱ���A"�޸Uɕ�~�<����R �&[di:�������N^ �}�M��	��1B�8$�@��/��T/��������0�9��� ��������Z-� ����<Ȋ�p�t�>!å�5�e�e����Q���T�U7(.%�bJzrQD��L�>Q��2��~nuYLa2�t�x㐳��t���0]_��J?j�&��(L$I(G��R�U��My�
���B�Z,x�ڮC�8'������2܆$6|�sN�
f�R�p�M�w)q��?�㱄����^�D��\��-0��Pd���)�;,r�E��;r���3��~UNu(^|B���zy)�m%'{�s�)�<��1�����B�2��xYz����zα�J�]-�8�����܌� ��2���J�^��!lN*��Հ���$���#���@�ZĮ�#
+x�XoF
0C�� �a�&�iv��9�Q�%�c3��M��pW[�.W����CퟕOOzԚ8̎�=200�	��S�>qx�����@F]���Q,�'�Җ�gR��4h~��*�4�c^9�M�P�)����X�-K"aF���|R��A�3,o��R��n��<Ly��'M�Z�G5^�P�!SN (/1����e�N�cE"4���VQ��|�^%���x8QU�sEV�+,[���N���<O�Iw�Qw%�az&a�5}��ˡ݌%?8V�w7�^`������
Ѣ�蝟�C����o_,��eX���z��-�Q��+3D�G�7U�&i���g�z��ox��U�e��M˘�Dq��+��b�u)�O��Q#v�Y�>��Um{O��Y�lD�	409�[���ޓ7�ˉG~�`n�wIK[1���yo�j\�4>Y�@�ɿF�P��߮&͑m2�eĭi��?�5LG����"�pH�R�Y��^����+��Q���M-%L��Cu�[e����8S"�W�/���,MY��G���2���n�bv������8�=�N!��c�U'�E��c��T��}^�f����
��d�B���т�^J�~�Mz���E�10My>�q)��N��NR��1=�\��S�X��sur��YV#[�T98 �,��YB�R4�p4ip� ��7|�D�-3�L���<�J�>�L�sVe�aa��ϫl�9b�AXL�OC'��:@+��aUμ��T���)W������K߿����Yv�`�����`�����q�`��r�8s�Cd�s�c�Q�_5����h�X�r�e	��e����<�;P"��oI]�S�S��������Ἲ#d#E�f3�[�b���l1[�^��6����y�?�>(*��h�����"8r������*d����rƾ}1mw� ��@`C%�>�!��u"f�F.7��&�Γ�3U�<E�a�؁#�?��p���ꉂFPL�[�2�n)1:�*�g�ٳ	��M6��������m�jw�P�����ֶ��8[��ɬ��aÚ�?��^Y3^Ru�W(N1���Ȯ��S�`�n{�o1W�=`K�h3���뤦J��H�'����Ӎw�3�UwI�̩$��A�����%tֿR�f�h�I^R5���`�����B� ��_�X�E �-���N1�R�����4`nU$��mp݂�F�(���7g�Qik��7���B�
���}0� \m��^���!ٛ,"tj��o���J�� I�8��bl��x�Ö]I��(��{`[APf����\'��� t
����cY�=�Kz�<�f�~�������J~�[8�И��3M����u[�g�P	A��T��,q_�UR��1נY���;�3�p�X���8�dk8D�d�#3�x�������h���CA�˹�(!<��ĹbM�yS4@w�-�*Z����PהL���C�k^eD)��hNh�,����~Lȡ�M���U ��
M������yu͢�X[�^�W���(6[PϚ?�Z�˫3?�b>s��"��L {Ye�=~��'�>�-+��ɭC�R�>?����Ȃ�.$r<F;��j�����fk�7�2���c�y��@��x������w?j�֢8tNK�J�s�Na��i����E?����a;7�t��i���>ql����Pg?J�
��ZYIT��Ք����� yX.�������ų�����@dD�F[��˲ʔ�!R�4a�'�#��-,hR��f@%�$α�7.�$_�N/yz�}f��
��?̣},��@�ø��MglMw�HYP�ۀ�V�4�x�O��zB��}��α�frQ�l@�R=��iWH4]��A��F�6�m�|�xrLv�B�;k����e��� b��Tw�(r� �	ǺZ� ���Ħ`7G�٥�>�M¨9�'ٽ�2FtsT	���p"a���S��� �ՃV)�n�m�`��
ms�:%aI�rBqTAc��w��=\��^�S7�dz���j��>_�WY �f㐖�:J����,(q*%}->ot��Q%<[�Ϯ �$"�c����x�m�F�A�H���Ӊ���	l���©����F�oy�]��9�t>�Dh�$ģE~�	3~�2�JE0�!�ZSq�nɏ�*�!�,}Ϥ�VS^Vz���|a���ᮣ�����|䋑�5'�+��Ő� ��伹�G�7l�Q��*e�v(��҃���aw����d"�S>�&�<�E . ��徲�9@s��w#����z�9�� �5*�i�NYgG��RM�7��KOl%� �J�Qɒ�D�[���n}!ĆZ5�:���Z3�ٲ߱=�R?,~��0M��2�^@��� ��?2�gj,��h��1��tZ�)���y��0����ۜV"��Ƥ��sv�V�Y�ӧѸ���2����H�"�`�+ٯ����o��vd*�%�����e�¸E���?@Z��]�V�G̓��8�L�׳�ܸp�� ��+��V�	�W�vj�&9e�����}�8�R��`_�Z�2�y�J��Q�`��q��mg(Mj����Ϲ�����/J�¨��ه�GD�K9��:?2� �oʒ�ow�$�����m-�M��?��+ZPM�f\U����^�9�/;�OB�Q�\�����p�텏ڷ�Z��W���V֚``�!-��mQ�Չ~�_�9j}c���-��W��l�K.#�t�s�L0wb��|����ޓ��w|�I����Q�f	��{��U-��Y+��+�j�,��3M��U���oz����wa���R%�K�x�<�����/��c-��Fߩ�8+0k�v�hReI����jf>��.ԍ*�}��-m� ��Y~z�#bX7y�����cV)]��.�T*-�w�h���ml3$�0����%�p����>���x����|}�߈rd�'�&�	W��֘b��G��S�B
�U���@fX䆘���ٿ��*B��7�;޽q�r-+��L^{!����-�g1�J�8iZ�7;AG��`�����
�C˗�,8ԛ��Щ�$""��Ɍq�յ��^��2���� Rr�IYJ������jD�0�r�l�,�,5N��)3<M	n��a����=N��V��+��u�%�ޜ$�~d�Cf#��������:l�B�MϷ�2U}�9G��QN�6�������65ч�N�tĲ�pXdf��q=  &[W�`��iȅ�ې��=L3��^�j$�EQ4E��J+�Wߖ�l��c��C���ƒ���o,1~�F]�L�t�A*VY�L劐�h]jF���S�;��{t��Ԁ�����F�B��lgMq.��������y�Xˬ�ӮnϪ����J�>�mqdH�L?�1В�앶ok>B�
)J�A��V:Z���:`���T^��a��z�|�[�m�*L=M:dI��ZRL@�I|���͐GχP�_��3Ft5���u�4΢�m{�)�:�ІM�4;�ء^b�3·_4��������(�,P҆Ǣb�y'A��^�w��m\cr�v�p��>S�0W���4O�ɨ�����g��8>{��@N��'@}x�r���nn>ms�^��{�j�]�v�x�����������
G����/�Y���g�IAsx�ݏ�W#NRiV���`�&��d�3XɪB @�.]#�~k����/��>vF�`����Y��JQ��Q&Z����rRǫy�p��p_�'?���Y�}�x���W�{� �p���_|X���GC�Z�/��b+��G��7�o�?����6*|��iѳ��(����JY�+q����Ez�
�J�0���?�T��G��?���\1�~�IL�s��[�ѭ��$O[����O��{�
J<�yqR�>TZ�@�.e)T���0r='X!8ę��(���I�L�1+���C%��'�Z��9<y&w����e��WEPUf��g_��{�`�Y8ڎ������C*\�;<wk@�Ƥ�4`O���S��^�{
��o76|�q�`ܧ����%���)@]�Q�Uب�o)>w�C��Jb9r��|]����忽A�F8#)���§`����E��C��ѯ&s	*���r$�2q'�&bܭ*��'z(t$A|Z�R�a�x7�`�_-�xgD*w�+�/p�>�m�q:M;mR�c��`��E�'�#�e:g3�\��}�ԝu��p����A�@5��m�(��P%NE��s�"-4e�rP��9�S�S�*�(�e�"r��}��Nv�ޚ�����?|�����|J�`u�U����D[��~�Լ������]Jy�8�MKU�v]Q��+'���o-?�s�?����1�dP�oo��]�L�YV'^��W�M{��'y/����H�k���/���uS��)������z��?����Mg^Z�8��b�@𥳐�c����1D��%o��7�����I��~D�a06Q�x}F�1!]�ԿdB�qC�Ph����)�"�3�2�����K�1&�
 ���3n�������LS�NB���Ꞝ�}�m�5d��!�UC��6৶�(_��Q`I�|7�R=����~�>B��U�ֹoI�iӷ��G Ö
�����W�KCC
��z\�ɧ\�e���~���n����K&���[�0B<ɛ���Ǣ������{��\�!��=ӕ�T4�:޸�0�ϋ\T=�}u���<;����ikn����#�s���">��}��U:A�Fp�a�[sh�.<���&<v���E�� �S�bh�QԱ-\��Ǳޢn㕥?v�H��N�� �����C�Of���ᘊ�<�(���������[�x��/��eJ����b��s����a�~��A�PP�)cY5�(u��;�+ooG� |���6#w[G���C�B\�I4$hYϪ��T��e²V��K�]���j�ޔ������� ��"��ܲD#ӑF��$Sۣ�q�~����O`��lB�u��HܠI��6%O��N�e#���J�N+Y�kt���G��Y\1#�ؘ�����iqo/В���LW�I�4�#G��o�T�����0ͳ���*#���3���Ԁ�h�a޹�����1oiS��ln�;� ���0�!\I�ё����ک��P�!u���P�l�ˊg�]��co�3韷?�k�~��5G�]���Jy�
��Qes�����.�H��F�{�?g�˳�V	W��ֿY/B�� �q'b��r��,~�I�'G�G\��T���,eF��'��z�9;�)c�g~h����kR�/8��N=k�j`R�5�V���G���?~8u*s��_�3�21>zT}ŐtF
WF}�{���1
��F�%!�Nq`F�@�_�E�z��Mܩ���+ċ����$�)��Y�^��>� ���1��Ur���9~��#�I�����sn9�|��~��#y��i�~[v�?�bcg��Sn
�?�	@�>��g40���ltr9��۳������^�ɼxG1�uhCc��恷piQ���Ķ�^�k��4R��ˑ$8(n(gͳ]Yj��+ ⯶�$A9�g� ћ�B�.x4���dR��kiG`��ۖ?YGcj��`bf���O/�xX�B��4��p$�9�E�8����$�W`R߅�s7�h�uͼ�ׇ'(�$�(��H��~ѐA#43���� Ry�=�w:��<}%���aC�iv�Ë)iA�Y�z�
-oE/�������8��;�:�s$����=P^,5%�� �K��
G��;���tO]��?�Ԕ׾0�0@��m58 �.�pE/U5�p��g��e<h8�C��4W��J�՜�Լ��nԷ������U�/)&��xꔭv�|���?�a��
�-�b$r>)�Cs)ծ�%^}��`T������D�\��CKR�i�ձ�r$oW=¥6��٭"��l�&���!B) ���Pv2V/��?�"��$� ���T��D�җ"7�5
;:Ъ�z���wDK���s�w>�kK�?�N�+3ת�C���]n'>�M6�=�c��+����?v�ag]�lc�y(X�v!D�� ޾�iKtƓ���6E�������M�6q�ٿނ�����{�+c��4�Y[�gS]m2�X�7�[������"V6�~d�?�d���%��)���m^A�A�����Ͱ���u7I7�D8Ī�s<�\������{�(�j,��	_��7����c�Xp��ݐ"=X ����7��ړ(��D �,�=��w�Zk���s!iǔ�y��!��?���J�;=�|N�f�� �K�`��f	�>t[��;����w���q[+n"��ۀ�歍5�t��Ӈ��'�%��C�j��m^�.l�
s�l���3JK����w��F&|�`ф6,IB����&��;���b����V׈$E����EeC��UE#���c!_Xs��+<V��Mu�N�Z����	�֪�]��j�t�'���!]�v��;hn���0P1�q`�sd�-ϡd����2����N��	 �egf8�&�������kf;�����S�8���U�_���,�U�}�1"fS�C��}�Յ�����{^�qG��p�kꯚs����f�H�'�Kz�s�T�:p ��@�=���N+߫H��@�JԱؖ�j�Ms�O�� C`0��8 ��=��@go}����4` ����l߇I5�Ѫ(�>�/�W�����{3:3�h�d��r��J5��Y$���^�ޙzw,c���Ȳ�b���ɺ�x�F�� �뢒�)�.V�C�ssD�dO��S���D�e�~��@:����T1j�� ���'�,��&#ӫ�-6�d��<�y��!���ġ��$��B�x�2�ؠV��1�C�%4�f|��᫄J:�$���p��/���!O&����Z=�ўhA�Lx��z��wl�z�*Yp],u�<L���*a �S	��K(�m��,y��{�l"�L.{��ͳ=!SMܐ `ˊ[x��*�-9�
WH1f^#�����9\��4b��߳/��J�!�,/��8�ip��2�Pي$K�3�[��-�r@Q^4ח�Bj�F�(��cR��{�� ����l �sK36W(�k�"V�F�8��]W�x�8y]��O���p�Bڼ�҅�	/�:�=��DOF�x\�pk8�z�}({إ�E�`J���,Bn�!�s1)�և�����7���+���a��0ۯ��-Γx�6��t�v`�8��~	qJ��$�Ζ�`�^�PH���� Ѷ��l�v5B�|<,��
�
^�7jaXFX�+̸�뼆<��s;p�s$�������ҫr�3d� ���<*)�g�2[W�E�������2�jy�]��P��J�@�~O%���Nzmj��be_�{��d16��ký��ՏS�1�$�����F@��{q}e,M����}C�L�K�� �A�~�<�a������k^�7���-�q�O�Q���dBVz��uX6��n�}���*S�"�7�:�<�O�n��m&l�8���I������@�v|�r�mI����Ifo|�;{*"�'tl�����x�C��HMMٱ��D´����AX�68"�r�
��ɧ��F#\����qa�R�[4�1qD�g���XY��a��ZJ�d-�~��5s������~� �g�#�1�65���K�����������N��`�̕�`�j�n����场���He�B�J�y�t�#�ϵS�����n��R�K���
��M���F��L�n��.j^оS%=,�K
A8vH$+'�ԛ,Qh@5�Z�����L�~0*#�(x4Q�u~�|�P������V���,>�N�׎=Ť/��/�|ώ9U�f�?,2���7dc��Nbh/^4�ǅ�����,yo#�G��T9���m}2�ߦZ���6V�
�T&���k�k���� J�J���GZU��J8k��4�wz�T���Аh;�p�j�gkQ�v��ƾ�$ �q��;��!C�	���W&B�{�!xn�P��h�]����N� 2r�X�K+Pl䯋�!��;�0_&4��t���>m.����}�3S�qu��n�e%��YʮD�D���{���N߆�;��}�-��Xǐ3��TM�4�V�vΡ\�Hv��ˍ���\RR8�I����)�w�����ι,�8=�9	桖�%:�z��\�w(�#���8�с:C�:g,��<q����R����)�E4+:(���J�U�d�u�`���"CW(>\��ݺ������*��md#͎QP�{�h<Xغ��5��h��!����0'�����h�
���!�2A��els9i4)��I�0&���P�����/Z�7���� p��!ۨW6ɥ���#W��b�1;��2��e<�Et�G������(��1-�ң����1������
����wψ��8��],���m�v^"B�u�f���]��hˑ��%��Y��Y �����Xg��,4�gyDo�'�VN�H���RV��zh���G葉a������&5ܾl��Y~78~J�ɤ]̉5ҭy�Mw(q�����p�	9GY�DKqN��@sua7�<��?!��.����D,���;�C����.-٩@�V�G�|�����]�Sm���&	����IJ��6�>JA*�1���͐���i0S�\Z�=��[;ʃ���'G����S�������%U=e:�d��w�o�`dψ��7�� ����V���Ǭ	�N�^�<I��j�5��o\���kZp�6����v�?�����喀�H��A�"�t7'�dZ��tI��N��{���Z��k�����~Z�_g�	^�V'p��|'���%�������yΑ�&���PCƠH΂�b�vB��ڋ٤d(�'5:�^�J�Lx�e��$I�@}����O���J�.�`���(3��@�۪��\3�9�
������dպ5�2����	[_��-KDP�
�Z���wy�Nn�ɻs7�u��+&
:��?�?�Uu/����K�u,
Z�x�Ɛ�\���R����/��!��8����
�Ln1��\V��]BSdjL��{ɟf�G'��9�1�h� h��v�K�P#t)��D�
��B�1��,��f��H�4��o+����7���wڒ_������
�#��1қ�f�
w���؇�o>̉y�,����<���1�~I�M��s$��1��p@w���fu���J��,���$�ވ#���XBVI\�4��8\#�����b��G'�T�N� Z��H�wD�������
�Ƨ���
ni�ګ�1%���pP�3I�5ΙY�U	�(�jlݒ�3����R`A� '(Z�q
���"pa�C��i��+�u�$V��);'����0|���m'xS���,�����s�L��{�Ɛ�+��C��	zk�H@��:gV��;��N�t��ɠN@QD��4}�~����@���O�B_pt�Hu{(��њ# |��Lz��~���&:Ki�N���֘_��hfs� �ߐ�5��1P0� ��Ur��}�T���_���ACQ�$Ş��X�B�� 'DR��E�����|y����P?�$Z\�.�/4)�]؂qA��@�.�Y����UY�e`ЬopA�\��Rَ	dd�LX7A�l��}��١߂i~�.�4�w>T�);:>�֑�k*1���4�M�68&s\|�����K \>^SGh�*9 O;]7���i �}9�Ng����	�NJy���U�\9@\�Jݰ���MA>�+�Ӄ<�VI�&��V�b���GT$�Н�'�\y������ZD�͓7#���X#N��Uo!	��_>Z<s�W!q��;������*2�i�w8NO�W�8GJs�jv��m;�j��4Ղh�I���$�C���<q�(fRjlY���J'�0L�ɉ�^�JQ����L�#o�lֶEߛ�<J���n)q�q�b���\����c)���MU �$9��#�?-�gյ�C[zMl�ٱc6�㓵�S�@IHI��G�x�E17��ɗ�(���R�2-F��B�6X��];�_�{S�8��d�w��u����1R�~�8ިz-&�,�6!x�V����?u�$�Β�ƈSF?��T ����#�Xg޾�O^���ŀ�m�P���|}H��0���cw{���E%S �§�eow!����o�mq}�*��]*�TU����ǚ���~Δ8��]j�k!��V��.�LxY�@&�a�X~��b(��V��V�����\<�)~	���7ANԹ��/(,��R��`����8J�F�p����wA��8��~}6+;��)/�E^2��s�jB� ����>\����DT��0Q��п��Ep��z�cX=$"�Og���s�ι��>�E�[H�����ޅ�N�c�
��^�<���*A�����r��^0�4��� �O�ȫ�\-�irrͨ��Y�6^A}�u�N���lWd�%K��)#�%��AG�Ԫ ���X_��
��򾹊�f��V:�U�z7d�t�r�yП���n�{F�1��:����m���.�}��!
��* �T���蘥�m��&{��;I�7��g6�Kk�;ݲ]�Z��� �$R�-ŏ�P��qT�1�*�RS��4���&na��"*@%Mo8{�<���j9]���ܻ��.}R�虖�~���J'�@������35�Q�=��Jt<T���5��}Xa��綜M(��j��.�ζL��qo��������N�l_��@�wS0��䱬�t*Ъ�)����{�&�gt2o�B��a�R����q�dC`�C��G��kp���txx�x˫��O}�j�g��.����]����>�H�D��9���5��.e��]X���$�k�]TuQ쬒��)Qق�e��R�<T
r�������l��H[M��c��(ᘌZ��՞|\��<��%����S�;&ڴI�I"��,�'*J��3T�L�����قp�m����(��`�,^����q�&>?�z$JX����]�V�%���6�S/k�/��W���!��k�ɿ�zSB�?���ƍ��VÑ#�����ry�?!*�����7��/�r�k1܇��)/F��G�Tf&�~wz&Paզ�!`z���;��B�����i.nt=0n�!�q%Ԥ��sW�챂q�(K�x��*!ϒ��Ϛ�4�bY]y�G�p&Rǘb��2!�L�g���Vg�Ƒ�̵��}#Q�����|�q�r.�(����K]��ʦY�f	��U8v] ����H�.�Ýlg���������yn'����m3EQ�T��M<Ҁ�#��b�W�>C�9aB��o����cKq
�vL����ڴ�)��[ܐ�j]k�:oʒ����0Y:W�5�Ï��Dt��H!��%.S�0\���&��e���~%ܡ�G�''����`@��v �#S��JQ�B�#n���aL{X!�����*j Q�6���-�^��4NJ�M��X���G7��'��mv#z�H�nU������A���W[��}��|Qp2����C��S�!8�#��趟٧��Q��W�V��DVk�>{�q���CO������O_��Y��kLID+�֝�}��{{��+[	�:��3����G�3���S�+ާT��	�c7�O4Nf�QQ�,��q ���?�>�Ë��r�qR���!:��>���;�
��~�_��'�e3��	��&��AUe�KAjeL���x�e.�T9�7	��Ϡ�q>D��\���!��f�]O�a���n~s4$d��G��̚�# ��c1�x�$ʓ� �?���Qj%E��I�z����.�$tʯ���ee����/t�x9P�C��ę��:�%S��V����]��a���I}v��:���p�Y�:��A�9�hpf��s*~p}>�ՠ��a���i�LY)��5��ny�C&ū��
�r��l�\k���3�7e`�Wj�D�j�<@�eI*���f���£��~��XG�>���oaj�&�������5�c�%�u
���bh��O�lc��~���ڌ3�*,�R�O�gn[=��������� �#���,w�,���ӔɧJ�H����g��T�����V0&���N�G#��	oQ%K:�� �V/��?=@�3��1d��C��}Q�䴏F�N$�br[XY�}��FwR ���36��4Q�G�}t��N���ĥ�b�i��;�yZ %*95��|�dq���*dgPS���K��A�1�@�ؒ��%h���H8����)l�w��~dY�\IX�>%ׂR�-�V�pl��� C<�O�)�c��
��p �R���qF��7�|�F���?���N����~m�k1�f�)�g@�=2�t׷;��k����6&<��8k��	"AvV�����Eq�"�qNl�!yCJ塌�M =���)_#fGwJ/�ZJ���+R}l�@:�c|����W�L��Q�3����[&�d�(ڄ��y��b�&[-B�ϟia=q��/I�#�x���n^���HT�9�e�{l" �f�agni��o��Β����4�̈́��<��*�[���࿠M�Av�p���Y�k9Xl)���]�ϫ�z�]�����U�j�H��Nu�}-��f������Tx\���5�!zHW�f��Y�KTc1����H�ur�Zk�ǃ/U皚G`�}�δ}�_�$]�Fb�b��#�����c��4�gig��Y��M/���	�����%whMr� #��sFV6��y<7`G���V�J]�![�C�����@)��t�I��rKz�#LØA��N�� �!�wo�$�� �e�(B$�b>�hZ�9߀��.B/�%8�q��:�4�WX�~�i,������tk��	��(���+`��PvSw��v�Յ��CDD��)	���:�%&ϖ�;u��1�`�(g�KB4�	D��m��i>�}S-}t^�W�52�S������;�S%���2n���t�d?e4��4zT�`�H�4α*0 ��i
��\�tTÖg&���d��� `Jf�4n��z\t(G����'��L`/�B=�W��7t��<k�жO�%кD�0���B�5��~ɭ;e����tnG�ٕ�J��n~���ⰨȪ�����V"�Y<��Z�����&u'�[���y��T�ۖ�{����4��=�2(=��p�,x*5yt℥��I)�mdP�oTI��+���J�I��:�cu�F��p��|j��ׂ	u�7�=���碶����.��a�� �ۘ%׾��:�V��1��u��[�/�k!z<�G|�|KQ�0B���~.�:�jp�X���	�1�H[yog�Ƅ�s�Cv��Zz�kWTD;�t��{�pY[�k�go���n��CSK2*�� ���˸���E��q�ޭ3Z�,jTw�qFڡt$��r,?��{�y��'H;!F>���B5T��Mt�wW����PYb.5�$�T4A�%�/:��c��e��J��ŭ>O~����#��2��E���%TdЇ�/���L'�C�yʱ��]б��wePL�"e�=.Q�L-�b�?*TZ��"�>la�o]�u�+�@�]�!P���8�7�#��5WehN�D�b��GZF9�H�/�L9f�΄�^XUa�Dl���W��Cǒ�,w�Ǥ�#�`�!����)�H��k���cגP���#��"���lFe���r��^|[ߧMI|	j�ݙ *m��_;e@K��]��8���br�������J�k�o��?[h�x�L������u*14.��b�����{���[�3W��k��N������K����z�E��0Wa����&�"v.w,�$E�m�Gq��Ds��L7�;CH�p@IQ'�0f�w��=���8��Y���rЀJ�'�@Z�	�ZŻ��Z�pWYD0@E��6jL�b�;��@������	������9����?���T�W��ZT;;�^�]#��ǫ�D�D�;�z�������DK�̴Е	E�t˹��W��sLa��!��'�n�>��	xhn�o<p��Ȱ�u���&����p�>%�(ՠ^����=m�8|v��2�A���'�JF6�X���	@����x7y��Q",AU�`N�|<������.~��|dI}�lp��TV�Ӷ1������j�<��KI\�'�9�[Q�c��O��q3����Wa򢓣%��H*�Ct!J�XU�s����Խ���&(ʙV�ůSU�ۥ-L� $i:t#���H�4=��xR}9�a�- ������D��$���/S�os���r;�A�~��F�.��ZlQ��?k�"��q}=�Z�1�u�W�7�2Q�^B�����1D��1�P	?+��['{a%�:9ژ�*Y-����&��{֎2\$�z�\�6����2�J�m�J���H��P
��m���Z� Ca-����bg�*�T4�������eI<�P�tԛw��>Ø)[�����z� �,?LN2�J�����L�n�X�/�&�� ���+�:J��c�&;�G5��D���0�������T0�g��ɹ�34��u��{.l\̴���':}z�	 �����( È#�lD���fN��=�����\DPo���֗�����G�ސ@s�����S>G�����J)�b���Pn� ���{>!Ľ֟���4�VI�4W_{J<�q%�}��ÜֶR����v�����J����#&SWr�ݤ5�h>B\	�{�%���ln�� �ܰy�� ë�vF�O����+d����{�U�P2�ܳ�S��x�O��e;��+S^xD���@�s��V�X
ȧ��T�/�n�P$ɛ�e����..OQ���=��4N�1^���a�����q��	2��jrLQ=6�OI4o�2C�Y �s�ҎY3}���h�,ݬ��x���]���Lރ�G��W�����G�#�U��:������I��2ϮcO&���3�R߄�bFb7��i�FՕ�%�0/rvazC��I�E"���VP�n�?��c.�ަ͟��!����"�� �Koj`�, ��:���c����vJ��$xX���g�w���k)[l#�t��/��}��Q��ֵ�{LxJ�Nջ�]�hWz�E8�IW0���$ۙJ|3�p��р���K�!��s�9(�c�](��Y�&;���`���%��h�|�`v�ሇ���j�-W#�%ڽ�������@M��)����f)[�QZ��{5�(����RU�W��l�S��v���P�K��|p��Y�Klh��u����i��&|Y�6
�(�kk�z�\f���
��7��xof"��2*�ҩF��a߯���ڎKs@���%F�p�y�F�X(�HXJnJRB$<�l�M��hٔ�f[rw������N���#G���P�Q��w��Wj,hF+6eՙ�/R*1V�l@�*�#�;VB����S0Y�C0so<jn�IpH��Ef'��%ʣ0	���q���U{�(g�c�"�#H�-f���=M�K�n#�՝��,J�kJ%!�|�����a��'`�B$��Y�/f�*�J�N���S3sQ�s�8��K��w����jJs}�E���s���v(N��lz�4p��1�m��	/�Ó�Y��q&�
S{���-������OZP�M<
�˲�6W�mR�݈���!k�����6��a�Kl�B����~ϝ��%A�6@T��xX�ٝ12�S}�Bj��
��C�/ 8�Ë�.N�S��E�Q�챷�T��ۆ���� ې)q�6�N�ʒ5m�Ҷ<-Z>������d�����X��� ���S�'���A�J�F�Ӎ�F�{������P,��u�KV�#W����]I��ChEڸy���n	�ėi�wp��#-c�����$>1�a�
�X����~f��D��T+����9s��Wp�i�`x�����YV��7�)��\��b�|�����x*�����%=I��*�و��9�|�&�Q�6� �S�X�E�>��WM��@x�/�<o�'�uaSP���5n�tQ��ˠ%@Ю%�.�P�׻���؏���4,�~q >������Ӡo����Q��eA�a��z�L��5�&�.��}������1���}�:��>�T7�n4c��p_�ֱ�\�vi���h���F\�_������^q?�c��{X��۹W2��F+�&��rG3Dzul�C���bd8�7�Aj���5��F�U��̬v�C�^���ªLJK%�;c9�#��	Xm���]I�=�rj7)l�~�M�3�eQ��W_+�`�F�כ�XԾ��7n�e�!��;��p�o)=�w��n$,�&�ze\�tP�H��8"o[�ߢ�.j���Sd'��@Bq��*��BL��W��F`�yR�|���}6~r�ct9�?�](�4�j��ex�
�1�?\p�K��1α�`:�L06���Ыߤ����޻JU��������6��r�D�	gE{q;At"U�\���3�$��րH#i۽:.��G~6�x�;�n�YZ��o��՗ɮ����Z:��j{���c��E��-�2{n.�`S�>�y&��H�u�lA)$陘^c���]*�Ύ����x�+�[��Ry��k�b��l��j~s�P�S�̰`J�T�L����!�z�vh�ĺ7�c}�r��	�vW�f��>u�(�k�ۻ��:��j���ù�M�G��1̥��pP�ۣ��;��X���mn�(�\.K1�t��U$]j�t��#�`1]nXcDw��qjC�.Y�P�L�rP���Xx��;[��c�w`�6xr��0
M�H�\*s<@�-���L�6rܬ�ܽ4�.@Z\��"�Y��}`c�9fܨ{��Ymx�\@ᯃ���S�)4��@��(�Kn���)�^9XI�� Ue�}�ܨ��=�:��d$ѝ���=�O[( �֊/�գ x8̈A1�f�0"�F�r��~�?�_K�(��\<����yE��ŅV�=U��#U��asG	L(B�L{,���W��GiN���%(_���
�~N��Tn����L�SZ��n�c"`oD�z%�g&�=����_�I�B�n��L��7_�|3ׯ�-�g��L��0&)-��%�3��#z�����Fz=��$m�r��z�ׅ`�R�TT���fa��,r(�������8�G�����u���HvZ��2x*�����V�F����9L&��d��I�f�VJ�m0����5\��4�� �q,�[�F��bX��#������ _��v��z:�ʑ�0��,=}T��R��B����]�h
�S$����R'�h�>�v�Jl,q�`R�v��	��ΕnҫH&<0��R�g,"o��*������ Ϋ������Q�ф���ڐ�eV 0�/��/����m�	=�>��r�~���>m�'i\��-��s����Ȃk��rmp�St��@�E��WM�G�&�;����<�t#����f
�ّh�V|C����.��#:�ûuj�j]�ݿ]����K�+��������e"�jg����U�;ښ3ښ�QUj�X: DO"�qj��\��|lt���\��G������ñk�" '�gܟ�K�w6j�GI�ɯD�J�5�B�HiCr��EQ�d��0P`<�����-��h�@�6��u��=��	J���ϕ@�41�,-觛�ϒe?<�����c2+i�-fY�c���_}	���LE|�rͮk��B[����\�X�@�{|gB�j��8��ȐA������m��
lp19{pT�y�:���W����|r�D�����&rl�����H��z|�󥛭�g]M�e�ACծ���,}l}LZh �R���.�7;�u&��sa�
�����^n�Mַ��˹4U/Ļ,�ڞBU+�I�PWTJ!��Kj��m�:���~M�^ �~�>G�]r �!�B=M��!�dl8m=�ۼ��ҋԯe��ۖ���
�ZV��2�L?vqH�]�4�J�ąX�tݡ��-�K�X�O������K�����<G7U�8t�Q�d��;6C��p��^�ɥ�h\����ZQD�||��f���3�q�'h�B���S�������K�gdj�GiЂg9Dw\��':3p��tOB+&a��0�{�瀏�fw�|�Em�1��T�Z>g\Dc�9R�(M����ц��o-y��}�Dn�Y�i+�%-V���R�FrzE��,�u�����[� n��!��.F:��C���ʽ@K�;ŭ'��d���������`6�jn6&l|��r��Z��)���Q���{�IRE$l����;����J���{��e�y��������@���ί<>ִ/6��b!	C� ��H�IF�R��.��'ކ�5�����å�����8��4Yg��4R�;�p8��⇨!�ś��q���M�Ȱ���$,�ݖ�!�1I͜W��*�󇅡���ųj`�cJ�9��VW`|J角v���C?�w����9a��l���Rݸ�ʱ�
'Y�Y*T�!�ȍt�n�+X]�KԲ��F/>�����F�[Q j��V:C���S{�> ��C��y\v�,xFMD�h�p#�hUf�������!�jg���5lL�V/I��5�g<�-5v蓎�P�o#}�Z�@�D��=A{1^Q/{t�/̙�Թ�w`s��vX��^;"�^�(>���/D�-�bx����c�_��s��زi�R�m�7�rO'��Um��.�J�`56)Z���u#Z5T��or�7�E�_�!ΐ1�dA���$Yz�gpT��8B4�sΊ��ҏ_[p�yp8iX��.9f�`<�\�2���|��13�w�fE At�zaL�S.��,����YSʈs�� }�߯7���kH鎫1ĀwY����~����TʮNp(��z��h0Fp��<�\���i5$���'��8Pمf��c����u�T$�t1�_].��Y-��J�ENk�A����< #-٘oi%�"��y�7�\YMQy�u����	����m���L؇}���n�XϏ�|�b�H�F'�d�"�ɶ���&��B�~LZ!��pF��D�%I�f�u��I���}#������v��JSƊ�ZM�зH�(�t�	���D����x.w�/x�a�ux�ez�T����&��^-�E&�2P��y:At�V�"F�Q����(�ٙ����M�Z7��-l�?���	Q��i]�w��&��G���r���I���n�ߥAn���>G�}��r�0���)�[��etcj���m���
�9�2"hM�M�Ϥ)�%*=U=�=RA�X��3��?���k2�k `0��#���1N"��N�ׯ-AZWi&��NO��,�����|����Ķ��<W��>�	;ڏ5��V��|P�v$@�46�%7_ź��"�
t���1�|v��6�{��-�Q�f5mb'rP�=�V��	`*�8���T�j|S�I�r�5?�"�b���%T����)X���d8�'���(16�����M���ŷj.R�"8�_��j��0�Ns��l��j�U8K�?C��~�T�Q9Qq��U� j�Yg_�^w'��c.g���z�'�u8;S"�@;��샺�7��|�2WI�o���:�y<zGӱ�U҂� 8�&	�1=�p�Z����\~�@y]����O��e�9T]��92�����M��Q��f�iı#1��kރ5L�=�>+
�T�(d��A�K�Ρ�}����]�F���{`���o�D+
�M�R|�(�w�l�E�%4NG�-/�xK^�X@s��b� '�z6�)�1g$ΰ>A�x����N%	�
��d�C���QOS�a���l�,U�������8^�@�@y�\_��2�+՟�����b:�:����Z�È�aV�++	bϋ�����~��x�vS�Iz�K��$��.�c�q�}���4D��8��g��C�\�~�<6,jG�f���ߋ~	ӟ��2�.L�=s�4
ĥE=Ԗ�#�x.������ĦC��m<h�;&��z;�G�bN���͕�<��n���|��ޞ�rmև+�4fǏ�W���G]PT5�KL�@D
���Z���r�ᕬ�ʲѥ���-C��,�H�X��\l���A՟
���؅��y[$��qr��lM\t? ���Ԍ�V�Gz�p�~��ʊ�|%��e�~�z�E��A=�Bo�3���$x���n���c@��W���0���V�^d|��5K��S�/��(7��-v���7�ˉ���\�u�9̧F�TM=:�U��a�H]�4Fe���R�b�҂5n*&��p�4���}�٪�ݘ}�z�I�[�qX[��o�Z���;����zQ�>؉�qb�X~��&yf��W|;����8���#K�)۩�|ghR��Y�[�g{��+2%������"�C����m=H�l�/����ߊ��U@''oY���ߔ��QÒ;/�d���d4O�Dr;:��:e�B�АQ�J��C�Q���#Avd��]d�-����s�w�+8O܍��<p�{1�K�?�d#���2%E�qm�6qu=��������Ut�U���_�J��laV��9��sScu�0�Z�h0�IH��Ӌ�Sr�+{�'��!B����w��&�q�Y{g�끡� l�Nr��so��uJ ��r��ݠ�~{��iNx��~��R�X���H�U�u��*�=�
3µ^��4N��J���k1�$��v��#�Yۻ��0߀Nb:q��l����4�c�Cb���E�v�?��F���Z5I�ǧ��? l�g���c8J�k���P*�<�n�g���"��Ȕ���#�n#ɜ��B�bgV�1.ֿ=�8��g�:�+���\(!�!vn福L��l����\��v]�)1�;h����J��h�� �B�ai���%��{�5)�p���0-"]J�O53��Og�Y�q�x\>v�~]��v�V9��ھO����i���g��ڿ�~'�����-W��T��������	8"�����O{^O2�4�� ���tУ�!�����z��0�g��?Ec�v"&u�c8 ��MDT���i8�1̄�C<_���z-���V;i�����^��R)�Fv�\T��n`��~�%����۠$�v�ys�M7$z�S+���KK�����~s��v�=9��;%��pI}�e%�>�%b��r�R���nh��e����W�:�˯����d���Ap�H�,8*[�j���BD2���pr��]��^�����x��#m��`��7j�*(����2�$ޒH��$L����'���n=��x7!؃�]�~Ի�Z�Df����M&F���f�c���;��ҁ�ֈSq�d��+ +V���㥭ω�ߖҜW�g��'O�c��G���3wׇfB�X��ϑ���lbL�f�L�]��c���z�H1���;F�3҉y(���އ7�6��}�L�b���q��X�S��	֭����	@\�:dя)�\Z�h��Mj��^�P1FE鿃�݌ޏ�́��s}��)p��F��A/���^6�;V��i�2]s��Q�.��2���QS�-�ϢJm���r6hK����2K����X/nL��9v����J���P�|?�g�!g���'��[������ҙ}Qs�~��B�H�N� ��x��B� -��E'�_����Hr\1�&���&�N�`�$��-Y���/�*�̧�����jC���x�U'�Ff��Wy���ֈ������BL��1�&�Z��4��:���P��}��\,DQ����ag�A��M5�n�����6(��[ո`�f�9r^�]YZ�I��Su��biWs�t�.�ѷ��Ť̄�ǔn�������Ҹ�+C�����g�)\�2����sH��9{�gH=�Y��6>��1�q\)����e�,C=�|F�qZ�%#|�8q���C�F V�'N0��b�gQ�u�i嘣�5���sJ.��d�K07��9�F4bZ !+�9���ι�j����2��7zCpf����o�@���.��'n�D�*ʧޫ0�|Θ�l�Y���P �?���	ZK�)ͨTm����,���,��&kZv�hRql�̎Dw5�[-B�&^w�'l���������,�݂{�� ����I˵
��㼩����<:�!��UiiDQ�P���Hb��3"#r�a��������OcG���9�"	n�u>#�
;�+Ũl���E��YI��_;T���ק�'�ц�8ߙ��@�&�����Nxڳzkm�zaO!�������'8=n��*C�*#5�zI@��W�䏻�����>bO5JM�����0����i�9Yy�����'�V�G�/�%v〳�'G�dB	��{/4�JKw���o�=O�J�h�߲�vI3m�ÿ����}�*��׉�4Ŀ	�z���E}�;���'\ te'���̦6I��t�wJ��Ǭ�	R����q��4OH{���m�´�o��>�e`{g����R���ʥ���1ޜ=p�)�0�[�bX����w�T�!SE� Vc��q�~~k��T�`�ȷ�ņ��:D�SRJ��X�{^�H\ �I���vl����ir���c�Ix�p����<�CM�U�0�R
����6�p�x�/tڕq�nIQ� \A�w_*�ǩCR�d�`���lo��g�t��)�8B����Yw�0]�$�ͻ	x���fo�[W�II-#�rcܬbo����| �E�)��_3~�9D���U&�~�T������'x���w ��
::���W9��o�a���Y�
)��9�\�:Ѹ�v�ㇻ/��<�~��]m9>z�Q��7��6҇D܇dt�`o1��8yV!z�PKC�"X^v+��V��^��\o`���G��g���y�'H�|W�.[nl�e�V����"�u����*[����򎡯e�6w$�@�a��%����^U\���nm@c\�T��`�%������(Vu0�[����p^o@ap�b���7�G�̝v��@��Z�W�w$�X7,��6?˓�����'Ց��b<g���=�:м�YGo@Ѧ}�HH�X�aW����Pe���� ���3�|�\�|>��h���b�x���V�}� ��z�0q�~�&�_Ȓ@�W)��u�'z��{�.$%�������A��5E��e~χ������7��\������ ��&g�6e-Ps�+��m+��9�j̧ۜ�e$?���	���ƀ;G�Ʃ���$Y����R�g�����j��(~�uu�s��b3=�Ȁ���Z�/{��{j�,�*b�i�U��&{�׭4+�3|٤ڍ�E��27i�0LD�BdA&os{��湰ߕ�{��"���N�BDQphMF�'\p����n�E@mڮ�sj�o�~!�z!+zcT�j)�5M�uƯ�*���GA;z�%�&U.w�d|>�L�r�T�gj�~��N.��7��i@���zĦk�:<��k����綁q�;�s�A�`��%��$s�A��jQ��x�+*e5��7��o�#�f�f�[������ߔ�-wJ,�ҭE��9�i�bE}��|A�d/'�]���u��~���]O��y�GG����&snR���������F��j�l+2�2SBŠ�H���'hTY%]�h�@����#�����)$�"�W��#�]R�UCj���"�%!i%�0�N
�s�~Q'�a����՜���K������L��A�ƚZr6�����T�e��znQ�2���?ĸ�WnQ��t;��k^��(���9��>)~��~���|z<r��y!6���Y���ek�Cm�^�o��W�QQ7m��o�t:�fo���ˡd��|cv�O*g�,�w�_��C��a؄Vd�O���&#�$g;�%d�^�V��q��L4���B��c��i_E�k�p��K�'A\�Fߦ��rV+`&�����T�ɦ�����-f��I���j�� e�V�j:^�[edsR���" .n���=���J���_�������	T)M^��y���>oe�w�7n�Q�����]�DA�1�_e�jJ��gN�%S�y�R#��O��w���{��c���'�"m������C+��!y?� �W�d.��j��K{_؟'�+s9 �=�V�2��]��P����GOf�yQ>2�If��"Q�����y���r�Q�2���ɑ�;�����K�X���J�X�uF��7-�Uy#0�;c $425��o�pw����h�w�䲞L��t�(f�� ʀ���q�����4�|h�__k1�L�+���$=��"F�V�F�ԇ��/z�Ljy����]G[�J�dA����pF~{Y�f���Tn��[�k�)��Ǹ$X��O)dV�杂��P`�2�@U��lR�� �>k;��ڿRQ�ā�H��)v���JȓhO��W��K��{X����]�5{���w�84"rp$*K_p���Y㨣O�6��0u�<~ݥ���7v2�YZ�Hy��.��Q7�`�~Y��K��n�L�z����|y��.���UU𞶨�29B���3������e�گ��p�C��H�C��H����������˶�2Kg�p̜v����4�L���*o��u�{TO�^�T����M��ꝳ��ɹz�|��@�M�
��5�8�wq���ur7a�71��#Q˰�ȲN�h�[u�������������1�V�d�(��y��\�A�km����l�J�kRw�FL��t8�2.�n�q���� ���Z'" ��I8�t�����9�R&
�������g�+�eH�L0�fZf�rc��5�/R��z��>N�d�IF���l,���CV�8����	)�[b�0H��#���h^���NB�/�βm���"� ��kUh��
 (���[�S�6��{� �T�r���w'Q��މ�ē~����GX��Q�ޮ�����N#<G����_��"ɒe	7&��@�̟ۆr����k����z���O4��ȋN�Ae��D�����5�d�#�c����\�B��L��xj� �Zx��]��^�.�p�K�뮚���/DB�nX*���5�	��F.Q�b�Ϯ�H�-V�.�h9�T�-|lN�ZþZfw��m��V���l��Ú���z��t�����"�7*��i@�Z�N6Ϙ�(<��;$���yôA���J�!��M���a�$��q�#$-�z�Q̡`�ty��uG�f�R��,6����-�ϖu�yN�c�In}��]��p%\���q��l�L���MK��n2l��,�F�M���Q~�7u�si�B���i
A�q7O��vI}O�b�1����Սz�w���wwک��o�/v�H+��k l��fױ��?���]#�	��. �m��2�4"{�g̛�ֲo�a�4�~����B�0
%�Pht�v|�ߴ��Ћ3&L^/��O��	�*�Vݧ��t�� "����|�����Y[�B�G�����P�|��ɒAp�5X|��4F;�3�}?��Eq�H<_��]�5ʞ��:�����vS��O�]�m"�h;M_��m���!N�~�Q�z\�?��D�@0�x�=j�k�2��ˤ���l��Z�Xq�HB"&g(����[ ��VM�ʣj��=/g���c[ڣ�ţ�q���\T9U��V3��"yB�~��}���C��%o3x'4��;�
,\�-�<���R<��;N�8XÓy�/�}(y L��9�en��s���(v�/�@��âmG�B�:� ˙���C�!_Uc���yQ�z�*c�z��D�-���\m�p�fHd�Y�\�9�y���"Vy` A���S��M.�ɍ+�䳂�ov:S#^���t�uG�eF���9#�oap�"�ԥ�s���PΜ
#��?�K*
jp��0T�`�{�.��Y�L�D.B�%vVƾD�8���#š�6p�T�V�n�@�e������ؖ(���[�/��̄�6.lh����&�o>�/���7S:�S]��;V]�n}���^f�夞���+~���o��هN�_��9m�ou���j��4�����l�����o��8o3R~�A�4���>{�������Χ��@-�9dǅɚd�,�<�8Y�<�|��`�`�׹}�vڞ�7l���+.\b
w��`��'���5aGdL�-�������{��ж���oN�'��]��A����-���ʫ3T�F������g.�kzɺ��� l� ���;|�GS�yVM��ʶ��wܭ�=��Dݵ�M�7X�u)v")&/�@M15GC���h;�)�GyD�P��Ll�Yk�^����>�Qj��n@_5�b�x帇���	n-�q�'@zS�l7��%Y�3�q���0��J��* �Q#��C���uUE���	�
?>�x�nT����u��w�¾�Υ�/{Z,��n�Ϊ�?� �T��;�B������geK#ҧr��ȉd�c?}S��Je�|���7��� E�9Ex;��u�_Ʀ�G%�v����ʌsx�T[E�3 !�"���X���L�AΒnqC�t���r�S����2+��q]f��D� :ϻ�K��]��S!����NϿ,b���I�6�e�o�[G�ﵔB:���M[��ߓ,z��2�_
@�����I���p�R����{�V���[�.���C���+�MAZLÿ�-���p��>�1���R��F��wxX�t	X>��U|�)~�@Ǜ�,�h��5�,��Y�tVW�7��v��r糰�{	+a�Ə���U?�φ��8�\��2�8?�P�G���ʾ0!���X��رͬ�6P!��{�c$�]�zc�	�7.Z�cE��7���_�?�:Z��E۠W���·�]��	�l�ם�y�ɩ�m'wN��+ d��5���I�3Yϫ ��]&�/KJ��!>}��h_ܰ6��*w:&�w
w�T���<�P��	��'�X']%rp�U���OR�8-]a��D*�LF!L���)��0˫1u�ns�ya��.���DݏH�a����G�^�mOGu7��Œ=�{�͇w<�y1�4B���#8R4�O�8Uw�B�6��l�%ǆ��k  ������j��t��Ae�%uZ��qv��a���c6d�e-�%������ݞ=W=����C�g݀��%�SޝN`U�=]6Y(
e��V4���59�
�!�x�~"x�從��W�y�������>��牰��1�ejCy�q�V������M;l���֢n�'���>�	eu9ebG���Q�������[�m����˩	r/x0.�]/;0w2y�{L�,�}D���x��b#Gde������نC�}3��c�8���q+7.+�g�:E�N
���!Vz���,���
c�-
$�C���my��;P]z��*q�7?W����W�%�L�?����dY�G5�g2!�.��Fr�W�]ĉ���W��4j�}u �ek�	1H$+��4>�����ce$-w!��AV5���J���`��N9�sG�n|�~�C�s`YQgM��P�O��2а_M�T[Y
���a��KQ;���<C�1�Q��_�>@JO�䴘���UM�A�2�Zy�m������xܦj��e�y�5�s!�U|s�_�s�D�~ss�B�����4���%�Qu�2-p�?8��&YIJ�r|Zֹ�z��pC�Q6�逨>�����h�H=�}�D��h�$dsFG1���wۅ�b��0�BN�����m�5u޶�O�gV9�a����ﾊϚ l���R�nQ1������"�X9��c\aY0W��"�'�M�b�bvn�(`QR������m���:�Kfۙ_")�=�U;L�/|:���;�� �b��|������j�0#�W��f�w9 ��ɒˌ����0@	�c�+��p�EM
d�x��b���1����aU�c��	L aQ�6h!F���t�$A� D��!����,���6�?���`�s_v� `��޷AA״�'%d�P;�5قpGZB��6b�v��p 򻟿|rd��t_�'X	��4.@��_+�Y�]s��U�=v2��c A8snuVz�:~�yU����-
 ��Eחz�f�E���(�( p�.�=�L��D�L�IC���u��o��y)U�
�����Y0 ́��w��@q9��	��H��T����e~�������CQDk|M��<|I+{7Ȳ�'�F#k;1����^�����b"v��c�RD�:!R���U�Bi�1^Y�2ȇ��P����?�.�tw���c�]Wy�%��ҶJ���D�U�TN�����d�)C�eCƷc�����o����}�7�a���mE�yv���˳ϻ9M��!-�]�E!���7M������U��2S�bQp.�Z2�{j���w��$w�:6��8�rƛ7���`�V�5S��v�A(uf�}�7�u��h$�Y�ӯAI
I�,�2e;�}̿����0��5d��c,��wӹ���^l�
5�l��X�з��i����7~"	����֜SkU�+��E��/TO��T�Y�fS"�c'W����;K�az�����&���Z�Xl��B�,^�͋U��ҵ������#x��Y\[���nxݭ���ۃ��u��D6�$u��(2��!JL�$��$v*iz�[�ͨu�14�lL�pv�2�������v���sEt�OS�xk�?A[����y�
_!*���w+�(���H	X���z��A|i;!�x�Al�I�,-�o�D\
��I�ن�q��>��~������c}��/��b7�����Q����?�=V��-�!��i�b�M��u�mx�z���Y>�ޤ-�_���������$��<�q�b��S��>������\p�0�^��x�	�L��L��!�99T�#��r2��HȚ�F&�w���6{��4�lԂ�ڠނ��򜍋�9���"e|^^�`w�~ �Kt,�<7��YF���1bd�D�ҧ�ؔy��B�D_"���E eR���Km�����B���!��Lxq��k8�����1�Pi������T�)W?���6L�r6-�l���	j9��ݏ�\YE�L�W���49�J��>����	�S�Z��Qg	�͖2���UT˺�	B���y�0�����p0*���yY�1ۇ0�
��-ǗA+�8��<G���۝Y���S���_�2|��o�C$U�v�{;/Q�F�v$`�5٘�R�nR+�TC'�Y���vZ�r@��B	����xM�D�}� �6i��@�13��(�8W*9i��䢗,_�Q�qL	�d�NѠ�Ϡ8�{�V�4��XK�5K6����M\��J̟A�f\�PۄT/���3�U���@��ʧNL6@FVe"0`�������=WT�i���F�|�c�%0_�p>�|l`�c��ԡ����(Y4��+ �m�%��3[=h8�0o��"Q���f�A���ŝ�n��3r�TH�x��3��vI�T[���+Un��E
�6w��zh��,"��:-X�@�qq	F�N�[��0v���r��ݩk��ɘq���3(�C���KT����HeG�=C�
q��m��j��>ÛW��UJ�E\u��������T&M��Z�kPqzL��6�B��q�L[U��d9U>p��(_�g�H0����=S�����P�UT�*Z��Ho¯�"'ǭ�W��T �P�ȑ[y�E+-�-��6�U$��=׶vfu,�s�Յ ���,ἥ}W�G�hVwIj`�=�7�m�[��է�O��������-��~Q���]PH���@�kb����\)�(�4�&
�AQkvp�l0�׮���{y�:$v摈���Qp��);%�ε[�]Ԡ�q�e�,}(�#�HlS�w'Aj��7��_c��;Ќx����6��(�6�y=����a�z�+2y�Ө���m��9'�F��"��]y�׏��v<~}�i����q!�:MD��>F�T�[Ū<�¶��2�ٍk�]N��H�pEks�8O1�������E���M�d~�▯&Ea�*�o��v�i5�{�0�mm���Wf#�m�١��R���5�U	|<d�%H��+]��-��܀x��E[x�&�T��:���F�h�^mg!kw�h�Iy��UqA����B,��f�,�Ys��+�qT-��ZF�h��H�:[=��^8�\e��`���T��䷲�CL�bde���8�%�A���#G��8�E���Y��^���`�d�Jk��'���G5X6^�j��k�\�8�|��qG�i��@����e�S/q���8������Bw�\��n�N�f~8�:�73d�j�r���C��5Ʀ��%�+V�YjK���I4����d����{���r{
n_A�$<z�E���-�1`3��Vc(S��s���pr��v���gp�4���Pb;8@�5��HQ˰rg2�<��Y�+MM�v���s�2�h��������/@����n� �~}�}�\u�7�D~�U��hOUxSਖ�Ek��V]�<8�Js[�h�CcNƗ���Ў �\5���K�i�V��&�۲��Q�E�V�o�/�8���`�2�Q�WQQ/��IG���@�hN����Z��ou�Iu��2c�j��\/X��"_�LnXj�����0k�T� F��8�)߬>�GB��0& ��!oUSj{�u��QWL1x�����X�bPN�����F)�6��͠<�ΐ�%j�ݡ���:��� nrr����R���� ���\���:�Hf��l�!>жv�?�5�Z/�c�WuXё�N?p�d֘]�]�P��E20%�ԺWu9.�$�ӟ�I^peٗ4�Ϝx�V�+�L'*�BӬּ������T�/k�b%�9F�3RS�k��W��yt�&����3S%X@������-0穖�S!��%v��Ժ�]���I>.��"����_���QL'n}>ӂN��{4��#����D��A��k��$)q�axr����'�Ʌ��O=�/��[ `���g>@���uRt�\2��1x�r�}4hݗ7�<�)nŞ��k�ޕ�>�\��B!��\qU@����b��J�OP�Q$�w�>����[���b�����ٵ�y����ؕ���i���ۈX�������Skj�ʮ�<�fh�-$�����p�Ho��tb䫋ʸ^��Bp z�,�c�3�(@\zR��#�>��� R�X�fIoE�:����Q������\dA1(	�wb�+;Q:_qV5֑y�A������D��'N�!��\u�	Ⱥ�y�*q��Pu�����?�"�	��W�Qe	E7�%�3!Rv��+��H@�ɝRx��l�����)SoюϬgq���Wy�iZ��
G��K��bv�!��.�
C������LB�wܓ�AvF�ڟ�8+�~�m��v��`�.�XF�J>;�\	�T�N���>�Gi����ؚs|� �� 2T˺	�qH&k���s�O`��N����Y�������gw9��}��>�䆎��X:��;�9n��LDn�*���3ցaZv/ f��V�b�Y�A)o�I�Tv
�P�p@�TE#�B�>�XȦ�*�lݲK�����2Yo�G�uX�:P���L��\�}P�v9%z��#D���[�EJ0��hܼc�T����jY��vº�s�a�på��|��:�v1��l�u��>\�R����	ľ;O*`N������U�V�GeD�W�C���HR	�%�c�E֏"��uv��!�	�[���@\����h�u�T7^ӌ*�a?���W�Qg�]Y�9�Z9zZ�Q�.�$}��r�)�.LIv@>���ʩ������n�}�U��j�+��|�Q�`���^����
����`�_��SI���5�"g�"H�����q�(*do�����@x��s]����zz��(F����{`��jD6�S��D�09�Ƈ���I"���0��2�0L���� �F[�����6�������ٳ:?���E�CZz�)��I��}��� 8̑��%DRa#�/f�~#B���so3PHB���A�m�M��F{eCm��Wf�m� 놙ֽ�:��'�بW̗�Bg��()�`���L٠z����JU�j�{��v���6�#&�����������	Rb�>�?��b"?�fz�R�����8Jl������:�"٦U�L���Ddvx���µ@��䒠��9���b��W� �u���iQr�R�����G�-u����.<�'����5�BcH��V�	fs2]�Z�1���i2��,�OY��0�,��ʡ������F��CT��������Z�A?6 ^��Y�<p�JB�!8����>p�I{U*�N�Rgh��۲b��8!0a�8*Q�95�[��0��L��4�}�o��vy�".��!��@.������K�|�d2��/��N��ɒ�3������y� O�����Z��mN������*��fdɞ�6�y���#w��d�]j(��Y#
�ou��A��Mט0n�~4�`�:�M�Zڋe8kq�^s �tV���=�FbN�d��b�"���Ykf��� �)؟m	\��,d"�a�!IE�\���l�tT�mo�u�d�� �6�ĕ��qN�ɦѽX?�R�[x�*��x�RK[��La|>l$��P3ⷯB?��*��v��y���v�;AI��/���QIG���W�����&ڗ�g�(��3��%���V�1��:�>�ХH���d���`���h[�T��N�{~��ߞ;�h0���R���O���D�_�����$W/��U	Ǣ+�Z�,~o���u���Nri�>[�j�,�HOTnS�����/$�-����0������O�n������β�\�d��(�%��W|ڂ�I�4\f[c�S��D�e�`����֩v<�/1,{����pbX��o�<��;�����E�V������E`c���:l��q�����3D�H���Z"�X>�����gwln���}���/;q�O��kg"*l���!0=�U&�n����س�H��9l|雦���y�"4�A<�Dܹ�����%� 0E��棕�<�[�����K���)[ppE����[��zt��W242�	\�Y�{�VsѠ$�y!$���BdS+�6@��Dޥ1�({؉�h�zM�[��Z�&X�2��	�Bv"�C|.����RSÜ`��˧U�Q�W-�rBc���E�	{���x�|��0�F�\���l�W;v(|��ӌ�T��l�#5%.yt�KD]y�W����e4�Վ��d�%�7���6���� ����c	�G����t{j�zn=�=�3���'���I]�1���ul���A���sRv �x*f;�$I���m���m|h"���F�m���NT���0�����FZ�6�
����സ����髢m0��D���_	����/kh�C�˳�\[��)Z�
��(���R0ܾ�,���M\^F;}t���2�L'}���;�Ixq��'�	����j����=�ړ����,�3��wd��˞��~���Ƕ��:tTK��]����&.h�Z��Љm�Vh����: �Qa�\˸is��������6|��`���G���2�d���������>�r3�_�e�_m�!vb�QU�U�_P�`*�����ES��5mE�yT���nq�5�oO��b�@T��fM(�7�o�%��T�#˯��R��.>����&%�S�^�w|��У�>�a���.`-"�{7>�$�N/p�Y��/�.���b"���\�~g��&�&������1ϑ�{5�u�m�	镁:QL�(k�0Ǎ���9]'���+�͏�>�Fw��7��0?B����M]��Q"�$�)����`�d�.�0f��_���ӳ�=�O��4 �ǡs��e7�4�y��a����|`h�ee���������A]_�bKǯJ� dNWڅp����AoE�m6Q�B06N��횻���%��dfa#�3cC�m�w���|�@^&hf���6u�~�NT�T�Q��+I�?�����d��a��),�ҫ6*����k�ː���:G5`vI��:/�D�b�G=u\ʭj�c���B4�����ͰÈ�����$�&�f�3�CGx{�|��-�`��M:>ҚPkh"�}�J�c]6;���Rxa�(y;�\�^���,�vA>��^��Z�o�o������z��xK��C\a�,�?��!�2`��p�$4��Q2�7V`�-,������E��q����)�����͚��z{�rFGW ��g��,87)��?K���������U��&��~ s�s�fՒe��O�
�ݛћ+BG*��г+,�?a�m������&|�`̂�Q;��� -��	6�qd�i:���s�JUE�x�R�ZR���(�f-�P�	>�@3���t�k6�����5HG�Q~P�l�a��GOA��И��`<���1�%��x��Lpͯe�w�UX3�Y�Bw,�R�����1��R�}N���g��A��s?�u���c�L�<�JZ�U@�����-f�F^�U�J'BK��0�R�
J_1�M��5� rN��)^�6ͺj�8'5�/�𐍥?%��$e�W���l.��V�i5J�[�-���<��L�C�:���& +>*��і`=2��=��r]엺!�g#���q�l��w����qeШ('@}�퀦�~؁�����W�>�G\r�[S�_��V���aSP[����XmRC8Š:f��IF���������fY�T�9��>�mȻ]�a��/1��9;�UH�5!��t��lQ�{�l՟�\�Ⱥ���w���:Y��:B��F��HM�2�+��X��֔&���.)��}�0jT�)�	Z�
���Q@g�7M�<C�)Ԑ���D�
�oc���?�P� �w ��ƥߎ��%L��&
���bOM�]����q-t�wlv��ķ$3$��ǟ
c�'j2;��j�Jq�\��,!�N���r����rsoR���A��,����3���-p����\O �&zދ����;��:r2M�2���#ۚ��艴&E2M-�:��?�{P�夐��Nu�ٌ���
@�B�(�.k��h��e�]�p�.ܙoL��2 �2��A�x��eư�ץ��n�ԉ�bH���HN�R!�<]u�f\�d���ZM2#a��,D
ĕl�"2�nY�S=O�0����%�"Ϊ>I�{3a��v{�\��A���woTT���nNi'��AIף1ZJ.��4� ���b�Ђ�`����[?�Ap ���ѹ��iy��R��S%<a��<����`��d���F��;���ʪ���x\��i����@Q��W=�ɰӎû�.j�e����_ꄜ����y��u!t��?��'f9��8Ӡ���D#��H�ކd@RU�����k�A�������gE�Qzj$]��ӻ��%�,n��ۂ>m-(π������b���bw5���]&h�#c�X#!A%.��(9�E>�h�u�rF�y�$��:�Y�Di�z�FM�F�N\��Q=4v)e%n���p'0�$p1׎�̨��4.���|��^,M?��F0Ė��פ
T��/�p���sh�T�JL}���E%-~���N��j�n�K�L��CW���"}j�ɷ�aYX;�eϬk���FC�#�����że'"}0M.&���C������?�R��p��H�3g7��*�����h�B@9����Z��#�aF la ���y�݋-�>K���:/i13{����������lN��_"Pp+I��dr�""�?��s$��?�����T�}���-(H�^2W���j���H���@�xgě�?��ѱo[�~X������76`8��v�ީ��Zyxl�M6]���)�F���tHW �ט&63��20���[�b�6�7�T��/u٠Hо��;?t��0޲���U�4�q��B��y`A%u���E	�fyoz��$��)�byR2�H�
5�3V~K�������8���Oup<A��Z���/�<�r����r�I@���\��<(��BО��3�>��!��Ɵ��H�Mo�ᨽ��$���:�iy�Ȧ	�Ž��W������2�N��HSr�rn����x�uq�Ol�p�੠ B�S"�(	v��i��v��i�	Hij2�՝�5�����I
X��1��	�EPk=�I�qa�fE<��a���~��|�u�����^vh_� �1Tr#x���ಱ�h�=��N�/�o)�q&l�wc�.t���F�����L(+������{|��r����?�e�k�{��˛壔�oHv
3��*��b���Jߐ_b��.���Qy�B���i�0z��=�q"����t]��X���Q��@�@��+���R	��o��f�r��=l�����+�茛�l��A9�'^���x~��E���ےs'$�o��2�"��p�껭����Zκ���Z�����_���!�?�|��в
 =�r�{H��������ݖ�;�x�T�[���[/����	Ք/��sYI|Ԥ/ֿ J·'�#���;�u�E��,C�je�Rԝy;U�_���У{�:Ҭ��~H�?:*h���t\���H��!�������%?�S^��n�߮�F�ON���w�?��8M��ífҴ8S�?�6������F�0���c�u23T��7M<���#\Z˙{����Fu�����lXK��9���Lle�+K�oɉK}�'��yh�*�Z
�,��9�#S� ��Ô�o�����j�^�.@��X���G����u`�3��ȗ�	�������p�����7,G�����ȶtl�������CW}��IGM:Ϯw6ВtDڹL���ֻiZ��|��'�����Ǡ������8�t�ͽ_o����0I;�\,�BC�	Fi4Q#�f��j�Qa��v{7��̀�@tW�L3M�ݦV�����-����xbMO�G��s^8��r���d����8�͛ �Hn�sw{�G���)%m�?�$�33b��;�������A�xY�����jb�~$�n�C������`NO���r���K&1r)���v�/Jg���+�ʠeT1�(�΢ʌD�b�KP���G6� ��y��h] _���t���V۔˦@�|Ff.0�в	�v%���9�Y�hyàj�AD���Z=KdսeO�5�6�кݓ,Q���DD�0+[�9#C���^��I(��k�Y�cQ[��0��rkT_����۴'���ʯ��x�:]#�d��ڻ�eݟ `n+�io�K6s�� ���e������
��l���OS\�>y��IA GC&w��*)��ĶZb׌�"��+
�v�L�ۙ�R�H���9������"ٚ����m��y�k�P�+J`	���gB� �"�-<4��9�"$1|��'��ђ�$�����uK�.$�K��B��X��Gu�/^7�*�}�M?�#���	9���E�)oD���z��B9��m���g��&��<C����҈ѹ6`0w�?����9�N�L� �b �HT\���S�KLg�Ya�NUj��Dp��w��3�&���bY�9�c�6Ь��ʇ��M���.0\�<�9�^Pp����Q��)���JKȺn�m��LHx�+j��3�G�����:K�G�P�����_����,��6��E����.B�?� �̩y��V�w��E�-�~��]X6F&�WSmn�
x�]��"W�aSL�~�K|��P]Q8: ���w�t<��Hw�st<,����!80������L�.��u,˅n����E�m��~-��i���&"]&�a�J��Y�+�(!������>Ҽ-��&�{�����D�=q��8�����{�	�N��G ��#��}����~:�x�_~������F4,!0��U��n+��m`Rm5\kSpZ�jO+-`�F���X�pB�Ukϡ|�������	(-{am�!c�{���ɭ�ky�O��I�*�o��Q��/Btd%	qV;q�:B��=����#/���ؖ�O�@:��'hBw
3�9��/���w�/!JX�1��Sj�Itw�����	�#��C��_ˎ�s!j5iCP�>ˬ�8[�>���բw sh����N�Ɏ�
n��Ao��_�ge�g��gIs5�zq�i��3�~?�(x����k)J���s�����}�j&�5�I���Ԏ�>��:��t�T%>�Ѯ�V��4r���0�f�*��iaa�C�j%��KJ�ƌ��2�.�k�E֙�j�翊���7��dzQ�=��2m�]�Q��^fp�¼7��,�b� ِEac���i��v�����ުH��P�Gg�L>v���Ȳ
�u�V#�3��W!��y�WK�V��ϖk��H�r���"^.?��#?
j�9��4���5�P#�f(*��SȊ�y�	3Q�j��C'�2U��P�؊��I���x�J}N�.��.���5G!��I9�G�����e�������y��s�n*Ee�=�@�Us&d�RTB?���e���	��eG�]9$�C����I�x7?a�����ou �l$(������[z)�����
k~����/MKĚ�.;h�::&�<���,-�G	]��U��䜷���Ic��E���Z/t�F����8��97u!��`<q�.��L�iQ���W�Sblg
�)P�����_�h�(rJ(����꬛~i�t�JC*A�,?&'w�r���>%2{�YeH��}f��H^�()!$h�D��	MU��q1:5��UJ���lA�V�<���/��Է*��+ȰS���k���F���PHE���큽���h5q:���B�pZ\Q*�JMX��;@��W���)b�$�!��3t!��z��$r�5?����F��;5lX�恄;�[�!�m�_5P�&9��ynY�4Q«|�.0q�ɏ���O�@����VꝖ�$����.�!��v7I����;t�|Ӄ�O���%��g�v��f*�P,L������*QU��g��U��	a��(�A��S��C6ќ���3��Qv���r��N���j���ڦc'��綑>���ƻ���:�v.�eK�5o�IK9��-z^�S43��5��\��� >��K�Yr:��B�3�D��$9|��w<�O�?�FO|�4K@���?�lՒ"j�-kJO���n�".��	#F	����a~�	 r�\��4IO��A�r���QF�j`j�7���'DPt9]����,��T�����OP]��<�i�Fl����`5���?���z"��)�9���=}���V���>��Xw�`m�Ecq��m0;q"vP�Tg���4��d��ˢ[/psI�^���x����R,b���SO���k�����Y�F]�Ky;����Z
��5�<2�U��IGy1�Flㆸ�Q����h�K�nu�}��S��JLq����UX#�h��)zlG�N��4�\I��:��g�j# ���Dؐ*!�ڦ�5ec�g����E=�1V�yR�k��e�sɍ��D��-t��p�g��l�ڛ߈�ó�p�Z9p��ڈ�J���l?�B�i�0�/:��ώ�?�G�l��@{ʂ$&Lv�ڼ��b@��z��Jя���)�M��X�=Pu}X�:�ю�ń�?���� n���YZ4�ۮw�߮X���)`��{=����`8W���-+��ڸ=`�S�]����a�M���,_�������P�EXh؉�Y�dW��m������*��ʹb�{q���w���600I�����=��h�R��;|,"�H�*:��X��V�THA�o#M��R���2�Q$}�YN	���3��9	���� h�����VXqU������ŗ�P�'"�x���C:�IG��Y�q���ylT����F>�9���u��D'ǉwm��8�I�w8��u3^��s��v�B�oS�m���%��8�>X� �n���yV��t��+�'p'��j�<:n2� ���V�d>�Lm1�3�EŸ�!�'�x�<�9RF��l�;L"F����7�H�dp�W'�R%�,+�O�[���Sh8l��F����dH �N�t{�;��Pp�߀x�����2��l(mX�z�_���l\�ؾ��n$���to�~1�8��}�CnDY��xB6:I�%��yB)Y� ���Tt�\���1>BZ�h>��|�φ纟�P���VJd{�"��Ps*��tG���&p��E��ŏ.[a���|56X��J��ç~��Q=b_1&���L
����fV�%��������IjNNVUP*�ٖ�%B�(��U���y�bj��,c�@l�7rL4�l4Q¾�����g�~@���.Y=��z�&�>�O��qy�j������cHv���aO����^����J�G��fd&=���m��U����"����C@��������J�S�܎�4����3F���2G�nY�Ԑx��:��p����}A�Tt0�ސ�`�8��l��O$bx�l'�s蜇�$��ң�� ~)v-�!�I�Š7������0W�h*�'	&!����JjJV�\1I�v�U�o�Lj\dQG¸f5|{;���i�C��n�K�r�yS�h���-�O�us%������й%FB����pAZ�*C�����]0��9��ިM+hg�y�ǟ_/ز��x|g�J�g���b��O�	y�d����� yԔ|C&d�Ɣ�B�c7Ņ��5*L-USD����(�>����-�l�T����|^�����^jp�eL�>�%{�]8�"ٲz���)�E�(�څ�xT�1r�v�4}�N�R��J����p4��qm���%ֵ�z�Kw 54��c_ޕ��,P[d����������ѹZ��黵�Tc���B���>�5�i8�u�r~���뾏�E��r��r���[�b:7�����u�Ã�������j;8���7"�<K� (!5@����]�{Ibq{��d�'��}�To����HMU]��v�� R��,�U�
c��a�֚I��p��Y�|�1��_�{�s�1q==Y%���U���×Ks6+���?�$���q'��^��2<e�.w�4�[	��"������,X���jh"�h�獓��!����:��JY�xlv�n�#�����v7���c��6�¤/|L~�����S��y�|� <x.��؊Ėj|*ɣ��7u�_�uqL"�k� ���]Jۂ�H	���қ�^��7	��&�O��
��I3�@=j �<O\�a+ł����n6��`�jm�AF�D .�ِ�������!�Uk�M�w�~Q��,��,a��e�����hz=�lS��ɨ����f�@�E�c���Õ���yD���Ku�l�Ov��AH�j޿��vD�W.�I0�ޢ�к��/����J�@m�g�W��`�º��ڗ!�i���h����BR��m��£r��C��ɹ�+�m��Uh�w8Ɋ.F'7db��ZK1
`9���D.Q�J3 ���9�N<U� o��r��=�Q��F�#��ų�3����9���e�!�7�SxS���!x��+��5�P-5����i@b[Q��vJR�*�a	P>ڎ�C|s**)x���0��
���*�[J��`�R��,��L�$��&���Hq�&OE ��9��kW!�u����{f��r7,������Q�3��s�r8���l�rt����mt�S~�� ��#6�?M��"�b��i��QM�M듿�o�w�@[!vs��J� ��6�:�i?$u:ib�wA�T�{�� b(�xõ�1�{�B�?����JW*���H�r��_m ��r�F�4��z�3⚜:���>���/�� tM��53��ぉ{�x`ox.�m�-dy��v-��t��? >M�q�������?����8�]���� �>J�'�294���K�?����g=_���7c�W��Xs<�Dgr�~�\���A-����zuL�tǳ]t(�� �P/�a����\z�}�*��|��7*�AH��%v�	�7�-����j�`�[�%}T�f����\��kF!D��t�9w���{���Hx��)���c�޵�WWo��I�����f"��ڶ R�d����,su��\�b�;��,�$3���8�����Bcw�C�;�3h��l�'P��.D�^<�Hu�J�>L�X#�9��������m���/jm��H�yk7 �uu��|��Lt���R��e�]��d�H��2����'o2+!_�آ���F_Aƚ;�P�C3���i���Ć�l��Jmli!w~G �K��tDN+ټ����p���ÃR#Բ�m�i/N�~����c{� �<!�>�TF[')q��*�ǛJ�I��y[�}9!��B4�x?��ItO⪋s��1qa�s�*�߮���ᮠ�P*�\O�h�`��'������ ��hY�@�<���i�I���S揼�=c8����W��:N��7A[�sk9����P�I����G�♨98�πB�j#��f���4�W�7;U<2�q8c�ץ�;;�����V��M�۠Q[�P:,De�%,Qk���H��-�0��Oo�D�8n5zx��e<����~__�M�ˎ���ͪ�LX�+���6 zp��g��t*�D�6GG��'޽�iL�@�P���VH�6����U�g�Nw �s L�"n���9��w�*5��I�U�����y��x9!����w��-���@�?�CVm6��0q�8I���ڦ�Qsθ2q$�3��fu�Z��Ao�gߒ����z���=��u�����.{���9H�c��@�XhE�d� �X}�(�ǧ�vyy�pf��!��B\mf��8r�X
h�%o*�ƜH;�nCx�#З^b�F`�moi��4v��7�l��I�؈�ӂ�i],(�e>L�����Wz�J��jw�%�^�v�W]pɧ\+���w��\�)�7��i�F�41���ď4�W;}�]+1�+L�k&j� �����;M3_�q}n(!~�����˧J�8b~�#D�uؤ�1��D<�S��T-�lJ�<;���=d�7z��ıe(5���P�4�kږxjk+q8��b�'	a�t�]<Ұ=�n[��nf�@��T���� ������ s����J����.�/,�%'�u)��4�DQvS5y���������R��Ռ&�Q���d�3dg{@�²�pq^��0����C4������ռ������j�B	�DE��Vn�_�A5�8�da[|�D�Z�n/e��7����S�r���������g|';�gS�_�\���M<Z�����?o)�e��H�mG�����j���-Uӄ�*y���I�S�X�j����C_�ՙ��^]�i�#r���j|~��	��F�<���Q�-%��\m�_�,ĭ��%��*����9��в�?��``�M�s�cq�M�Gꢽt�^_���{�׼�4�V�NH#���PGT�-���iw�L��+���=:X1b�L�����/͍�A`�F�H~�3WW"�9��E��_՟0r�{AA����tR϶ڵ�%�b ov	�7���%d�IL�ͯ�jC�~s�&��2u`[�����G��}�����)A����d��9(z�}��������H"9�<�%�2R����,r��
h���A����x͸�MXT�[L-�J^��g�<!��T3���W~|��F��<���>/݅��h�U�f1����hW���n�M ��}k:a~�$�V�sP���	y����L��DQ�ڣ�L��g?�9������w!�HE����+�<�f��Ђ|۽����p[ƀ�u,�#��J�Xp��M��m�'��y��b��1Yx7zɎ���"f!
{:�T�Y��)X�6g
��4�4�C��k�����!0�e�0�����@0��} ��R�`�mKzu�*��j�E5��
a�����t{�<���f<J��|#ڙ�{������+A�?y}�@P,���X�>�>$��;Ze��܏=!ѥ�䣃�^-��p՚�k��Y���EM����f�-cq�
�󌌇�?���Xy�-�ͱ���+�BP����#���|����6i��-r��L
�>����4��g�`��׍�yA[`�R���j���M9�0'�|u�c�GXkR�K�{��=��y�����^9~b"�h�e�����B'��\�/g���EB�;����.�`(�m{���J��ι~�96B3cʎG�v�etdRk�+�����A� �'��m�Dpy�'��1�1s��L-i!r\6Y����E�Y�_����a���_����;V�Y'����֊��(t�m�P"~Ք���?�nL���=��w�O3��S��-$'���άg%�p�\p���xQ�,����������J�{��o��v�zk�#@sl�u%�1��_2}�CɞW��޽�3�R�~M���@��þ#�`�? a�ƤP����B�p��B�����L��Pa0�ǳ�3�9�3�� }]k����˥Z>�ξ���AX�=�e�4�[_�E :��4���k��!���6Xz*ڸD���b2H�Qj}�r*�ic"������{���;� �ҿ�K2� �->G`NR]fIR|T�C�\����uQ`(S[Y!}gKڸ�A�m	��÷�'(O��&eZ��]);|Ŕ��%�A2[�F���eʈ(nB#pf�o|VT;Wz�1��6���j�Z&qu�&���B�Zr1s�l���c�=0a-e[�������Ե��%W�����)?�e�5�@��D�Ǳ�u3Ǜ��^�h
�rE����e���m�m�M\�����o�tv߆ݤBQ/��2���h?W��Ee ˬdi��}����M���?s3��t�5d�e�p�i�q���ss�����V��y^�Մ���(����*b)�=S������/CN�Nj(��%�����}�*s�v�	M�Q�b��j �������Np��g�N�;:m�=K�̺��}.�̯߽x3�("G�|��	Ոā�.�b�x�N�b�Nm#[Ng�}ec��A.^qm8ܶ�8?��y��G�'���Ҵ�3#��g�ez�!���v� q~�/a����#�U�m�#���c�cʍ����|IKT>'j�a�������Q��]}��"�wy���6��ǔs.'@u��a�2.�y�˖Y�6���G� (�D����I)���U�d�*(r��
BΕ��gI*5f@B H�v�fզ�7�Ǌ�?*�J�󮬼/,��mg��'�����;8�/�Ɂ�c��N'9u���X03%��`a�H̷d����T��bP��"�Qro���Z�]�:�� P4Q�Z�|l.�>�+�{^�̜���+Sx@<4ȷ$�j�;q�If�ez�CIx��uhƎF����S�ctL�O�ӚQ��o�/*3�����R�G`������Mv2�A�2��K>	8�Z��bI�-�bN�N7e�Ŋ[?
�y$Q�<
�L^u\����om��UׄפVO+��f�Po^�8]�޺�y��-js�x�ow�$$],����kZ��;tl`��w��:^��@� ��k삝��c� KӠ���<��]c[�k��^����o���х��p[��vf�3U{JQ��a�Է�n��6/���e��\D�c�m��s�r�(nB6��a�j��Ҟߏ��Ԕht�Ҝ�X�-��j̓ 0�����nA�,�r��U���d�7ǹ�N�I��1�=}��D��D���"c�J�`.���?u�Ïc��'��o��s韨W�\�L�W)���SmiQƉP���P��;�0`B�����Y�!�4-W��kic�=3R�
v���Y����8�'9r���9I��v��>�Z�jQ��P��|Y�ݎ��P������� �l;�i<�×؇BKt5�C��V��)=<���Nɥ�ח;���p���2s�������u��=6�+��xAGJ����A�A�	oAa��-|��$�w�sub��o\f��M�M��6��R��1e.kơ�W���ѽ�-��$�ZB�C�3uثӧ?�!e!S��VgE��;$�i�vUO������o��\�.� 9`
�"��ׄ�^ߨY��^Z�iv�.ޫH27�Lp��f�����y�:k����D��"����>k��[H�U�?��kч�}�#�̃��FF��k�"��A�V�M�b^2����9G��h������'��b����h��O��n��Q����X$�AWD�jb�-�����[A����M��	f�g��(4{�͍����-��󫨐�i/��L#<#䐉&�G�a�3��X���*{n�T�b��/@͙pUI?)\G�rq��G��:�~�'W��38��ɲ�Q��h4�` ���dv�k_�U�3u�"���65q��2 Њ���M2t������Qs����:ۖG�<�T��:��1���lf�J�+Py#N�i��cNQ�g�D��y��]O�5����[ذ��$M�]t�2�m 5����E�t��{}<�g�(���'��1��y��i�-y���FCZA�~�ߒh �
��͌�<-g��E�� ���������tf~�Q��j�8��ۀ�Y�%�o�%(�Q������a��z�+7�D=��]��z�k�w4-�/�:�b��[���������;�!��?|�{�$�aI�.T4���Iz
B��=��J��\��"f�3��6�v.�ޡy����\�v6���!�A�����S��8 � Z����_:��V��Eya�]�R��g���^3�_	��o�^X\]r����6]>g�a<4?��r�zG�>����낏��dh�s ���w�i
�>:�A���Q
���VWRC���Z��΁X��tt�]{���󳗕*�ץ8�&��&�u<u��6��rSp��6<tO�M
R8�3	���Z}�F!j�^����;��
�|i~^�ه�+��������N��e"�}zW�d����2�61q6,T?�+T�֍��"9�ϝݼ)F��#	�*C}�5
�u��ꍚpTq�DS�[� Kxz���NX��A!��
~_��Z�[���_�V�N}W<�cOuI�Dڂ��*���َj��$b�TBU���1�`��f�k�l2S��U�"���@dL��*�����c�a=���<�p۹���4�����\�� M�����[��|�Ρ!���a�������E�����sq�/X������{Hn��)f2�$�'����9��a�/q��A���Ngm�X��|�ۯ2��Y�����3��3M¹3�r�c����uѳ�>��SQ�_��5`ow����f���;�Š�8F��K:�q��`!��F�:����!���FG��#��s���;��O��pb^����{�Ѹܝg��B��f�P��a{�|�/C!� :�-s���Y�� ����T��s����A˾L�{^�i�G��1J��R�fl珧�fAq��
�]Y�na'�u�co�jW�'!��՚=3)w�a�R�ć�Y�B	�/��?-�l&�6G���e����`Z\��ʪjLu���9����0��a����(�;K�s���HʁB�*S��Jk��jc��5�V��{��dN��IE��c��Mn��Z����g�Z��S6|��g����*'��
���9Î�?�.[´^�'/+Ə�TX���K> ����6���L�9�aj����I�t|A��,Z��B��F�z�W7������,
��1%��v=#?�"D���e	�Ĥ\�zjL�R$l�
�̦�k����+.��ǯ�����6�W�eeJa�h��:�ԭ���"窢ڹO%љ�ORb~t3ݰS�.n8�G�d�J���ڪ�kJ���4�>W�	Q�Q��E��?��A]h\�����/�ft�����+i-��oaK^���D��7"[��ˋK�*�ֻSJ#�7�Km�9��+�籨�ʆႺ&��X$��uЫ�$o���m�)�?��?ί���Rvp\V"U�
��w���-њ�IP��}Ȱ#���q���B�&6��襕@:'�����?r5G��g^��-�z���?����qS�w3�����[D��{��,�V�v��]����8bf��$�!�}�-YӸڛIj�خ����46��rՃ2��}��ɰ������.0LTE� 06>v&�JzY�h��7Gu27�ld�)��Y\��3��Cܰ�f5�.㻷$l��;Px��b|�"��\h�_�Y�������[�`���+� ݘ<�G�/P�/�����Jʷ��6�h��@��Ý����.���|����y���(�c�ɮ�;� ݪ���/c��m����ºwMB#Ӌ
�Vz���;P��)H�2��>�W���^e��?���G�g+�:â7Nfl�(�������gf��xy�W@�LG��n�y.���\j�v�����;`�T����AQ(��⹰�s�W9v.�����l��F�_�N�R�ʭn�7�
���3��5?���0ٵQR,��@2�{�dP ��xl��3��>W�
W�N*�NP�{��o�1��Ȟ���$�+���9��Hw�[3Jk���FS��=���Q�
! �K?e���d�m[2���xy�_;�[�zV�Ո��pڥ�Wm�����R�
�cJ�4�^P�O�(�T�#Z�>��K�!ߐ\栿�c����@r�����UL�X����3%$��'Ճ�3f��c�!�3ܢ(V3wH�A�ۺh����.!춗��)c� Ng���=<4�!�ANv
)TB��F��4~b--H��j�1޼��.��N%�H��]����W����I�	q��i�b�[aD�t�Ɔ=ؽ�?5ʥ����b�bx�W�R���x�j����}���T!�-���)%4�;����,�	ɐ)�����YJ�{�ϑs�LlD4�܆��Ye_�=�����fϐQ7��z��8��R�p )3���3���Qpq�3\��C��_o�O5+����jI�4����Ԅ<��qgM�9�*��0]?�=�r�`������,�7ɒCW_�L'°�� ��C�y׊K�_V#w���_�N�Rw�C�)It�����5���S�j�ɗ�܌��Ah�0�YČ�z����(��lO��9�����ncL;g��_�b�������q����B�)�0z4Ĳ�!�Pϖ�ny�����9;^K���t��3!}�Nu�k����yi�c��/kf)`����pFP��-"�L<ʫυҥzM �[?;Ϩ� OE\n����LY�s���DY�5�Gn�FQ� J'( W�&(je��D�n�7!Tg�g�Z�m�e��\�WUGK�Rn[��Z#��<�QZp�R��$m�$�qQ�H�3��;]i)6T���.�8ʪXά_��֐{h��%p��w'I�Ç�ODZet�O�Q�������i#(6�*�����Ym'%.�D��Yp��zjYe<MV��ӗ��H�R$���L
��h�r��b:�����	�8�d)�By�%π8�)��X��X�UP��x,bj�/$K�p;�să��P�߿>G����f�~(��w\�Nk��X�e̶�����ζU|��g��9�HD��!��(��(�+΁�b���&:x)�Z����_�+��y-BZ�d�6�Y!�
�F
�e!�u�0�,5�gi)o��)��0�Bݩ���2�,�8�ElFOҞ�gQh���Y2�I���]�+�Etta��g��X8����R�T���Y�p�����;H�8��c���9݀[�fl'A@�lt�ף���A�t_�[�^�4[ Lp�L�pKg����^RG���%=��yO�J��	�"��uV2�'l�4'�Qe�����9��*�|�x)�wd|����K�ۓ��0[o�:���~p�o�*C����i���&Hn��M�;��`y���%cZ�+�Ti�Ѓ��X�3yyN����墳˄�����s��^����sD���5 �Z��p�
�EPk<@_���޴x�����k�$��%�X���Ra�|M>�Y�{m�����в��O��[��Y;�a1-�"��8�F��]�f�� �H�Yk��k��T�>u�h)S����Ţ椵*�1��+�X���p�^��+�v`HX'�i�O��5&�&�ɀ:�y��g�k���Uk�U ��E�.�d-.j�3-�ֺ�k=&���ř4(�L�| ���{U��� MG����U�{ۅ�1�o��8%]$��o]��P\�$��D����+g�h���e ��1J�a)���R;�\7�?|i����VIq[���es�:mf��:�2��觪�PAON;.���]ؘ&)�a]��؆�r��"��إ����!���Z=`HN����}ŝ%�|�ݷ�Oo�LF��9u�F���e�DN`YSCƪ��ӆu��-R<q�0
��� ���V�u���ڥZ�QYמ	���Ln�8�.�O����l�R	��Q������	�A���#�/B�j6V�>�-�:>��94;{�.O�h�BzTϫ�=��@9 *I�lx�}�o�M�Љ��텘ŵ͢�
?��fӖ$m�鵲�k�1��F�s���t��(������Y���R�MS@-j�tl�R���g�*���'�(�:y��$E�.7����~��^��c�z��Y%�m9]?���ΠיSD��9��M�	S|���U�7)v�)������$?T��Ŋ�=�o��g�O��us���^>�[��hF�:8.����y���pd�u�^\Ppr��#��M���Jg2���(�����K���ҩZr-���U�(QƞJ@�𛁷f��T�aj� �{�:���ۙ�}o�cmz������$��j4�+�%�rma�����`�nv�,����M�����Ad��b������Ԋ��Mޝ��\U�|F;�%��_xn��H�p�F���;����o|I��b�Q:(Mh��POÐ�'pӓ0���y���/���[��B��81j#+��;_Y�]|���c5����8]����v���=]x�*OsĬ�DV�M�̼e��x��!��f9��W}f���'�A�}�j߰�����e"�V��K��&���o��=���_%����S��VA�&�1n�	��w�jr��Rj�f�3u���NX���M�y&�	,CJ��J2D`p��e����K���z�_�aTC��dMu�F�P��J���.�$tD�3섈���������ݧW}l��
�X���ڴ� "��i���4�}\���3��� $��L�&U*�	���A�W=p���^��]7r^?Ԥ�g0���=`~m	��^��S�g��
B��fZ=x�ȗpa�R���ٔ�c�,!�pt<s��}o�M�I-D�R?�Q�7��������y�v2r"96�ٻ�+s	�滴����H>,����qid�\;ql^H�Y#N"l)�Ix(��M�9�wɩ�y�����3��P2%(uڞޛn�WQDlpq-3�L�q:�Yn��I�q�zG�pM���9K�5��֠���Q~%��"�Ѵ:�������p��G��,Ӷ1�N��ߓi�/��
k��Q���j�(���s��
��f&`F$�+�2�z��Z���V�����~i���O�7��z� ���#�%�޳����������&��� Wjy۵���%"gc�� FZW}Y���fuo��"]��Y�4!eBM�f��[{Sn��Q�lSX�?��`��̩^�9-_��B������v���'L�����u�&:_��,�X�6p;dS<-��"����s�ˈΩ��$腪y��V<;{ ��Č���M�x!:��#;�Z"��!��HU�ZG"�6�?n��_�2�d�%O�5S!X\,��w,<x���ms��`SڲG2m�ޭ�&��*8XS��H��X�,R_87L�L�n�v��[77QOǻ^v'�g��m�.��SF
����V���;yz���x�$��[K�����_�3���z[�׹��Jx�|QE0�Sן�z�Pwq��߆�0�8W�hL^��� <�TB��3�V2�\��~��VD�`wȨ��u'c��,�)��D���K���O>K�l\�ˤA��{� O,nY�)�����(>^�������Aq��2oCu9�U24�S���T�� ���@�5��uG��d��.�AF��/���ۡ�ۧ�P�D�D��_%5<�ҍ5�1�x�H��NqXD�e� J`��N��7n���ۅ�����g��~D�Z3k���� b|>n,c��U�t��3��{Y�2U��=E��7�����Yŕ#����іL3�a�_!����YEG45�ƕ��d�T�}���`�w�wX(�ۛ�q!5�M%�<A��_�u�fg_,��Ae�*;�?�̎(��Man@P6c(G��Y�;��8��v��o����:�����!��Lq�#��yY�<�@o����C00\��Kw|\�O��e��2�!��O_2��(h
8��A�5@�'�f����7���x����ke?k�vԶ��1��\ʦ\�p��sE�[��{սtE6�o��+�ߐ���7��s���&�a��~�k���0:��K���h�f=��d��D�w>�[Y�����w�(]y�������gC�J?q��.[���z��B�I�ֲ�L]��v�Ӻ�B�hG��/��%�7���7��)4�>h���oV�G��v��{�-(�F�^��I�	͍2��{�'I1
1C?���~��7h���
�"����x��2͵ci�cZ:�]N��X�@mk��@�Sheh+�2N-�8��`�|<��� fj��� ��Wq��>;��ӝ= >���iV���l��%���;���,�H�R���s��i縈&�vX�ئ��c�'��`4���"��T������t=��-ɖ�t���|�M�!�z�g[Hr��N����r숥`��3��O~�`�\��bc��pv[�1��-��.�_�˶�D�G�_)MPfI�p��Y�GO�:���=6�)7�U��Zò@U1~����Yե�lK9�C�7mK_1[�
k��w ��Li���0K��.��.� ՠdRp��U�󪎩'��A����&l_X�JI�ڭ��TP<�/��-=j łvytPQ�TrJ��s��T���>vj��S
��ӕ8�?x��,�3#���[����dԂ���,���8� �u�:�����kh��ϻ�����i�ta�T�c^��m@96���U|i6{�Fdx^n��6���!4"��=pd�kR����g���6
w�ZR[�tY:�$-����6��:k�3����f�i>�������|B���2V�ͳ�r3ׁ��>�Hj`��Pf��̼����.}�0��Q~W܌_ו���gѳ������D�����Z���[���!��d�N��Wu�&댆�S���!L���򅖮��-+~;f֞V��M�1p_O��y[OJ!(Җ+��Ri�a
��[��0�7!%ZQưF��Y��wd7���[3�S��iSM��.�.�sh(��Q@͐-HO�;�*��y$��P��t1� M�<͜	�-j�G�Ә�]#)��|��F�p��#�4ņe;�N)A�҇�Wz��;(�d��y�Z��;	�\ѹ�C	�h��d\�D����J����q]�4Y	�)�زb�}�u�#�^��'�������<�9����J���R�މ=�����3<���D��<� �'Jo���N0�����ҶV����РD���i�GL�346ц���9�BZo��꓉H_��I���-�����H�$J��Rx��X@��<�a!5F��Z}�F���v;2U.�4��7����HI�t��l�w���Q0s�ط���=i��W<Xv��'HF v|PJc�Ł>�-�]P��k�O}׀�KQ�mM�uv�����Ր��k�QG��R��~�<u�E6��3��u�vvi���|l�����#C�B,��xIYn~Kl�{$�x��ٽ��W�f_݀�us�..\�X*(�bԷy��裝)Y�nqL��o/�1?V��+~D�����s~����i�.CN�B�����j�>����2d�Ss8gecyy`�#�T�0V������eFD׃���
�࿛�Q�f������F�21��vѐ��[|�v�x}�:�����A��j>7�:��ܱ�tB�]{�E&���d��,�;�֔��^��i���@�eѹ���d�h���kJ��*5!��g!����i �A��� 2o/�^�Hl�T��j�:��E�(���6K$����� r	'f�O�l�{+*�W>��h��|^�o�t���`��h�~�ӂ��������1��r��=���k�7�`�vEI����o���v
��練=ګ��:�m\i�����exO�D*
�<Fd~� s���~�t�'�Ԋ�]����9�_������jU-�qK���z�9�,��?O�G�Ic��̔�U�^�k�m^�>��E�Z�m��6�u��{��"n��_�b= ~Ш���h��60�{e���l,.���c�'�g�ywIi��=r��-�p�B�9�9�J/ �1��)YѲhI=8�0Z���am�,����9�j�ď�����	�R��K����%���,�PAظ �@�<n��5�ϵ��|�ο=�'ż���k_��g��ƍ�u�A�P�	�6�瀔<v�wzs-:���-���] vP�#i��W��x�Jj��o�k�GY�ހ�xD���d� 8�'�{O2�q�Cam�f�h,�&�-�KV���IÇ����W.&�S�M�3�ք���;�3y��/g��f��c,��
��m�#��_B��2�ǹ�>�,��G&�G˾-+��+�B(aԓ$w�SsJ��K�´m|�%	kv�����%9Y�yla��_�q�&2� r4p���d�v���j��Ň��iNˣƚ?�ig��0��6���5+M�q<��2HB�zU��ԉg(��Aj�����'���i{.O%>fש-˫W����j��	==prMmUU��6����ı*#�~���+M�v�2i���*�87xE�PQ�fC�����S�pӢ�z=�Q�9C�ge[���qe�Tj������g����i��Y���[&��Dm�r�/�ftD�5ڽÓ��FP!jzL�<B��=�[�0���!7'�u��Ÿ���W��]�]X�Q˪I �!�+���'#Hކ�ݛ��G,�|����g�8y�7�5Un�5&6�8��(	��	��d��M�T���'�0'��x�%�[��V�_r{ Dj�s#ۅOz!���~�a�1��h�,к=��l��E	���Q���٨��	i��4���%Rn�W´��4�/Ɣ�)��J\mq?XU?����P���.;'N�5S�y�Kl���<�#�e�EUR?3�
�t�"�V��8�t>�a��5�
��1Yx~����u�!}mQ���2���!��V�byt;d��ʀ^�����R�c�T���WΈ���8��)����3����:����m\^M�����^WjeHOB��6W��!�$UxC�]�mBtw�ѦPC[����e�XK�d�W+Mh����� ����ԏ_z�3�nr�u�� Ir�������#������b2q9s�R���(cd��B��3�&\{|44���|����o�-���_��i]i1��	��ŠF�	��[x^.�H��	�|�Iѯw�������z���yU��=+FeCiU���'��(��Gh_����:��^'"�(�B�u�Q{"F��ft9&��_�#�چVӏn\�ʡ�Dj���?�Jj��2�+�7��8ր2��D'����j�et�����'��07i-w�чG��a�`� S��	�����MZ�N��6���v��/v�?��&�/����.�ܤ�� D��ԃֶ,�������j��g��r��Tr�~�]���3�m��~�mi�tm���L�X��}GM�]��Q�ыH�ʕ\�|�%��"À�0y���,�w��:O,Ԙ#��x}������WG*�Mm�
��B���4��u@�/�E�چ��b�o�RO+�V^�kez�G�&�Nql���M�Tn��[�A��}����Ŭ�m)y���{�߳�I���"7��4'���=Xoh��h� Pc�i)�	�=U4F �-�`����=B��P�,j)һr�G_��"Jb�L.vxCp��xm�R���Dl�:0�B�����A�_���xԢ�ZE߬�#�³<�Sw��ag������߽����*O��X��N4'�ۣ"�=b|i4m紛n�d'�)/�/d/��$M����׼5?(,5�),}:��L�-���r���~��8��@�W��
��w��e=�� Q�C��M�r�6��ce�L�٘�	+9�԰V�}�m[��*f8���x�ޟ`��k�UZ}Qn2w���xz�7���q� �=��Y�O.�b?^�<.�3^���������&U���<�7��t�1/Z�P�riF��6q�mf �N��f�i�,�Ý�r���6��AKm�|N�w��f.�ڍ���H)���#
'[��fL�H��IX��y^�w�b��Y�Q���m�� E�y��.����	e�;ϛ+:%hl�^}uj��]�~�j)#q�8�V!���I�͆=�A�ָ��v�>��@/�<E�����~훿��F��9_�����(��َ�
_G �������*�@4�!��F� tg�_��[�t^�$���J�E��fF���l׈���d�uCQ����Ϟ/�d����R ��&2��W��w��Vt�hL��D�m��h�~b=�_N�{�+}�U��]�����'�R�@�ޞQ���eB���>��	����ϱ�aK��ED�7A:�1ڷ��&btA<g��퍷�\P����۔����S%� <��fy��3��D�F.8_d@tڐ5�eS�_�Pr��gh�l81� ��_o��|c������h�HV�a�;@OV�s��`��q�|A�|W�7��[��H�-Q�ИopJ�����ϼ-��*��OQ� �|d�So/@e�n-�k�6U�ř<���
�{��NT$���#%:�ٝ�d,l�(p���,C~cC"���s������f8WV"���� �dʸQb`����< C�1�>���X�'�$������X�q�J�2U?��CvJp��2�C�lZ��,����Mm�a�3 ��V���O4a��j��9G8����c"X3 �/�?%�V��HtQ��8�gs�ӈ�W����B���v����Ǵ�5l4�::F,q���ʥ1�m��!צ�x}��mu�%0G*��V�Z�}�T��;�	��E���g-��4�;�*w��X�9�)c�<�a���qy����ɥ���\A��6`%+�/�WO��W����U�2�$RH��2*��V�VǄ�Ϝ�w^����U��B*����l�Y}�p�����)l�޸�����:�j,ω�!T���;���.�լ��AV�췄���b�0L�8:���sL���Y�@_*��mU#o��Gܰ�p�����4�V��
t];���;�����������ŷׇ,��ΚhO�������� �N�G�OYbN7g��
M���v��Pp��<��5k�t
M�pe6ѫ�(�p%���MFe�w��J�&�����=�\�d�9]9�0<�p�C�Ɣ{�Ӧ{�OФ	Z	ʍ�^��
��S�K%���Nm�L#
	��8��BQ:
ߊ���	мl�Ū�	�֐m}$�5����J�9�9![vTB���t��5j@�����C	�����jՋ��� x!{Gc	���]s�4�g͞��5��t0�6&�Ra���GӰ�V��_�����ep���<��N��<&z��+�y��h���ZRC�I'��T���0�2_6/ʗ��@1ڛ��}����Yjm�F�c$܈yA-�%0��W�8c�-�ޟv��y^�űά�%�&\�ϥW�܉��E,��8��T)�����)C0~ǲ���Ș�yAm���Ϊ�v d\��i�vB(e�.��ހT��Ʊ�CD0V�{.r��5��#Z�0j*Ǒ�O&aۜ�K���i�	�H�tk-Tv��z�==��C�Q���8�ީ~�hdL��y�֜b%i|Y=��u~׎��W�o�����5[2��&���Vk��k��P�$�q�]�/::�pw�H�G{�T�l#XUh����p���I�?��vvV���ׁ��~��6d�mC����nբ�_ʌW��Q�2_�a���M������/��	j/mj�f%z�4l�d20�OgW$e���zi/
Z)&Q���O�1�Vr;Y4��Ƥ\�Ol�� �ϰ����X�3نM�����Q����'�v��62J��Wv�J��{r����[͆d�QS`�U1���ψF�Tpj>�P� �td����F�/)������+���X�/���Ω������<�g���wT~B�V���9s9jڄ/�KE���h�96�?W�\��i���5���Y̏�&�+w�`l��\���E�Ϭ��EZ����F��Y!z;�joxW`ϑ��5��l�Qk:���X�xh�:�����*����U�;�,����ET��j?#Ȱ>����C�,3�Ċ����W�g��f�h5m����$z���\��Є���^SU��(Ab
��œk|��,^\u����>���=�w��n%P�����5*�/|L<R��TL$~I���֠�b�z���|RI
�~Y,�/栢*�L���n���0�z:B^��#��c4�����@4b�K�W�_����ߔ�dӸ�Z�=��c�Ӿ)s?�8i���N�'����x��*��6��W<E�v[�/G�ʵ�Js�����l�-��iT D��ݮ�=8��A��r`PZ�q�Q�:+�����sr��MR2���[M~�h���P1�����4�iR���܋�m�s�D��>q7o�zk	�ѽ�vXx���}2��Is�Oˈ}�p�H�bAh��u\T*ʪh_���_�@�����]��[�$�("u��Sp����MÙ}��ts����>IR��B��"<�JF�{�$����e�B}��-�����q�zs��8�7�</S�**9կ�t�v���ΖT��u������� ]�A.a:��]���aΓ ���J_x6� ���і�#��Y�@�mW����m��[�5%hT�2�sa͖��c~I:��69�'@]F���oۖ�4��}-�p7?k��C+���I/[�=����O����M��%�洳���ʸ����躗u �׫a���m�U��<�Mf����-�&�[���q�5�$�:ʵ?��]1����w8��V��0f>��K�?��H�8�bt�F��c�k�����8��%���J���]0oUC��7�d�H�W��I�����&w����y�a��'l2F��/Ƭ�s�e�� Ө�.*8��4z;�g�aH��L�:9׻��2�bu�	�Sx��zY�n��]�*�9��Sh���%�&��bAfأ�ՁC�J��e���K����K�L�g11h2Q���|́�ؙ���r��:�%�@s��9�e~3Ź�4L�$�E��P5�� Rf��K����􍟺�?��P�}A�O�=|;��-�Hn�r������~�V�>���'IUd^-��{"�k�'�����_�;NJ���_��@������hi�菎B�~_��F2nֳ���ұ.����l%�hċ ȃ�=kې��x�����{����rd�Y��[�󺤹EU�g9�-�?^~辮�!+��d��_����`.(7E�D]� ��$_;c��=�ڭ�}������#��(r	Uk@����(��4�
jÚN��9���A�c��/v��C$ܟ�M��#����������	s��AW�>�������t��/����y�p(s[�q���e�N���Q��W�4�Bo����*^bq�����p*(�3��_�c�̷���>�.�m��c���[�G�8rh�%bZ:����xX�z��X�V��!s�DZȌ>y��"%��oT.[�2n��&ΙYk���%:���W`4_LY�;8�;�WER<Uˢ%` gG�!8>��U�3�O�\|6�U),o�v���k�"����Ěv��ـ^t���#`eU_ T:��Wf�r�Rv94�4�@V*EE=�c�6��(T�<Zg|d��I�m�\!<���j*up��񸚋\O�"�K�A0���d#â��O�Z[�C��õ�#�ԍv��Ϳ�%������V�yn �:&����b �<�|( ���� �޶��������WMW[��8!4����l��Rh�ȈD�RPvV����$��{k!Ls�3����ſ��#0 �:	.��uoEy�����Z�}�z+tB|SH�i�Nx������DT�JL�DX\w�dbyc�f~����r<�Zo��6ȑ�ҁ�-�_�}�\G�oh7�hߓxT� 
xz��I��KG��S� �r��0yS���;�!�#��j!`����β��"ާ�
Qcu|y"�[EA��d[v���ho-�%��І� W�,b�e;�%p�LeW�Zx$�u��2��u�S����5��f�#��zċ唇����ǋ�t�fr��9�z�·hy���kq<���1�J���"w8�Y�&�r�Se��=2��X�F�,�fG�$�si�텴��{V�3�11mӽ�s��
WG �0:"�˛x���I��K�'��<K�'��ϓp�" M��Y]�HsAo�3�u�k�=��z�7�5Ǩ¨�4.9�H>ň,�g�!
����˒����~�i0�Z�,ᠼ�"3�f�|���&������t4
[�l��������5A��)k8V�*�{�}Ey�{gw��v>'��^�+�NɤhOi�������H�='{��w�����WT�M���%�e�e���yd98�
��W8a �jTV�H���l��^�����A�x3����q��+��I��g��w�o�,݌��}�FˬLL�W�X��0��|͵�Y��k��At^2�~��(�ʔ�6���҃��|*��#��Ra��t�����u�S�ߛ݁���a<I��(��	�C��y��T���FӾ���p�!m*��Z]�x߳<�{��v�7P�����#���{Z&"[c�P���L%��΍쾧��瘷d��?0T���f8���q����#d���L0?���?8�?*��n���1)b�7֨G��ekn/��^o��c?���O<��+��ҧ�6Ϡ�h�� �ۢ)��@J����"�nlL�:C �/����ظ=�˝ҿ���#���*_S�w_�|��1���-;֪�]�U����ڷ�p��y�D�DYm "�D��U�'E�NS,�-i�Irڱ��j���#:�Ƃ8���<MW2���"�ֵ&�0�e�J,<R;���	o�d?$�D�H�k`B��Ja��_���ʲ�ؠ�	��)5�Ո��!�����M𲊬��[0��U��C����OŐ?F<4r��za���*�/t(�2���<�R�.���[��j��$^[�t��}��gt�z�Ǵ�Mre�TV�0,yU�QLi��OI���N��F\x��O� :���1F����������0Yئ�T�[[�v
�<q*�P��~��il`eR>�̟����l��-��m������ܢ_�JV�<v�s��d��3��V�4z������z����s�XS�S�8�a�������9}ǒJ	�o��Wq	�2Q��U*j*������힐<#���1�!q�����;�=S����UdA��#6����
a�&�"�Yk�A��p�V��<p����˴��,`6$ڠIY���R�����^�s�[J���v�2�@b���o�ӈ��gK�(@��qyTJ�`����qf�S��S^Q��
k��4t�s��N�Y"�/9>l�%��4����&��H���}���oan!�h,]��v7��#|9]t�pc	���8+6��#��`�ö��ߔ�B�� #�Y���H�Ȭ�[��QE�6
���B
"l�+��r|"܆3��J!�C��rR����V�^���S���I��`��`,QH��],��B6���X�i��*to�:L"�ZK�뻅�{s���8��6s�S:}Ƀx��=!-8��
��!(y����U�g�	r_���V-d�o���+r@���P�Q���Ya9��!aZN��� �n�83r�����q�T%W�����-f���F��(N��I��4?cm��r\;�#L,+6�G�Ζ����W���]�zR��x{�x��hۢ�xs�L���=�C��@�����"C��yyeq)�,�bIk�@ i����#�w1��x��V��K|�(��7^w=��Fh�VA�}0@����h`�3k�Fh��27�6����L�`Ɠ����=F#��v��6=�i���U܌ZEy�l������ѦO�J~�@:s��	���9�\y����H�GĊ��?�y�r�'�#i�4xs���mF����J] �_�.o��ώ67A��2����dF�#/9�+gh�M@�j oЧNb�[1��[�06�EC��ȶ�ڨy�~�;�"rD�j��L�3#ji��4����]��_���Xe�0��˼�L,�\�H�m�q�I<,A��x�'^�t�?'>Z^�5]Bc^|"��2š8�t)=B'~�̲+{���&�i�(!�S�n�lYwl����g ���ҙ��.�^�R.������!R �ԅ�b��0��KX�� ��(7�V�ǠqT`����孧!߬M�I+�|T������(�x��KL����ϩ4ۑ�v�G�	I�%�6�A��%HX`���:)�|y��Q��FX��8����&�Q7���>��J��"�ͯ�����D� ��Њj�%Ɲ�F��~��fk���L��Dd��A~.�M+R�3M�Z�)!���~�oq&Zq�A�w9w�vVT�w�B&���sW��)��=gT�Zj�[�hҩӟP$�
�y����G���J�v��"��7sҤ�����\)N^�d0�V,��S�7�G�&�t�`�@yXu&Jn�(�э+�*�d�Y(�0R���aS<�wi������s"����ʄ?x@ф�s��Y���� }��G�7`Dƌ�lB�
i���)$c-8��O^�q���f�k�BH
,�5�H�q/ze�`�G�A�|�l��ݪ�uhj�G�~�|}r�Ε���^l3!���B�%�fۢ�}F���.J���s8i�Hbf��dڇ��D�����r?�qE|���E��T+.���eS�Ѭ!t ���q���2��d��xkx,�v�g]�>�\����֜�
'*:��������
�R��Ζ�+�z-ْ���������$���K��c�sv�'��S*lB�2R&�}�J��(蕥T�Νp��s��f�R1w(�cv꣹!�4��м�t�MUHek����G�8�7|cQ�����x�_�ں,R���ƻ�Q'���m�;RC�"ܿ��R�" e�'�Z���.V<������i�V��P*Nٸ�"~y׼|ՄwPK}6i��tko3���/��BIL=����T�Y*���^�o�v��?����W�a��ekf��FO3�?��XK�D�/�u.7��h����YZXk�|��Z��g��H}����3h������v�t�>BEwm|Pk��wA�F����W"�l�J�Q��j�;�qۋ�� @Yb%?rUS�o��.��:�)M�0o$0I�j��&�l�kP�O$ۈ)�"'W���.�1O�����̚;�#x��z�w�A����95�F!�Md�A����e��NO�I)>�����p�2|y�OBM?A��2���?����ߔ6�� {���O'Y�E!~c}0�IP��A�ϡ@���[\s�tV��OAW.�
�4�=�#m��1҅l��`���������չ��{A��'��޼>#~��^�fXD�68\I�������&!�_�-B��9aM����S%F����f^X�#;f��%=�����1�s�D�?��$ti�3��q�RW��m�a	8��5N!, ��!�v�h͠��=��-܄�WfviX��{�>n��/�͵�oc��7���.�'l���6~X�[)�����󷿫�礵L1d�Y���T���j��E�TJ��	���x��]��,���?�[�!3$X�?��J��T6����j�x��G`#Yr}~4R�^�~
��eE�ecI��X��5V���H�n��P�r�s>R��A�@����{�,�+���	�Y���F�N�Ҕ�Z�m�B���ef�"�c��Ҥ��^���'(P��J�	����I�������)���>[�E���t_�
jv:�8!ۗև��o�R%��_H�)�h������'[6�]����HZ�ğ��'x��9tvF$a���m�x�r���5^��I(Sr�A�V��K	�qX��:�Fl�ݿT�
3O�����='O��1�mKqf�U�!��ە�'��Z�r��X����mx�X���=�^�LWHz C��D��GO=�2IC�Κ	�O�$tq�y�����iHi1B��%�A������f@0�=�Ʋ�z_V��;z�ذן@n�Q!}����7 -�~�����+SD9�W�^�Q�(�����~,�����d��q�"�~U ���R��arR���O��!AK��址!��x��<,ҕU��v���1Kn6X3�Y��k`IHS��3g�r����Y��}_tVn���c]t!���1N0�ȶ��8��Зﾈ�K�n6SC��f'`x�bt�K��٘���0&W�,�n@+8]��?°I����@�[7�RWeB2C����4�=��/=@<+�BЪ�ǘ=������wt��(�h�m�	m�LX"����] b��w=�1V��	�����ڱ�����!�}��G$���H�l�rq3����7DA��p��hYh�38����l�y<Ԟ3f����S��6
��LR��:F��u�)�cY���K/R(,؍J�]D�"�&�r ��8���DH��v�i��y[�z^�ۀa�+�Gm��/<"�y.�W�{`w-ޠHC��h6K��TT��M�W��k��K�u>�B�D�^�
�s\���c|tz;�%B��T@��K��~c�]-]��6�4s�m[��>����z���~���:����Y�G�s�7I���dxGH.ӭD�2F%�d�����Fv	�zK��-��Tٽz��6� �m~J48Q«��y� �f�ӷ��QL#	*,�*����l2��4�i����\U����<�W�8#�6��n��	����*��[���5%!�3��2|�"�3�����n,�FY�>2}%����ӹ&AA_Tyx5�t-h>�b�s�W|�]Ң��S?�mR��$�>��]��W�����<go�ȯ�fn�>��x�g�䏀-N���$�v���Lyag�G��)����r�d{c߰�\�N�Y��cm�(7�����y�XNsK������i�'�T�#������J�\�A���=C�A\5^�EU��vʹ��� ~��8'�C8+|4~������C��w�t�۶��#�q��i*eS���[��'���#�Yj^�ϲ,����x�@�!�̉U\�9�tJ�}�VP�Fsj��yI���/�U ��2��h&w�z�Ъ/�%�cӆ�/�#�rȡ7�rB�C�M�YjO�/�`C}P>pr����ؓ9Ih����������f�>�=%`�d�0E����YN���ob�V�V�*Q:A��L;��߁%!3P`��_�ѭ�[�]�?�/�_�%o+-����V��i�ɚT�h�j���&:�b`�N����(?��`��H�w#�^��3� ȓ�il��K�����sQƺ�����;a��i[S3�2Q{	�� �ԗ�ݑXJ�޶�|��^(inV[8�޷:��W�'3'��A|���Z�H�� �5v9���a2�r%���3'q�ک3��\M��{< ��wJ���_"KǢ���^� �Y;;���2(��0�M��x��H�mO%���[$�ƍM΅���Y�Gu�_��q+�8IxJ�u�/�3�/d!�ֻ�z��Q\��*����BS�\�;}A�ZDw!u�g�����fyAF����H�fo����"9y�"��Ϗ���X�ԉ��
|!��f�����!2�V`Q��E���<Ӭ�=��/R�,�j>�����䖃�&�P��Cš���b�i�,ߋ�� xaP��9=2��<��$斅��(0GJ0j���3b:MgT����~���e��,�n�vS�%G �DDJN]
FX�$J��Y�?ؖ��nUr��~ j����@	��������4���sӟ�E����g��I������(ʍ�����"��;� /[�/��yu���'�N�oC��"��Q��h������Z@��=	]fO�l��A���ۓ,���H��.i��> �T�(Q����U/� G'Z\4Hs[g�7xtE)��x��5��iGӞuDqm���U�.o(�Jp������d���s��4��{�?zF�����X�Ym����1��p�XD�E`/�{Oj&*�LI񋡥l�:Vx��0[m�D/k&w� e�L��j�_��C�a�"���3��cC(PJ�Bw��zaݯ��Zv�b��xp���Л7NÛ/)Z�Zr�ذ�3u�^'Rw��`�P����m�b3�-ZUR����=Evk][ӂҚXK$��mrb� w�����[X����Ω���rg�~�0����~��*�b��tx���oe�0VL�D+����ٗ�!}�����N) ����q�[���Đy>���25{�e�B�QO���3yN�"2�d����;x�\0(�O�8_{���>�iǬג��jP�3+���0_��1��+�s�e�M;5>���u��*"аJ*��t���R��ӓ�aRS�[ej�T��D��ѯS޸a�k���m��!�=Z��x��Tu�?I��y�Xf$z�����K)b��'qC�D=#�z[��)/�rE�a֣q*��s4���'w�H����hP�7iũ�-��,9�������5��o����*���*��Y��ણ�
z��JeJN����K��/�Ҫ/��X� �兵�K�ml��WAM�i�:�YQ ��"T�Y��u�=����-%?Y�&�n`;3�އ�~�R���ڥ*���||'+�j��r_�|��#���g��ɚgYo�Q��\VA7��j5�[9���oY�w����h���sYjn�,���y�N�\9��P2>ܳ1ME!���6���f*QK�8�I[�ĥ��E'��TO�ŜF�fb=h�t �j{�ze�Ʋ���RU:�;�)�|�
ð�I��ф,b���I���I��6��\�z�2K���=����V���vxG�Mp�,���įJ���WIִKB�܌�tn|��2�1|Y\�|+w��=��QR晴�a*e\���vv��n9=�u�Ї���_�L���l�;҄�(x&0���|�-^��a�"и�]�#��]�S���㬲gd���\����s/�d�75C�7��D?�	n�+��&y1H�wޮP����#&Z��WQ� �9�Z��$ί����O8v/�xm�F%��[H�ꃰc���W�JNcT�4w��V�5��ڔРU�c��E"���/R�Ľ�N�%ۡ��ПM
�Y�������M���u=5�⋨Ρ�p�?T���mO���ʕ�{���XBV��j�g�Xk-�+s�A��<N$ ��S�w��L�?��QmL�l�;���N�=�'�����h��Cp>WgǢm���3�FΕ�\P��`��|bD{��FuJ��z��W��V`�٫��A�5��G����C�ř�a���U��������G��z�VWC�%�"������]�<t�%�&�!���;�k���Bϥ��o��_����\��Hʣy��y=�$Og��g�E� +ӗu]��Y��I��z��[/�N�Y��?x	�-\�c��ɏDP4��\��,zx�/"���"�~�����<�b�{�z\Yy

G
���a��ٿU�[˳2�yJ�n��'�%~Dm�%�J����^L@������a�&fU.�;�=��BƝ��Dp��#XAe��ۗض����µF,f�&�?���Qz�t��A9Z�E��\*�XtL^@��FG�:>c�0���5��J����s��aw���^\b޻U��b�a���(��@�N�tB��пu��1ݸ4���T-A����S?g��ð�-!��"i2::�A���f��oh�ÕJ`B�Qyp�Qy����
͂�wwo����>}�L�P�����}���u���ؙ
m��#��q��v�F�tۂ��x��z�A\0S�����(x��C M����f3�'��ə���[�4$���P�	��?�O�sn����$sp��eZ�$l���O߁`�h
�.��v�4�9�CC:p���y�C��@f,�tЭ��\���z8S����:ܦx��i�|�_��x����*��べ~F��⊔��D/���B��%;�;S�a�������/.I&�6k?�z�M�[.m�6q�]M?�<P����q���Un�\���׃��N��,|�bJ�{�P�@#@�'h^I)��ui���|0�wg�Ş'��W�����^<_���y��#m�ñ*��@���%�qk�>T��]r�F[�ث$�����i��w���a�7��=lج��K��t
/79�JF�݄���M����ü��a#bA��Z��na���]��+��!D��W=�n�eN���АZ�h�'����1J��Z�?�ڜ��&)���}�p4gut�E�U�v�o^�*�>�m�Ll��ij���k�_*�9>�����M֊�D�� ��m�D���X�y���qv�t����00ñ)0�	�~��~�Z�Q,�q�V4�ٝ�/�
[5g6	�Ϩa��+&H���UK�tRhe�er��y��T��
 .�OS�ͮ1���l���qU}�O-@��a��� T�?r�8�t�{[��\����,�D�5̡�����3�R
�q�[F���i�oZ��"eҰ�)Y��F�-��q�b��2J��1�eOZ!��ҕA����h�u=���͠��(��2Mh����U�)�8�҉�ۣ|
B���`�pn��o�jd�"|���n=Ъ�]|�S��Z?9S�@���]�׳���o�W�8���|8H�u!��;g�2�i��GS{��O��5@�G9^(zXwg�kz)4�+��e�@'����̈T������)�&��=�ӽ�R�X����~Te����^���e�.ݯ<�l��ڟB�n���"�C_������a���9�2m��_�%���m�`'sH��YI��O����q����c�W���{Z�X�
]nS��"�xztDlf�R�D�����:�r�{�d�N��n��
޹-k�a���{�-tm�#�J��]����D^��ߺ����>��k��|�p��N���y�w"�$�ѨBͯ�7���(1�.Ӎd����u�'�:�m[���+F�T�!Z�Ɏ�箰���Kq��8wxȑ?�+s��=�g|�5_����6:>���)u�{
@�[ػ_�ؙn��6rĕ����sc�h�[��� oz�4a��z��<����'o�p��54��J\$�p�gU�� J�#YPʅ���l�ȕ@��T9�������֦<�1l��N���(�T��l�scv�Ň
lKSS?U�sy /u��y����EP2��S��tR:̤Fr�I�=�D�3���^gHS�9g�,K���c}��v&�8mg�z�/_oG�/aF�����Z�+6����;�����m�T�~��884�xh�?^Dt���|6O)��z�[%L�é����ee��|������_ -�e?V��cX�)q���|ڙcĜu���fIrw6�1�{4�%V$&�nv7+����<Ӈ��¨�#�)wћ��A�e��V�z�fW��4�J��
r49U�c��w��E��e�wz��Jt1�Ԍ�`�D}3P	�r�UD#X����߻>dT�L�l翃��.���~H�KtsZ.��A��گ����3J>�/ǿ�2�Tָ8GS/a�66�-��b�[u���j]'�&��<�fO��&J�/��a���7�V�KZ�M�'Q	*�qp�:��ՊVz�|O�Q�����v���{��u1��b��4����K�0E�%��&���6H�y_ԑ���x�	t�j#^�\�[qHYd�:���3,�ߖW�]y�4��F���;5 �=�\PYV^�H�>�E��h]n��/�"^OX]'D��C�0���u;�g����� ������u	��5�j�D�@NU��=���J���,[͞ܠPFk�V�*-�K[@	4�xk����\~R-�\VZM+����a�^d��R����&����/���K���^Q(�^��M�a�#HO.�k0X�pr�Z����c� �z�0H��Ia�m6f�m�O Ѹ��3%!�ل�Q0���
;K	)������	Av���k;�:��!�k�JĖK5@� ��*Lz��5�O��ܲ{��c�����ޭ�Vɿ��MȇP�	tV�5�<.�2�WQ[�`��
N�vP���8�ix�>�Rۘ
��Ŧ5�l�SoC��lo�D��Ǳ�n�*�g�S�"N)���x{��TC�D�tC7N`�l�uZ9�b�h����T;����?�K�xJ�
�v�P��s���(���62�~��@Oϻçx��T�*-�yTL��'����n��n@ݳ���%��K�����~�e��� E���UWx�����a{4���})҈�w֯�~H�Y+�E�ζ��L������8ݽ攏_b:������_sae����F�S3
0L 4�̷<�?5+��? Hs�`�9�Wz�:,%wh��4�e4����>�,��m4�+��CW_���!����uC���	,�x�ҏ���&� ��k+n۬l�'��K~�x}�����~fy�����߀r�y�V���J,`�1N}��r�m_[]��cs��v�a�+ӫ��5u�O�Q�w@���f��p��$���ΟU��1W���b6��������q�T�Y��'+w�7�S[͚dw+P� �N���r�T+f �Jp�!�:�l��>���4�16�%f�A���6��C�oLX!$��?	��.�bs�Xֲi��^Ѩ���__�B�9%��^:`'z�a�_�y�7�qM���V�?��P[�/t���&�����C4W9����|x��	�*E��Ni��؀RF��	Єy�SY=z��zm����'�:h����K�77v��y���T��M{�лC^�{[�f]�g�������%���'>*�Ar��d���e��W}���O���ɐ~�T�I�>we�+A�ܦ�rj���� �2�u/�t�����������F(�};
�'#�L`(�������1y�Q�r�/�w�L̊���G�e��ٹ��ȓ(��g	R ��6����j�~�"����9�&\�����x�/"�V%�۪��l�4.,��L��9��	'���2�e!u7-s�{uB`<��@Bni�$��.��{����u�̨r)�j"^�t,k��SY��H�l)��Jgw9G'Y�m"���7��p2|O���a��(����L[���Mu�# kM�\��0��ŀ�x�&r�7�����6��n�8����tj��E�tjق�S"`o�M��A��*��@|D���4�G��I�K<?B(p�[u,�|��HaT~�&�g Hgz�ςY�*d$5P�_���t���Ysy.��� �~��E83���w-����ϱ�m��6��"8C��<^��U��U�;1�5L����
��*�ă\p�roO��'} ц>,�8�}�J�z{��H�O���g��%�� �n/u����	u�#t����1�#�{���۪Հ8��;���)DLf�(�{�u��ٍ�h�v�D�t���%�o1+�����XO���(-*��/�m�Ty6�Q��>�L�-i��я�����|�a�Ǎ�i�q���P!����)�6�(r��T�=��移)tu�AYT�VuO��Y�6��7�0l(1���0��\I���ܹ�M���ee��(?&��v��Q�؝:����cಠŒ����kr��Hm"�0���;V�U�����ޒrQ/�W`Tz��i 㳇�}�Ėnpc��MDU5�|`�d�e8Z��4��B�VI�y�p|<�3Wi�8�P�Җ��>��W�K�"�]{j���
���ü�}��_Kܿ��"��C|IB�A��>�#�
`�Yr�h���W�0��
������r-�8UHP���-ac�<��HϨ���9�\�ԭ�
@5���NL*�*	q�f��D�U5T�\u�\�k��*�޿fyN@t�Z�
�P���p�C�d��n�ḥ2;8n�2n�5>.p+�IS&�J����'O�3�}���.�����>��zxD�=�����f��������x0>�;i)�	�S-4�Z���?_Un�����d�������>T��}4�S�n��2<k� IyrrDL�]������.cV"��:A�itëW^ъhSE�iV/�D�$	�?0>il��FS�-j�A�1�.�j���7���W�&sF��U�f0�-qF|G��ز"#)��;��<P�_n.����et�5O�Lv�wHӖ���أ�����I� �>9�;�܆��~-Ҋ����o�?�Fb��c��1[+C~;a�Ue��U!�҂ϭ�m��4=��;P,3w��������!�ٯ�;��$��Ж�E{���n�ǩk=E�(M}ԧ�+{e��s V ��0.�guv�T;�����[e�Y@C�Z\}��4�[L�t��-�X��Y�^�vS�")�Q����%s��������@�&��%?�2�"}`sb�n���$4y�-��W�*��jb��Ok�����p��/e��u��Fs�c��#�ȁB�Rᢧ�0^��|0��n��];�7�b�T
:�;�(�n���ܕW*ڔ���Ȥ-æ}���J���o����?W�KMp)��h3}����w�	?��7ͣfP%U��W�At4'ýZ�Y��Zd>��*V�҄���|x���:Sl ���{�Z$I�
M�R�o���rpSg�;�xO��<�?|��7���V�x1�pzlVeZ�sG�8���ʺ��.V�%�ƭ"RC���F_ĝts��g�*J"W��`�Ϊ�Lc٥�(��0�s� ~	�o�Yp��ܳ'�Kv�+��~�łL�@��[Q{�����;3���.o�����/5.9��\��ߗO����beW5�Z�4fhc�k��q�J��P���J���I�ˢ�l�l�qp�\%�1��+�ܘ����4 �S���%���c�ݩ_@����;b��&�����b��7*������P��ˏMRt=�j�E�]em��L ��=Z��:ck���z�Dﭐ	��'�|� �� @S���Y�Ȓ�e҈�d�8}��'p�#���.Ƭ�ZE\5=�o�Aw�b��Ų�e��s�⤝w:������-($z���M�O��i�P	��Jb�a���w(���7G��,�(.�<� �:עmZ<�&�/o!Yhi�v��Yh��t�M�[�U%�.,{\���5.]�BɾȞ��Op�dR!�j@��z�C�WH�����Ʌ�I�g�i��N�;�L�K�y�m�7�$��}
 �k&T�ŽB�X�S�6� ����$6��%�����ױ#�=ͽ�" �P�πrW�v�Yn��S�ʼV~G?n\YKo'e�K�C�vQ��^n�E��ৗ����Ձ����W�~�hfv���Ӥ��r�
#8$��8O`�/x���Έ��a����7ZCA4�♯{�&�g�줖�?��ߐ�Fi�d^n�Y��M U`�.�]�e��=��	�J�"�85Rŭ���\�-V�GJ����J��yL&��WM�
J��E�F��z��`�5�N���b���3�yUz	��9��9�߯��g!�C3�=y�MŵF�����`��/f(9�ũx��]ӽ�*��j�Q�G	𕖩�� sa���]i��Z���ͺf�fm!^Հ�.ALB�����! deY������~ƣ5I���H��9�B�Ͻ���������뙙�46�ʨ.ȉW>�E̹7X!�[������Bg��P�[?Cݩ�b7��YjfP��D<s�>�;�cs|Q%����&	~Y�>ɴ��r}J�A�9G�j�c�(�UVџƭ;{OR�{��x"�_��K�#����l#��A��q���i�w��-e�w�j����tQ����noJ�~z��b��~}����^�8E�j�L%���;&/��7���	�����
��5S��*7,-v���<�FK��,sġo�,COb�вP>�c�3|���E	b?���/�W��p ��dE�Ә��S�Crs���
�����:�(�2�<P�H��d���Zp��R�R���-*b��_��Q�SL#ox��~��C7��L��;G��bH~.g ~D�id@�(��1�[%��0	o|$����+�}8����?7��?��Z&R�����4h'mY �W���k{=
���:�������G	`�b����U#吗\@�Df�a<{A��i��l��+�����݁��/܈������2^!>p(s2:8o����"2P8m���C�vy�����3���<pV�E{w�·ph������KN]�|����]1�ںmF߭)&_/�d�,|, Ӗ��p��,���Ų�K7<�Q3��5����\H$�,:�Vzԏ�&1 �S%+@�u���o�<Z5�����uZ��d�:M���˽�c��On�Ĥ���/���i=�4�Bߒ��I샼?��h�%?CRs�t�5���!��,�wRĝ�|b>�\%�e�|a�L�le�;�0덩�{�ټ��ݍ��?�R|�N=�����D,w�>:��1+�x�yb��[���+�Lw�WY�D�e��&�E�Dȵ����܌M/��@şe�����.8M���hk��!`5�m��G��q4��
=X&({j�|��֌%��I�"�ly��9�A
�������o=�R�?���0GO�_�Ap�G��4��E��ǜ�bhW��f% +h]ٛ}�H�M#/~Z��W[S�p�L�UA`�MtǼ��#E���n'�g0_����Q��89
9�݀-;6yпouwHa+%,x��33��Q�`�;m�?�U���B��K�V���v$��X����b��~q�b#�h�A#�]�t���Gr����A�:Ws����׽N�ĆOz{W�n�j���6u�`h��mCg%:v����4cr�����.�0J���0���h���I�ȳ�*�����WX ��dMՑ+/�<J3�M�qo�Ϛ�š�O@*��R}��)!˻�w.�=�'��U���$\�9��9���c�b��M>�Qx�zZ��ܔ���y�T�[*�jd�V��[$�V
h8J$/��V%/��2���7H��ҷb_�9�f�QWO�r�����SA\�6(�<�:U��10��hJ�p��OF��wI���&Oqlh� 69��E�,&�`m�D��Ak�S�R�7�Tˣ�$Lr �WLJ�!�Z��Yl�<�r˃�i��~�Ȯ���Z����c��3_��`�Ep����`�f�`-c����8�w�dc[r�J�kAU�fD�~0�=��q�@�|��8+Fa�u> m��+��>v��"�og�ܾx\�jڥ�����C���<�@��0�i�S�B8ov]}���/W�72=���uTPU�P̱GĶfħ��K
����[ɃG�Tp.vH�;�㻣�����&��ӱCΪ��v/ou���!C/R��%�< ����r-��A>�^YPc�/B#�Hp��V�LB$jm
�O Nc�A�+��f�!��F�"�B�C�Z�^
�i����c#�p�Q���B&�b�vQ���C��_�� 5�#�� ��7xo.�;X}�{�G�``�j�x�ÿ1r����
��>h�G��a�a���G{�1���#��c6P��3����P��<�*<:����P�J�|7W�ׅ���k��u�&[̺*��:/X�E���CE�(C���Z״Z	���)Y�-���Į9��/P��� Ncd4���8 �f�m����������2u��VE@�'E�!m$+�7a�jJwk����dњ �r$�VnC=�vlLە���|f���iR�Ė��$t�zvg7�"�8aR�m��΃��d���lТ R�|W� �xs�D�
{-�ҤJ��%��)u�X���@������ih �'g=��lr��PB�H
�$>�+ި�?�)�Ѱ�Z�"����������_};˗ 1f��	@�����U����P>�M6���z���יrr�����ٺkP]�6�7�~�M�h��*�׀�1Yɝo=`�a��ĞF�K��d��V�)�2UVz4vv@r���l�FP?ԓW�ѣ�9ܖ�N��R�#���]��̐S	'z3]c��>�R�$vk�?|�1Jn{�w$�*�B�b�z�)����͵�??'G��.
�'���8c��-o���Q�B�1�h��&�����5��-��o֯:G�q�a<;�u��vܹ&�1}C"�$����Vw	�BB�����2�F�p�:n�Tp+�1��!�e��CA),���CQh��'��=��a��z̲?�}��""4FD8�3�p]�>��Yf�kyt]��_˜|���j�����l�����>��ג�dn3�[����i�Q]n��%T�^za���=�om�>��=����,}����P��@G'� ��Y����_v��d��'��f]�ۇE�H���
~<%ܟ��ɧ6�z�k�p����_Y�Q��`x1|JI� ��ȪR���V���LO{�c�h2p/ �I~�?�'�1�:�'cȼp� �:�=W�J^���S�`�xIZ>��P6w�U�>]wC���"���^�5 �����w稭6��dU���%�oV��6I�YZ�eЀ��H�D���evz|(%���j�P�mH��b_�p^-��&�Bh��$f_<�l,F�q� ��E�/iȽf�CҡXt�:��ZD^o�偑�k]:�Ɉ�T�ºIv�f���L�J�U��*�s�7ܢK�:����B�RoG\'��<�.y�@n��8(���g���@��wƆՆ�	mF.J]n��DY����by���g˹�����Q�|��( 5��W���a�K��p�W�~��lj'2�Z��W�=J�ҊN�WJ� ���`�����2��w�`�t��p��L�ӌJ�9Tē�q�N��0j24�ZV�,��]�9|��G+}@�L�����>wY��J����vޖG�E	�@���j��!.����~�.�e.��wj�]�O��,�#�>��<u���ۗ��d��Y�����6K��3G�|J�T5���j�`��rH_�$�����L�N�Fކ�琎���ذ{����u[ȟ�L��]��&J���0��Tl��H�����ɔw9����5�8�V侕(F����d���Q�V�<��,,��LE@u�:<.���Hz��ݯ>���5��R7)�
�T��$�X��<��fm�"?��w~�,ƀP��v9�B��K�up�:��-	�3Jt:�l�"b��Ɗ�j���ڜyQ_ 麈[�]*{~��ΦMw�3u���7���K��HoL.ԯ�� H��+�9$���\ϒ�=���aB&I�k�1���nEW��;�$m�,�C{��&�	��1��, ��i�k �N�%�w�ۉ���}�<V���C��Ġ
u��2��2a�-��S���f�L$���cq@ePq�m7�e�-�;L�H�^%���m���[�nnT3��|OR��3�K.*v�?xj2Y�ˎU=�4 �h<U�uO�����
��Q4�|�����3���O�F�V8Re.��{��=1۷�PV�*��/-5{Ԍol�c'����L?7h�:�ɠ2'������TN�H�I`!��R�X���6�Y��[�mznHM8Hۈ)�
	G<Ɍ�!���V$���V�o�>�eQ+|��Q{����w>�g����u��b�;����`�<�Ʊ!pl�X(���O>�$�')�cCYb��XR���� �G5Ŗs�لA��F4�B�����3gV���T�Fr&᰾��Es��7��� \�!��W�lM��͇�o�����e�_S�ii=�NJԓ�a��W�I��Ns��\�4���? ��	�3H�gW�W���g��6&�'7�рX�Ĭ� �z���۵>�e[j��wK(�n	-�E�����S�3|���7�r-j���~�h��JSE��̤����R2+':����ʹxb�ǻ�w�;�j���[w-��( ѫ�Ľ�6�-�-��LzŸvƂc��~�x\$S�YY4�3�k��Ԣq ��õSp�q"lg�\?s)��W����>�
��ɧ3��ds`P[`��xC)���J�$�OU�����'���5�k9�?���[#�6������k�^�ܩ��
�`�[$/;L��l =� �C��w�y�S�X��~H��L>��0¨�O���X�1�j�b������^%l�+���:)0��p������$��ƅ�Ȏ��$��&���pG�y�З���;Y�Z��6 �L�@B����#E_�P_���+_�Rx�6�I�$��L�5+V,RQ�{q�`^�J�����Q�<�\6�4�XOҰ�F@ShC&o�n�}"�D0���D���] Å�#�h|u�S���QlB%ж�. ���ް�[�!�|:����F��:�����<ߜ�c��p�n�V��YZ�/��p��A\��e�?�ǠU�`c��d�E<��;y(���� Mb�����Z���@��d�\�f��z�yȠ�/+'.�[�R!��Z�X�$n�xU���UҲ���րD���"&��v���3P7����,�4�ުrPp��:��%R��M�$��L��3������|^Q��(���&I a5Q94ޞ�0��������7�u*�� \��}�ض$p�Ru6k���gp�E��Q����T�P�|Ks�\5�
��ga$��{�v;�������ۓ�\ͮ��qb�a$�_Ю^B��r�k��s'7)dAWW�׊0_���2�Ov��K�%����2M���@�r�Wx+qy�z|���7>W��/B~�09�,k_�ȿ�5Q��A�zǴ�7�\�C�^)�i4��ۮ�y�f#��CUte�U�U��uff���9ث7S$����ڕ���JfڴlM~3;�&2ʲ�o`%͆����N_2䧗����9�+r6�B��߶�L:��*��M���;�l
�ו�U�b�$��X�&J�v��g�{jH���8��DlYO��+T�E�M�"jM)(��kU����#'��2�<��D�l7t�DQnW�c�lY�{Jd����'��U�����g켖�}(�ş�-H+�h'p(�w��s#�b�ɼ�?0Y·B���-#��0u�T
z�ߵ\	���E�o�e��<J"�_ݡC2�4@5.���ΐj��?3�eķP�O�wו����~���G�VE� �8�T}aA=��~��>�jBH5��	�	��'�=P%�+�]2��i���n�w�]���9�% F��gW$�X�̒ĺ��.< nͱ�!�fm����-g����������{�D��l`�}��� |x`��~�g����Ť�@��uA"���#��,���=�_?MKP(��1�k$a�Hp�疟���V#;�b٭I���0�P10�MLLV~v���w�~�5?���W��i�wxs|3X�c�M�Bx�Л� %�;xI�K�"�+�="�")�+��A+'�ŸUz�����n=� �'UlIO�1�4�)�]'���g��V���K�φw�c�ز(�K�&������*hL^�R�Ɋ
����͵�<��灵�r��۪��&.�2�D�463ߐ߷vH�ӱ�)�1�u� ��bEŖ>зn�,��3nN�z���$.�b"�ԇ�V��f2.�)+X`U��t)y|d���V�2�7����<�i��LF$�T_+ZG�����n"1�Pg8����@���X�c%
���U�7����0u�me,ހ��X���J,�L��,ȶjY),ܘ�`�ݤk�'s�{�����o��~�Ѭ��\��e?4�D�{kB'�
��>�9=N|�4b�fy 6���~C��@��~��*��U���
A/��1��*-G��?�d�!��9���(���TFS��i� �3����d&�����p���oq&��a\]4زS�1������H��P�u�_r�ָ8�$����gW@�/�b�dE��۝���U;*��D�N{�� ��'�q7���e�3m�%re�ۿ��m.��<&誐��ɜ��lB*�)^Él/絗*A����h,^&WC���{->k��Y@��$l�>¸X�!y���x�A�bb�#�7G��$�L��&qM>Y�p�^��3���@�$�GZ��^ �RE&z^�`�en������P��=�Rr�#�x���Kn�Ω�s����/�Z�5i"����W!��'0PҚ}���7J�	7�u�	���;�&���s�}�n�[��z�t�z�|�X��z3�]KA�Q����ru��\�Z4��z���Y9��������>��Xx���-���^<��Kl/l�R���bR�C�����h�q�:���D�5B�7�<�ݱmJ�zxs�?������E2���n��0)!@[��I��/3\�>s$	�~u¿x,��;�h{��e#�JimDd�SX��ݓ����r��-6��BiR�8�-��wB�\�4��N�S��Uǟ�4�1� ӏ�81�nK�^�0�s��'7w0o�yAK�'�#Ұ#R�upU<(9�!��ZBV���d���e(U�)�jn�1o&�0���=�X�ŵ��0K��s���� lO�����PE�"�o�8�#e�#�r��d�-���o.F�#@&jvoB�˪��wR�$�m�J���|g�^�.��x��JM�Ǘ��O~/�z��7P�A=1��������Z���E��̹E�s9�iB݅�t�������r��?�N2�K"�X��&ꞡ�"����=1�Onr���scW��"��S��'X���:�Q�K�vl#�Ј��M`]#���q����h�t1����g�#Ð]
 �'YD�=�U(�R�hPt΋����+uZ5�؉��a{�v+C�)�?�b۱�cj��P�����L1T�0|�G�) �s�2�9���=c��OI���⺏�Wژ���f��ˍc�#��$V偓cȹ���b��}Zd�v�/��4�ԭ�����7F���Yq�̳A[[�H�)c6�6��l��g쾥�+�n&$;�#r��z\X�F
�6��rC�9i���se���N��	p�n�B$NA;�gr]�㐦�>�JFJ����qʉ���C���v]D�x�:2�H9+->aZ���&�44F������s%=��B���E��CE'd�v큭n��K���dy�&%����G�'L��_CWă �A� �g�"���$���7�>/LU�����4�D}v,���U$Ix$�v���M)p���[i�S�rǶ�P['��S�!�>����xh&6l��K�������՗;�kfo:��:Js�b:U9����H_���˟��#�Ѡ�(cf��kH�q	C	��%�z7���P��Q��sptL�� V�B���hm]��*	�����mA*��`0�%A���eb��K'e�찯���=[�dό2���!��[�[�.��q�j�	��u)l�M޷Ĳ�Dp��<�b�g��N��r�d#���"�Ҽy�1��� �z�1��1D<��zY�J���/��,���]˸�V���q��@���?��"�/1�D�Zr�y I<Q�}V ۩�f�;nF�د	n���(w\�Ŗj�����)�.y|����9��DmN�^�bJ�׫;�Ғ�4rR�D���QZ��[�kB����8�M�71�Q�)�V6wWFeE���^8�_vߍ� ���ԑ�ToyYw�o>}���{\�k�%
j��mM驽�u-HL�ڵr
f�9Ѽ�x��2=�Y�G���t�F���ˮ1S����c/v@�_!����D����9��8e(Rǌ�����dn�boõ*d��n���3>?0�����ɸ�����7���#�gK.�Z�����+�I"T�,����L�F/C�B%?%T���I�a`Z�����3�X�i��6@Q�f%�s��[E��+����PT��|K�vֻ�_G�'y[;���nT���
}c� �ӡ{��}���v$�l���z�8�3=����~��Ef�z����PxT��T���c��!ܴ���P�;q�p�P�� �\ �?���u���"у��-�YE<i�5����+'���q��SC�a``��@?�>�{��̞�Yi��-Љ�U۝�}z�s���>�tZ��%x��LW������*m7�<D�R)�@�]����<**�Ǆ6��Cqz�s���yi��c-7�����������<�ޖ%��������ɻrn��˅�Q�y���J9NL��!��J����n�в�h ҬT�"M�q�d��d��@��G�\�X=��z'��qPt�!�i����8�i��B��q�	n��ޔ����0X�שt����ک����:f( �[�/��.?ON�i{��.�}T�
+� �s�_�}��P1�Ы�HJ]�K-�5ڤ�����M���Z>oj����&ku�ў.��K jHL�d�s�� x6��g%A�5!"��BՒ8*�P �!S��MJ�S6,5�A��9u>�v��D�T��M���9��U� 6�ř��F�x��G�{�k5����:g���]����Mv�o�.���(.o��|�tŤ���d{e3\z��(n���s��-�ЀL���<��jq#zvp0�5�,����������]>k�הT���#�VG-����4�;�ǻ�\���6X{=|>�L6N�4�8B58�>H���/��Q0I)���X�����▐��9p.P� {���@j��k3�;+Fp/���T�̬�lv�[Ɛ�<bp�O��KK]iB`��W&Q3ʖ�/�j�Xiֵ
6Oi�1㢑2��ꠔ?��񏖦��ۆ0�B�ћC/��O�x�[tɭ2L	����ؐ2o���9w�Mj� +^`9�I9�R��X7a]1Qn�$��s|ٹZ��.5��E@Ưvp��r�%���_'���YU�>�#>\�br��Kq��ި��`�?�v��K��E��FB����'=���ErU�m-�FK�qE��5�M<�
�z��d��I��0/W�9���;��o���ʠ�O����v�Yd&B z����E>��ɕ��}�#�D��L8�Z=�f**��c�>�%�z0�F�ZP�*��SK�����N/!��u��}rq��u'�kgV�����oC+h�~5@_(4>����plb����5����߅��(E�p���i�16�����o����_��V�����| �c�l8Q��v�db��u5�ZgpO�m��r�s�$|�m-gɻ^u�Tȵ ���diȅ��5�4��i�=��/�rF;|��W�ןPL�����~�y�v���{
@�{lu(����:���f\��[E��Ë�>K��e�	�:�sfڵ.�Z��k0b��$q�n�8�l�xל+�4�G�a� ���%�&���	^�P-���5X���f,Fj�(Q��J����`~9�jn12�Utfq��hH B\NIA������-�"&N�����ͨ(a�%�J����Đ�Җ-���dV���&�C�&c��;~�/GXM��M;��Q�������MG���n���#%�>�w���R��rP�i�"�F�ύy3�֘`�������A�s�94=!�{8�D����]�,oF��;a�O��A[�ߜ�'&(Yoۗ���'�9Eã�
��X�/D:n<�H&w��*�`H��)?)�8.�H��}@��S)�f�N��0}���q��D�s3�Z�jN������H%��DN(����w�:��� e��,PT�����
ۄ���M�@nU�ul�#�8r�u�D^5R�޻��`G5�#���ƴ[���Z/=tI�qr��P)b�p��U��V\����N�yd_��lv�A��(���j�>������d���)x��D���*y�?^1B�u�M�g�L��R�����Z/��=�����ɫ�|�A][S��*�5�pՓt�Ct%���B����ݙ�^%�"��C-^p7M1���r��Cd+ H��!�60D���L���_ӥ��Ӯ ��W,�wGS%�_:�ǡ����n'���o�������y�l�Q}�(�ޚ��5��7�'l@�@��ɯX^�~�߫�ܸx�-P!���Ql�Ab��CK��T�N�6z)^ԑE���_��ׂ�=m!�t7L��8��S��T���o&L4
j3]x .B�^��7CZ1ak/��0���G+�r�����H����hwl��;��o�SP��o~a���*}٦����������6{C@�@�"�Y�C�@\��S0Wm�^^����]��DTѾ*���=��#�Z��7�e���wv�g��[8��S�`3�}���@��YY-x���/CxX��_ۃ�a�b�q!���顺сq=k�ٯ~o<������;Y�9�Z	r��?�QC��1a���h�F�V�#��E�y0+/,����sC�'��1KwX��³0k��?�.)��7�m`H	��;���"(�Q�f�� r�N�Nڭ���IÃ?�f6�`�����A{*�zشySy"i�u�9�rܺ�F7��I�mZl��^CIB�A��7o=|���m�8���0�K<uD�*b׋��mr�yW"�,&��ᷭ�j���lUqّ�}�8;�,�C��;5C���1`�.L<5m�%�xXu� �q<y�7!e~9E�b��nQQ��ێ穂�n�1���	����|Rd�Q=Y�g���B��␴�9�F;�c�����N�PĂQ�Y �3� 74��X����`V�Q�}��(�=�$�K� v6��~,
�@�Zla��~	hWV�%V����O���PY�E.x&%,C� r
��G�&Wʫ#�N*{��G{JG�1�}�*΁|��:�td8�!��?'�������e��Vr��8��僆����Q��B�r#9����7��O��r+a�h�|}�M񧄽z%�GÏc�hIN���},�`[E#�s�#ೢ��q"+�d�7�h$�+<rȱ@�8^3���8"��@L�x��L�Z ��)��|���#��&:�9S�o�q������W XV!�
XC���_��o`�7���ލ���(r(�kg��/
��<���QW����J]��8��e�#�r�v	t�lDn��zr��u��G��T�h����!o�=�s#�t�@�G��f.I�U�jQ��0#)��T3�יFӂț�4[�)=��k�׹� ���ns-��I;T4��팸�a#��m�&���c���Z����[sz�P܈m���u�3����6�,d-��1����Z~[�������U">A+� ����o���L��̺R��7�ڞ��,��P��=�Wdf�����RU��x�W���[�S���lQ�?(є�����La��P�;hB�p��{B��/BВp��������h��r�Z+f1�-k� ���-D"oQ�3�3|�T�����ϥ^y���)��m�/װX���t��gM��.s���`+��;�7AQш�L�NKY�+��_��I�
sP%z� c~Oe<r����T.}^+IQ�x�x~<G�P�XF>�����L����i��.�D� �1��1��hB��F��+�!l��|�c&�6�JEF�)(�P�]ԉy��)j0q���в;���>�A� ��� ��eJLO>6�p�"~�8�z"�=A��Ou4���O��o��3�9�׎B����+��;�s�H����nTuR�J�����h�Ӱ��wh%��'����Ɇ�ɸÜ�x��D���{��7�Cm�m�#A�D���y�	�ޡ����!��S�X\�5�a�9}���ilk<X}k� �]?!���W&�U�%�'�:�9-uF �IMe-��N߳��`�Qi�w�UIH�s���h;F����H��$����QN�c�7!��f,�n��z?U��g����E��&�A^yCG]`�O�!;T�0b�N�2�%��VZ�uٹ���E%��M�@5��	k��'.\��@�N���?��XEy�m����������ˉԖHG$����L��6s�Y���� 2!��w��=�Uw�~Ę�I�-�*���������2J0�,��,d�)�{3�D>�������ee�9�e,Ĺ�M8�_@��I������t�g�av�C��JZ)�8ZSW��*ZH!�����2�;�ͣ�&z*�o�U��QۋOD�n'����S1�)�6R 9~h1��m������&2�B��M;ȩ�@5�S�V4p>BIxd��>kuQ�n�N����I1�^?O׃�%��2vL����e`���_�+{����;D��Z��^��������)='����j���7�5����:Ƹ{��OaM��8�8�uo{�+
�Vr;�Woh&�,{t�Ⱏ���	��؎��]V���@I|FՃ���M+#�gK#<�������7�ޛ�Y��sh�Cc�Ȫ��D�j���aæ ��}�G���� E���[����$ ��#�<�\&�� ��Do3�q����L������I�Y%Ѳ����J達����Nf{*�����9�#�.��z�q��^��o�5�t�K�"�`��\����+]�xv
K{~�n��*ж��.���&N6�S�"�����w�~fݥ���I'�Y��P>C5m��F�L��,tґ���g�"��֙4��T`��n�:h?h��+#o��~�����XP��W��-Aazlp};8�W2��u��Y�����awZ%Zx�]�;��j'Kx^Y=��E���Fe�z�;ov��ֺS-��'>�oN�4?o�O���{,a��Ż���C�D�u1����R�H�\Af���WШN�|k.{M��7Y�%s���~Ne�M{��$*�ۈ��AX��Q����U�-��ñ�<������zPb��l���
7_��\]�R��'�B�묻��R�����6��z������1�q!������F(�E��t��I�y�u:lj#%�bE��u��`�����*"�������A_S�ī���jD��
q\(�y)�����^�<�UY�'x�G�3J�/�h/���U!�K�?���wU��R�քv����]�Dd.js�u��g�@��"���4�o��҄�#f���C��&�_)��R�Z���.��[iR[��P�IC��m<���S����K\)
{�I�'�?��k+V� ,�N���k���u|lD"F�a�mɪǔ��G��e6_CA��@C�:�6�}���v�Z�<, �*&���%0����]�܈��o��Ed�&I�;��pP����$]�1��_-�#�3�P���@Sy�	0����jT�C�}-W�iﲚg!H@n|����O�쀃���C��(�Z�F���0����Z�2ǬQ�e��Qh��G1e���xn�������X^iu�ɝ$?*�pB���>})�F���n+IO�w4dYR�fݱ��(�����2�w�d"?ڥt$�w�a�ۆ�OE�:w��~7!���k�Z�i`k�4��bK�=�b�	��c�!!����a�w�A:�ӫ�(eL�6<�L��4�C�<�>ДG���j�,�]�N7�Խ|Y�o��Kea�K�����QxuՒ�-���Ž�E���.�X���6Z��b�`2V*�;O�xP��hUB�7��H1$�*	��7��4*ی���=�-�q�$��^�k�]�'�����xa���}#a��{�^�6c���DV�W����>c'ʑ%`�9��A�����gL��<o�Y<��Y�	-Z�!o�X~)̇�N�¾�!-*�w�,�b�ܡ�m�d"q5�'K���x?6BK���n%���nP��"�&y���-��r�:�!��ߟi��b)���?p��� �̍P����KN3���'*c
 #Z�W��\�J6i�9���82l� ?��2`,ag�h��Fp"�Q�t.��u��ႇ��`P��������,��f��h�[L�s���b����4�u.���-�^�:^��N�}�o���9�_�)��@�Q���P�K�<�+'�8������,�k�� ��ST�M+?���!�)�)����ڦ5ԕ�~k�ihC�3�%	,
�3���b0Y'��WP���X!}�������"[a����3�i�*��W�'*��9�Y֨D��������~�p�j���g;�ǈ�K���n��=��W�>�n.��Ñ��j�6,)��y�]	���\)i�+�2(�8덡GH/�[���;����GӲ���b��*A;g�ș�Y����������fv�(����Ո�Ño�N�3�ͼ�>���5*�7���J ��z�a�s��_(�`�f�{�Eژ|J�6�Y��d��l�aݯ-��$+C�!��&(հ�]��Zc��ʡ�s3:>LO��e�v#x�T�)�E�I����tZ��GX���ߤ�$��!�>R��
�浃lt����-uVڻ�LH=Jt��`r���v��z�	��c:���"��ڗ �W�&~��gu�y��ِp����,��O�Gc��j��c|��c��n\m�����4�H�/4(��#f��b؈u`eqg!���W��f%
�w�Q �Z0%�#5�r��-�j�$0���{䥼�@��	1�y��Ջ���_�f�P��B��"����og����#�]B7��*�$��zn�&�`��|(�fo Cχ+;�Z�d��=:P�Q{G���Pc�b�<\b�΄����U�n��ՠ�4럓<�q������is�U��o%�=Q�L#Y��|B�l0�������x$%9�9��ŋh8�&{�_���ʌH��Wql{��t���A$��� �xhĔ��Q��<7ݧ|���%��ns��~������	�U��!��_�]�v	K\��Cy��j���zx���
�� ��em,��9{1n|g����)��gTk/[�Yp,蠆D�0LQ{��<CJPג����]�ݞ�3p-��$�v��N�~<N���5�t3���ʥ��0i�Ja*�W��)-6|�4��E�U=Rٚ~�˛��N��~�5�}��6�~�v�`��k,�$�`"qX�$N�y^��M�f{A���*�Ӿ��Bf�2/��0|�۬���sSG��M�ԗ� _ܩ�?�A�����6:��M�� ^Ww�����\1h����b)O�4E����� ೺�c⛚�|)���vU
z��Y3���.���������1w�k��-��L�$�U��w���s*̪{�H�C��s��NJ��:�vC�F��Ң�WB��=��G�I}��Z��bխ?/�^���^��M�M�h�¸D�;��t�t�:���o�R9�<x5
��EX�EKU��}ѩRqGA&>^z�N�ɚJꆐ��� ��L7�l̆J=�4J}~bm�o���f�pK�0hV�o`g��[dn��/�LShL�9Ң������_��̙�v ���AtG(F���V�;@�ҥP<*P�.��J�倚����Z(xc��� M���
��L`v���?��!o�R�����	�m���p��m��|!s�2e���J�&�8���Թ]
=zE�`J�j{˩�K�p�����>Ai|������qhP�cHC�{T6�M�iL��:�b�D�����3��#�b�D�N��N7��~Z�~�eJ�vG�P㾋�9�T�����S�2D�Ak�����3��5���{�^�tY�	i�C��bB�W�Û��Lax�io�W�Q�q50r��Hz����{X���7��j��`v����?�%��:c:>�dF#��
�O�,nSkV
!Z�Bl�}��o��j��K�[Q��s(U�Q���2��d�b�5�n��N��|�)��6��*)�v��E�s�=���Ԥ��4DaYZ?�FO���ɒzi��UD1L�v�-�c�13�X�i��b��8��ޒ�H�'J>�⹵)�}�����5�7�;�� i��6�/��V�B���Le�H�|s��I����$�g��DT�e ���QJ�R?���~Է�Ϟ�9�o�e�<&5��CS���Q���N�8�H�� ZkT����[kC����´�B�3�`z��]{_�.*�{@J�l��D�ú�<$�`��(���*5�ɞ�4�L�?��V���9d�5�5��Od��u�;�z�xR1+� k�$�!�t*S(/�]��L�DA�}��ν�Ig�e#%D����p�l�W����\�t�b���]��G�)9�\Z�K������˃�`�`�K�X���ץf��u������d�OHy�i<���0�`���V��~�>J�>�24�M3����X�|{~$L�����J����Uυr�3��>{>|>Ǟ�D�)����,��0Nbq�P�H�܅��:ѫ���:�l'�IL�Xl��3aT��'����l"t�b���bpԌwK]K<&"�@��܄J5=����;�ݵ�Ü�.^�}���u�u,��t�h�yN"�t�W͆� B�3y�"�R������D�#C=2���v�����s�_n����s���d���3�aP��˺�`ʴ�j^>^D�Y��
prd�:�a\��{�+��˜a�阌N�8���6'���>�T\)"B�;�!щvp�%��֋��N�p�dbd��v���(��G���$��$)I��n���.Ug|s	�m'�j���qd�*�w��T�c�(���e��rƌ5JhK�����;W�볂d��`w�����=q+C���ߪ��X�|釦�l��}`�	�L����
��A�o��w�3	�^o����W�kwc<4'��jC��B��t���l�3x��M	�K.�*p�ƣW���R�s4��N�Pb�2"C�^��(��|N��s�,h˻k�l'��]Ikbg������)��) D�����,��?7�ź����@7]�Qe_p8�ݬ�Yݥ�d�Ʋ����,��b��<�����ћ����*y:)���3c��*�L�*` ����M����?�Ճώ�M}���z�ݎ�E	 T��K@[�5l����
��5'���� �2���Ě}���|�V��=��K�l��;�R=�I�$�R�&k��-������? t�������1s��?��� �lW�&,X�o)���:s��	��P�H���u+��qrRF��+$.�&� [�7V�먺t�F�#'���YL�z�f^E^���S�c�0�6�C�GgF�F�̀�<��,��.���͵�p'�0V�Ċ:���-�9X�GUP|�������Վ���Nڇ���V�.A��K3@&����޸�y	��w��_Y��Z���s�M}�S����	�%/y���.r��C� �k����Er�P�J�]<�k�0G'��o��.ِ��ĦK����	,W�K�٪���]f��c���� aū���V0���L��̡�n�`U��?�5�����d4t9߆,��x�2��5��Hs�&��4x��%h��je�f���N��q�iò� �!
W)m��%_���Ը�`����G�Z�>dĐ��S�ʆ)�gd6��z�