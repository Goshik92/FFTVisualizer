��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]����"F��{��l^B��i��o�A���Ȉ���F N�
jD��w����KS2JB�!���>�g�3p���9i��o\��;����"#�5]JILcX'��|�������Csg�JV>�j��G!)������<�5���(���V�d�	�$���/ly��p�o�Qn�+���&�/�h�1�����m�#(���XYJ����	�#T�����Lqڮj�n*�d �M����i�D�u�KC~��1n�\U��^�C��$0K~C'"�,�Ʋ�YI�'^K�j8O �Y�C ��Ǌ���̪b��i۪!����q�h��Y��q��g�W��/6C�5���̴F�_�kC���Y�l�Lg�����r�\:�������OK� I�M��	��0K���9DF�>��Aد���i�g0��UCi�ҫ�$c@��cj��o��y���!�5� Ă+����U�yǗ ����p���H��AϦsg��˭wrs�V��«�H���y�����q�gx� -�U�����e�����k�$۪��𭿍^&��D���jx�
m�Q>�����(�����?�P\�Gd7��}��7�܀.��@j+�'���u�X��O��.N��mD���I-��0N9������?�av᠅K�G�4/��Vҏ�2Hm�d��d8%��H��� �Xy��:Z�1�=�?sY��c�5I�]\8�X9�����dV	��ңI�B�ix~�顪����[��x׈�]َ�<y����*��l�S�4�k5n)?�!�l8[� ҳ�E�@�)x����O�����h��ݏw���GX Ц[�2�Co����c��Q@��-Ynʱ��4��.�x*`2U��y^E<:�7d`J����MO�G���j'�C�	�G�tQ��~���^���\���'~��+�����U-��l��޲����\K?�zx�� ������B"�:�ц�v��7ܭx���@�.���bE"�Q�d���t?1q �xD�K}o+q$\M��f���[��j+��򕲈�<7��i�w��8HZ\���_$��@�Kxo�" `
 �ghPL^ouh� #��^�E^�<xىv1oD(r��[�H%R{��{�J`�$�C3.��@X�D$Z	̈�_�ƨ����Q�����*�������Z��0�j����.��g�+���|lpRDd_�n� A�=t)�m�[֊x:c�^��a��$�|_�1��Ŝ-�'�Rۮ��SՐ,S�Y�vU�����},-�:��L�`e��"�1%�@T�b�C��Q!���:��5!�;	ٲ�А�r���#�'׳B|�f��{�$7��g�����.}"�}6nѽ�*���`ck/mȢ��M{�5�H�]��{��K"lʑ	s���Ue=I�m�LY��by	�\,⨮�r�H��2��hH���9r?�x�T�=�4���?I)���tt��t�L��pD�$���k�[�%(sA��F�U�v�	a%�⾖9L�G��:��B��nF'k��7��I.�D��?�h�K��,Z=f�pU-��3�S�f$H�^	�{��l V=����@7�/���A�����9�v�[w��9D~�|c�{8���Zy4w�h7� ��`���~�����s?�U�k%��:�b���B���8Jʹ�<��a�\_�{V�z]wV$GT�K�_�4o/�>@Z�1��U��l�"vzb4#Z�e���L�A��Fm�w�7�����G�efP��Q��{�2���%ݪs ��D�Е�N�N}׬��_�Y��߉�����X�ZV�͓�-9u����V1���}�F�%��β���>�0G����䊆�i.8��j3/�(��q/��]��5F�v&����D��1�c��h"�g�b�Ot֚#�{����P��B2h7�.!���<��*ңD_�ؔh��;�g]����HȐ�nn�R��� Fc���1*�Cax�)�V{����`ۨ��N6�|����ْ.+��+���ūuc�8���-@cr�y��*5��i�4YS�>��"ˀ�4�d��V����P���btNR���W�0����sC[����Z���37t�ˈ��E��8�D�,���#���%��w6���E&O}�}��_{r�W��H}�늻��UEy10����Y����('C�˭)�l֎Y�G`�~�N\���� ��β+���쎦@H2���~���q�2�]`�:(��H���(4����ω���.�a7A����
,��7����E�7r�@��8�L{��2}r�K��+�ٙ�64=H|�2j� ��Ki��Π�����	0�A�|��4�{Z2����O�k�#��,Y���){���Lrb��j��f��� X��>yA���jC'�p��?l��6���uq�](d��n��j�C��B�7-즧I$��C���qM�N�;'��ǲznf{���T�Q����h������47�S~��������	�e8{�~��|�R��ek*�߯ ��� �i�����f�Ɏ�<L����d]���[����
��bn� �<����4%i!p}f�L95җ�"D�o�W�gY��R�V��6�=F�'�K��֚����g�1u��|�9*�Z@c�f�(��R�G�4ic�DI7�;�J
�v����$�ވU��&�	� � �(wWC+���_N���t�Z��ζ��O�����F���N^�����N�i��������S�Hv�a�$ �&X)C�I���pY�4���_Ex ���0�g�c/�_�=��=t�Y���(J�b�'A1�B#��^��d5�O��c����g���`����!�=qmeE-�a,E�e�-y���!1��yg.�yy���@N�3ʶG��Dg��m-�����6����h�%�v���k�4�0�c���`�m>��Г���*�����}��W4YЌv�򀏖[�����N� WFA�V�ye|�y`����2t������SPa��S'�ô܅����d�Y{�An�	#}�x�X�νN�|}��F����v+A�������.��N(x+��|��7 ��)o%���IBؕ2L���5ֻϲ�����u��oԩ�4��~���JY�H���AT�A�p��me{��>>�iʛ����%��¸��Tl"���������šCA�V��qP�ZwAq�
+x�����
�t1N�:�)���㼎ú��֥��Cl�(�z�N:V˙���r�"��T�s��0XH�I`��|�➉o����s`#h!��W�3���l���H����=T7p���lu�f����8�T�s�n��	�甑T?l�`6j)U�{�-]�L��u��*8��So4�� (����3n��m4�)� �z�Gw�Ƙ�B0�7HI��UͅJ�}+��I�􎄬h��A��Ͼ���?����v���y�P)��3Lt�\���L}oj��֧��~�����O߼͂nU\И����Zw�%�-�e��@�?�K�	���sVK�ρ�Y>���R�@�gRt�4�V�I7��c5N���Q�##�=G��&u�Eڲ�7 �)�yE�r���u��A�W�6�X�bN=q[��L!  �݉����E$Rv�H/�>�'ߚ<\04F,1c�
`���0Öö�瀔�H:V��^�gj9��a�� 9G��,8M,�Y��cy%��d1�a~�g��-q=����yl�����M=�d��=0�g�4kW�����22�>B��.�o�d�X��{~>��V��e˾\���U�R�|��"tr;ӎ���]�0�ORۥ{�[sB�ޯAA�6��3v!6��t�γ"�O�sp��-���5xgH��N@!�M�~�|���"R)�*6	�Da�����	��m[��O׫ˌfi�bUoȉ�O3ݓ{aR�0���S�z�+���X��s��n���Y^F����7?>+��N��ȿ���V3{}����}7�᫠%Ǳߤf���*�J�?c�VXtz�9�O6�
֞��[)� J�P�諗���k��?��'<K��3�Q^H��>Xss�NLP|������"#](t�M��'X�}�A@�w��C�#�K�(>םZ����h�$ƛmz�z�0�<[��K�)���(�5{q,�X.��E�� ٙ�����	P�>M5$.���'�L�� j++E8}��mã�aQ��m�%�='����S�i�g�F b�X��-'!����y���/,���{�f�&M0fd�LƘ�� *G�K�68zg�S1��"�_d7K��"!cY�~A1���%	p�t���%0�k4�T���ǎ y�Xzu�vCg;���+�iơ"������?��ϸ��Ez���[U+�@�����+h���t��5�vI��+�_�#pgGPsNC���%�U�8YGX4���TT�?���0����(��3�������2S���u4t���������`����,	��<<W������ļ��%���?dU����>ϳ�����C�K?7��qL��ٌ�T��&���������*!�g�|�e�}�A��D2D`�۲?f\s%��o��x��!ej2؋�*k���f��^eJ�#*�s���c�V�P�jQ.'L]O/�{VZ�u��KF&lq���-g��c�^�'�+[�MZB�Ҁa(�~��&3rWj<Y��<&g	bd&7m�+�Х_@�|�����-�g�u�p&�$��kݵu����Ya�6o��r��2֝!KO�p�i���Q��?t�J;��,���cM��D	����+X����������p&�Kd��'��s�I������#���;s�m�V.�1�ξ����Ćj�p-���q��|��tA$������ �=*K���h���D䞗c��kM�F������2�¸��_*:AŮY�%��T�A��@�XH��GPn�ֵ	k�YA�+*+q�<���9��-�'��S�F�Mg�J���>s�P X^*d������� ���/����X�4�B�'w6|