��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf��4Oᐢ��\��1yfMA�>bpAo9�f<]B3��SN��T_�eI Ya�R���p�K1p((���*��?�������[x)�~��}�t϶��\؉�bN6%\�~�+���X�+��P�T�������
�lGi
B��}�<�(��{��B�0� ��b��!^�*�>�l���z�;�������)#/P��D��sd��N�X�(�e���*Ӳm�g�W�:�h&�a��z��|w����L/�Pbԩ��g�N��n��T[�a��$3L�O�ׇ8C�ǩ$�l�$��g_�*������zh��]Ƹ tf�)0*�{��<X��߉S�@�����{��"��s��`�̫�y�m
�� m�ϧ[ ��LR�Y�Mĳ���O�5��^���&v���L_��}�Q�_V��?	��@ӷ��<<���mDf�l:5oA�`\�#��ţ��POHo����~t��ֻ�DlO��l�Q`�=S͓�����cB�Q&0���}j������A�.��?m�k�z�L���׎43�c�"d�eY~ (��*����e<x{x*��e���[��z]i�b �q����rՁt ��~pc���mx���W�*�EH���`4�l�bYQb7��6<`��'@'��'�yǩ�ʐ������b^��M���5�<����v8�AL�R����d}�[X�C`(�E��d�1i�e�-4�\"����������mAGx+f�������EA�C�@�9��H�pf���O��-"�T�꾍�K;w }��ʁu��Q!e�BL�a�(�F4d�����o�P���	B����U0A�0���n�n�<G����Phm�]6ī�M� w/�;gҒ�E=�3 �#��I*�b�s��Vv"s Iye���@J�VN�1 y�o�`u$* ��&x�/�;�SJ����%�����!�+��4�"p&�����&C�@��������}ɪ*(�%�W�JJ^����R��=�t��3�7�����@�yQ�>���VD������U���r�Q���[���R"�9CnMq�ʤv���Z%3ŇG�>�{X)����րȵK�8�0�l�]�*|�h_�9}��%��V⽡�z���i�y�,o���ze&���(f!A4n�~�J���hnʪ_���ڨ9~G��~zp�j�\��&yS���s������z7�n�W��1��5髿-v�Q�vS��+�}�|���m����G�u�P�ΖXN�ٙgY#���vqR��]�[�� WDQ�ll�u�g*��O5(7f�̨����U{�=N�� �	��{@'Fo��uԭ�3O*D�KA�q���_E��`�Pr����}س�B)�<1ͺ����i!��dji�I��0�������;���+��0ދb���/Gɬe�k{�|�p.�y�Ϧ��~�w���ǥr,&Z?DI�`�pj4]��'Q5�|b�V�}���
���s��^'�xR5a�50n|���[}�L��O��UI�aG�L8qe=% �>e���j�������Dϰ����w;��[���w�G[<��O�3����j�dV��ju���k��<�<A����|�����ѐ����% �������J�`�b��B���g� o���H��&AhuT\d�%�{�X�X
;J�Q"P ���..�v���O�	V3m�)�q�PR�ʡr%�5ߘrq���-���|�`�$�-�\�􏊉�9$ڒ�_�	��+�����C��7g-o��L	�"�ڗz,}�7�p+�����ty��]j
�޻0�j�S�����Ee�ҿ�����lh�Ob���5�S�O ��C���\����	��:����w[(iU6�������%8��B�g?�����n!B�� �ʿHd�\�۫�#���"+�`�o�"d8�`��������q�Mq��0��~��#�7f#^��ᅉ1b�C�����S����I=[�^(���GLh$�Ue'�'E�0���Iɘ�-�����J��0%u��\0�S�U�, 'S�Er� R�d+��"�t�e+) �0��-�@<�Ɛ�f���dF�x�2޴��`i�	6;G�]��$�Omr?� ��XM��j� V�S�w�T5M�cv�p]?)�&��*��#=S���`�A��g�N���0�nW��hhHd�եt�Ur雝���<�f<@��ö�U�$�ں�'
����0��3d�鑆-��I{���P}Z-<����hl�r�J=?����tB��𳿏e"�͟�k�E��3�E��&��z���5�:K/�jm	�u��f.JW#���m��2������oE^L��k�9�=�n�-�˶�c�lUw���῭:�_� �!�2�r�8��I���ht���Z����b.���W��Z�)T#�xXTC�&�U�ICЪ$z~��@���)k��i�'c�������Y����nջ;����27oBC��,�f�ř(�������L��eݍ&"��V�!�����@L�����������LƆ>�&,٫F���3�m��
����~u��������dΛM����ƀ�[��G3Nb��oᲘ�3�K�����;˭��W��SN��anw�dcZ(wa�"�5 ��M5��ǨJr�0]�^�j"^`�E1��u2��K�/��*G*--��C���7Ȃ�T5�5��m���;����Ď:d.� *�-�4�~�m�\qS�X!B�P2�PG���&�3��
�/�L�Э���a建�o$r�E���ݧ	�%���M��H5���q�ݳ�Pw)Ȼ#�A�������~���P6\Ƿ%�P�7	� 9�]�f��L�cI�2ە
�`����G�F
9s	�KD����9�W���;�=�"����q�:
�u��Мei���e"8��}�$��ut����ZĀ0��`���Tt���Q�� ��Fp�að��X�?���=��Kn����R�>���Ɋg5����h����xb�� �X��#މ�5���R|��?�j�:�a��,��2=%Msj"���a�����E\���sA�θ�B�R�
1�N� f�}������v�����w�vt/��n_�����(n�U�ŒQ�͇i{�] )^k	T����s�*ĵ�B+�����ߒh�J��� zm+m�9�%��<���yT�i�C���Y��7kD��	׵�Ǭ�f��S�A~Eu�Y������l��EV	���<�\+k�Y0vRν�P�T�8#���o^B=@���=��[V,��{��?��󜵑.ݫ��A.`;"���ׯp��0c���f�6���~8�\��M���.n��ӎ����hjy�Ĉ��,c�Ī����ڬ
�o9�^�~@�����3�[��/
Ƙw#a�8���%��fQ𘬓5/B,#Ⱥ?�ܫ1M���D��t�F��mb�)P?�Ȉ�K4��[����wz����U���wx�3��p�;f�W#���-�F?+���&[&��Lu_QUz�D�t`��Z�a�-=,�d�5c��󖩫e_)¥>c���
G�-]�U?��7,�K�����BZ35��u�F��P�ze���b|�%=���K��A��=+�Gu��|p�,h������6�{0AI�v �dV���Ei�lpZF-�x�]��q?,?�B�;�Q��tf�< �%�T��&�cT&RCx��������5��忟���A��cR���x%��}3xJ@��pN�?��,��I򫍏�2��q36��ǵ}��X'��[U0._L]��ݴ��0K����qUy� �bM�`�ԼcaD�:��|�T嶊����i�������6��:��;�"�����Г�T��S�8:�������.���K�����ԟ:ҹN�<�Z�`�H�aݝ-��[���R^��"�l�� �W,��'rS��7�?��w�$���Pc"6!��� t��i�#��4�����$�-}��
!8[�tJ�^=���L��M[�#OJ�Tȥ��]�tw4)�[M���ޮyY���.�|%�W
�����q��ϰ#{P?�l��\7�7�pnv����gx���o}���S���8����]�H2�hx��&��]�#�!Ů��+��{�akw�.��F߀z��A�@e���u���]&�}�e"�36Y�O�IR[s,�L�ׅ;�x����
��ᒬN�'�l-q�2S��q�q�=aΘ�L�{!�W/t.>6n���"pz�.V�DŹ9anKPm�ͻ��o4Nʝ3`�Y��ñuTEd~����*�~ Jq_��0����<��ÿF�?Sd�B*7�6S.j���1�.g;i�T��'�1�Ͻ� 'h��$����R?�^�xC�cC�ƽ"3P*Z�V�6�>:��$M`kC8�,���xp��{��&���b�h���ڔ�)
C-�*|�k�(� $J���J�Vy�o�����n����ͤ~�����mTT��'���N?�kI�����TW��˺h�gb�������Ŀީ�F��"Ldl8��\�=�X0���\�Eq���A�5�S؎ʶ����3ޤ�W��(f���^�xel�g���&"ˇ�Y��y�M>�W%A�Fo5����K�w�i|�3�USa^�&6�c_�aply�/Qh�J��$��_�FB�5}P뺨짇P�W췆��E�BV|��t�;�"���ڗ�ĉ<K{���Fe��?��3��,���a����vy�e��g�>�S���L���!��Hd��X[���{���w> v
(��|�����G>иq��?JZ�<k��!��z�����;R��Ȑ���po9�6�$����0������>y�%d��WF���R\n˚��*�]�3� �����D��Y�B�[�)ɀEW��J�xKx�N���gF��P��~p���M�	ET�S�Q7G������%ް� `�0E5��P�;�+�!��r��Di��/}�_۠qx
���u�ѫ+3������'z��!�ݞ,�+0�x��-7X�X�n�)��c j��Eo���'īݵ�i� dIc2v,v�	�rT5b�3F8��X��i�.���,��u�+�����1�[�����Z�Ac��o�.H�mCy#��P��]h$ݚ֭���S��mb��׷_ �����N'�Lu4Y(�e�����9$/S�z�'F[�	�C����e�a�i��Z����f��!E��eE�=�жv0�r�.�!tomd�f^5�(��>����u�ٺ�e������A�胳Zo̰��������џ����b����(I/: ڞ�t|)���BJr]��80?�W$&]��	��]��/^�����5[*0�qH��/ph����� �j;=���M'k:���I�*�2�kl�J�����6=��/���W#���+/����nl$`I�DE���͆��~��%~�R{v��ށ��YZ�v��5�9B1ir��Щ���<e�l�.��9�֔{ӎGsĐG�	�$���R�W�d���_`c�Oa-		���M��q�P�R�鵏�	[%.�U�T���y��̙����B��l����:�w�KP�Zl�9~C��e��xqZ�{��J�� ���<�t:��W�8��`�n����Ǡ4H���|�K��̢��G�7�
p��FC��_�l����xkb�YE��,�Spǭ�F�bE�Z8�
�`x�d�-J�:��C���8^U�U���t�t�|^�%?$@����8ŝ;k�)RD;㦕P�큎-�X~�h�ba����VOOcV�p��Pע�Jő�[]xA�Q�(��C| R_�>1u�q�����5y���+0!���'�h��oH$*�LgbZ ���fF{ѥR���.>�����)eѰ��8H�ס҈�>�j�=����L���
��.�hjR0�Xӱ8fm���sEwi49��7H� ���J����\��Q�6ٞ��WT{�
���ԳBΣ=H��z�R�kԧ7����\Ӎ+��L@D����4�֤f����]	M1�vC�#k���A �|W�!/8FzS���~��c��"��%h�A�ƽ�)���W�%�Q���T?�{�Z�v��v�6Q{�%�n�6tu>�F!���ˤi	v�D�����`�a��׼6"�l��^�镽e�RZ��"��d�e��h-��٘4o��������E��?au;������?lB(��.d���I��٦Zh�T}	+ˍL�Q�H~+K�,+��9ש3�&p�ȯ��	�e`K��C��:0<��7) �
�����$�y�	�d1FQ
����
�YJG���ս_�f0}�4g��(Hӯb�Z:x�uxm����p�E+���0�e�Y
/K1ǳ����{Ё#G$��qw�M���*���N��\Ɯ��g����M2&Ao�#Ɯ�{2O���/a�ˡ��W�h�@D��Df��S���i�{� `����<9Q5���U;&S,z~12f�GPM����I�Jl�I#j��O�I���&劼�% ���w��&����9���}#�w�a�j�����A*��PJ�P���'�A�̯�x8��V��Z��	�����#Z�2X��c)i$��<n����A�`�^'<O���9�_ ���5����ۆ�k="vn�Ȍj�ˡ�Hv��d�y��|s����3����,��.N�ڮ�oS[�Hr�x��Mٗ�Kd?r5UC~�g��{ƌ��,ԅ�ˇb�%/���S����N.���B͗�Ve�߫sY��I��5v�-�N���*"�`_�?n�����N�W[(p�r!6_��j��"ck�i�U��ؾ8�{5�����7Hd�&�#<c��"9*Hi�%<����-*�1N�����X�M����K@H�E@�����;g�B��U��������I���,� �]J�ȓ��M�f�5�T����Ϛ�Mx�fܱ�Y����rգ� D`U�c��akG��Vu��;v
�*>2`,�nʕ�U��2�Ą5��~�@�(����G]���;\�i���A��K�)>e���3n�B��|d������d�>f�#hFT�IIM����at@N����)o�E!���*�Һ�F}L��{�� �8�R��F�{@Pdj�s*�ލ�ŌH$,$��r�ڃ�.6�����¸�0��~sm8��*) �9(B�]�	;~v*������[��4KE��9LN��:�#��1�����#^��f"�������4`1�֓
�vd��t ���N\H�j��n�k�־y
���f�O�j�
�r���I���䲅��~k2�ʎ�l��	�6���7bg�{�i��q�U�Μ!P��tz�m���Xz�T�R�c�!�g�nd���kMO|؟-��D��qD�l������=C����P
Ѻ�Z�븢~1k>Y����t�P�w3Y���X}~.�'�����6�z9H�����
M�?�~�� >��<����H�[q�*��+G���W7-�08��l
�� ��nT�0��M1$Px˨����?�o�)Z��Q��� x0��v�`x㠸��;��svz[���=�M_�l�z���g���I�D2�v��u[:M���aC����A�����[��I��V�����-� �NC��!����X�KO�o73��sl�����6��8����P���f�8���"��eb�{�jk��tX�����#�w���1�g�a�b,u���C+"�z-�w=������%,��3�a�������7k�\��*�c+�U/UE�P�lĘP_�䪊�Od��:�I
F���&f���(1ɑ�QX��=�tIU��V�y����4�N�aK�TǸ��������D�VWP�u��d}ײ��_��ז�h���P�F�=�`_�q��\-�DU�����#�6,PŤg�E�5�X+<m�tЉ��%�pӠ���%yo�Ju�>��]�煃]�ne!-��2:�����	3��M���e�*���Sw��$u�2��5Z*<�U���B�����u���^�����AzڵT)���\� l�>.j-gB ����|n�~�)�%p���V�@m�9�T�XbUO��QP�E�M��k���z��������hHD��{���z!C��0�X�\e�k	aƿ�.8d��p������K!8'�tYS�+���~b�tle�cc-���x]�ǥ.H��x&�(���_��n��tP�?�-���d�e�х����&\�$��o������A��X�W�#Qe�
h����n�.���!���wٺ��oG �  )�g*��c��#���A�D������z'�>����;{�1��OԑZ|����;܎ڑ���78���%V���@i���	f�<��k`�{��eB۠�1���C��[��%���v����]�Ugo����H%J�������YՏ���OK�3�w��c��wIe�@[(-��Chf7�� pֶ۞��CF��+nΪς����ny }H4��9 �
��:�U��R��?���d���X�7nh魧����l4*�u��*^��.��eٹ��a�g�W�����Bq���L9\2�{�3^{$�@�5MA�&��}d��äT	���톡�Ҋ���f�R��j�_/�^�j׮��W��9 �R_�.0�=�9�9�N��#no���=��|�$Qr����X�c���^�&�\A�ܪ֊2]��%�	?�'��CU�Io�Z�[�]-g"��~)��G��6�
�r���)2�f�� �B����,n����c��c>3���0(Ҏ5'�=fU�9C#-&�f7XV��)Q���~F�(��θE.ӌE"a�g���?�a
�~��a��������yimeJ���X6��"#�М��V-��T��3�%��
�	�~Y��+3=�;����5}��5z �8!�v@�%4�h/	G��6{�d�|6:o2'�G������hR#��Rc@$�F_�X4�W{���t���w��F":o
���;HBy�5���@�����'I�"X��D���/����,�𼓅��[��Ly��`�@3E#� =Go݆෱�|�m�΅)|ҥu�CT&�p:�|2#����/��7?�y��<f�|�Sť�ud�V� t�2@DN��,��J�1z� �Z��(��Kw`�|��FőT�}:"�x� ܡtY��.�	�B]��RF�͙m�T�"V�����㘚ױdtV�f-I�T�����6�Z^�b���\�o�!+,��n���#�/#�.�9��b0���$�W���u��;�u}aw<��u��Ӹz
�^߄���$'�Ԋ�rު����UK)C�j?=�hkX��gWm<���O�q}pO�v�͚��.�z�G����Vl>�"{�ˇ�5'� �?���Ĳ��{�;pC����MIK\dMȦI���}9�;�D�P<k��������7�����>J��g����|(s_�2�����kv�����\T��n���}ʉIU���S^kҝ]�W�UOܨԿ�dQ�Cڷ����>m�1�xrmRsrJj����i�/��@ư�Q/�����!�Q Jj��}��F��o%��f�+�c���K�+ֶRh0f�74� ���kՉ.M�a��������R���2�K
�%V��N��	IV�6��D�ů�`M8�6�����y��;qd��
f�5fd-Z���sp��G]J�S�vh�
��+3��y4`=�=�[}�{*��>��sG�,OE�_4����t��ZU3.A\T�-40$*{D��_�Ҫh��������qӖezn<99^b�n�y0����2��{�� !b����φ6�rwWl��q���fO\cg� �D.L6r�Ib�k�ڐ�S�k,���u��{N��ߴ�cX�Ѫ���i,�x#��Rv/q�ď�:�/_�]~�L�tt.W��*�U1��N��Q��+�ɰ��1#R6k�)��?h���ɹMq��w�8��8��2��ۭ�Cv1�}�!�-��I��H��rs���-٩�leZ{�^Y��ڙ�q�u�8.�Jq�ٻ~�9Z�X8L�o@O!!G�|gƈn�^r�Gnyiúک|��@H��s�n|�����3.w������}¾�����>�H`Ɉ��xKiB�ޔ<ŢC[��du��&�I�#��p�Ģ�M�(����Cy6�����G;f��g�TJ!�lu*��F������W�c�C��w���wiʗ��:֜��5W�V�2��nGƂ1Kf�~%��9}���G���<�CB�;��p�f��㈬��_���V��#$�Z[7��2;�O��Al��䩏�.p� f4(���Mn��g/Ly����R��¿��2�e�OŔ9v�SI8�����V��C@O$��Q�s���
�~�!g"���.�VkEe���B.�|`�'G>:�p-F\�������M�a+t�����	�"�*���]?.���T����i�Gf1�nd���,ts�ܽ��w:�r��[7���r�r�%�� �� � �'CXv��M�W��6��)6���+��s������z�~V����o��K ���Cث��X)4�r��A�80��7@�C�cia�>&>i�����v��)�K��c��̇m��t|Ѻ^�eN[�D�����F�<E?|'���ב�����.��u_��:	+��V/t}�	�|��`�;`vh*�l�X�U�����zz�����W� jq�2�5���R����LՏE9ͫ�j
I�@��2]]�-9���]�w ��D�	����Pt5��,n�1��\�;84��8fXf(���P������z�1o՜̢��7<ǧ×|ޣ	���~�)�u��1����D�2oC�ݰ���d/�����U�<�9F����F[�S遟4�Bp�S��>gރ�֊;*�2l?���>g���6ZQ۶)�6��w�A����8���8Q�8z��̯{�CjF�d[P�j*�gE���c֛4��",慬��HI(w2�!���-��z�C���ˋdhad+ �ABIS4�j xE�<M9�`+���}��w�w\5R[0P}6�Xÿ:�#�7&r�r�#�0���A���&�F<}?��a��dJ&��φ���F���V��M�h���BqA�$An-�7�e���#�߿yj�i�>ʅ�0K:ϙ4��K�ѻ����}ĉ�����}Lj�eN����T-Q��(}d�XݞN�:7�g� �&B&�I*���C \ىݰ�c�����	���zM��G�WXm�46�oa'�5��tz�R��U/�\,.�8a����j��Igqf_��x4�cU���?Y�c��?�#���hq�{9>��I*�Yp7�%m�G����D$�7L'�"�����>%�]���/��A����T�:���n$iI'DuE�G�xW��]�]�u�]�_��W���f�6�����9A:���=��Ea�!��W�s�:A��`uND���!h�S�HH*s�c���`R���w�]a��]ҿŇ*����)_HR����|�C��J����H݌�7�l��0gU^�2OA�I��?��XЭX
4���ʡ�8�2�����M�\���i��;��y�Օ�0y�O��wJ�Be��-�/��O�\@E2����W��ڳ��<(|�%��ޤ�'n8�����̵����}5�R�S�������%
�#<Z��y�߸l��<emt{v�� �����V�]@lɕ�_w|>�d�9CO�1~j�x���l
��uOG3�֤�5)�k1J�y��_���B�~�mԣ�3o��1�A���q����3x�`;k�ɐUҦ}^Ӕ�ـ�
1I�O�tG��5�7�u�"Ǆ����?�F�f,�7"J�x�����[ q�C���p��������U�fq?�Y�/(9r�o�d➁H?Co���yƔ�4���*�Y��
�i &�h&߯˳V�pd�����lp9�p�v	�uxk��t^��a[�iC�j]�l����w��Z��>� �qE��:��74���w��k�;8�d�'�XMP
��W����ë�Y��?U�}!�� n��w`u��4���G��3Đ/J�������n�t�n(l��W�<6�4�ѦaN�0���%��3e8L�N�:
����VP�p)�=��
S����v!i�X������4af��d�W�TR�\)j`0vF��o�,����<W�0"*B�����=�|7#����ړ�OSz+25�u9�� ?G1$"4�uQ��<����X�����=qD�h�y8c�)`R��S��&2��F��<f8��a<Մ�[��1�,��)}y.{d��B9���ּ��z� z�x����g˙�BW�
����A�C�Ⲑp���o�$�� ���0�묩zD�%�$��sS�ш�U���(���āIH���|x�V�2�{/�sr����#�vV�@/r�FQR:�Dhư"p0�0E� � ֘�
�2��dװ�Lc	%k\f	�r��+B�1��_x1�=�$_�q�AA�-�R��_���)�T8��A�XU�d@��&;��U��=!��:�F5�x0������r�y�<쌚�`Ө�RKGߥ���Y��k\�B u)@���Ai�+��|H�^	]A��>�ӡ4��B��V%��!����K��oT��O��8BE4��\�Y�I�L�z$r���V��f��54,r&{Pi����7�I��r�WH4�&�6M��n��3���K�q�^��v[�pܳQ�U�.".��6�U�-��V(���d�=��S�z�n����\Ѭ擘b�8�	��3ݟ6],Z�Qģ7���c,�����h��(m�L��W �~��S΍	VןK��2p�QL䜲�a����� U{����du�oN�~@-L��HߜZ��6�AAtrw�Իy7����l�Q_tx�
,���e�����c<��'��Ł5{+e�#E+��*��J��fv!�+��B��R|���7�e�5}��j.a]�:u`I��>����͏�n�)-�^�
���צΎ|�W�5���q�nV$��8t�w��D��̠>��D_��=�Z1�8�1`�Yο�xg� i�/��]J��,\�п6��e�����X��2�"���q0)2�f���*!f�m���0���=*k����#$<5q�Y�Wl�I��������a8ȍ;.bC?`�&��mީ�H_xƲ��j�w��@(�6���=v�V�	�/2��>g���j�v����l���S�L�#M���Z9�uf�+d�`FBd}RKq>/:D����`���Xu��rJ�T̕m�X�u�Q�Hqy��B6���bQ��x�����x9]�1am1�:�k*�l����d��Xڌ/�<ݢ᫃���^�g��pQ+#��+-�Q��9��d��4QJ,ϱ;�ɸ��n�&�U��ך�*���E������Ĵ�*BOQ.��p����N`�oZwg����/��jߛ�M�ى���#T�>���k��;'C�4񂒘�.sc	.�!f�,L�R&���u�)p /��Hd��2���"L'7jE�bĸ�ϳ����Qk�+�T�qۨ+��8^�D��m���y�$�����`���kZ0��a52�me�P[��Y���Lb���e���x�5T�I�t����]펷v��L��ZW���{o�*/j�y~3j��8a�쭬��>.�=����=��w`
~���ԋ���I_�}��)7~kU
V3�1�l�+���\�=a-����D~�_��S&��X��V͏5
<����z2��#"xD����4m�'��Ի�%F,�Jt��|8Fs��27~���E$�5��j/�����f�������_����5H�0�����8S>�ڴ����K���]�"f}������h��֤�}\2��e�э��>��T�$Kxn{�d�)���o�@�����S�ј��~�W2�	��$����jBn���Ӌdo��el�aA_�Esc7mF[�<3�}:DsB�QUS!�c�Rx^���ϳd���A�c��'��;�$x�o�F�{�����ְ ��T �*�8;m��:.|�+`cҡ���6Uܬ�k��8;t@��9	!������Jғf�)��_R���S����@���2�w�A���L�AW�H��ř�����)�%�ԍ��!O/�h���·�|��m����������	.2?N�K�^�*jI��aT$U*�M��!�N������L�w���`5�g�6�¨,�kE��'�m���06D���6��8��<��Q_�D^�}�=���9g%o�ֽS�0�>��=���/�BZ���f�g$'�zL�Z����r��%�U����T%�
wɒW����HЬ�Wl�5���4����ȥ�{Bơdu���u�93U�8m=�a��=s6�](�L�_p9%q�܆�+�l��Y�C���)Y��r�)͌�J1�$�O�8�ѐ��i*R	�1~��H�ecX���Y�N~�Z:���+�K�!��Ȟg�4�׽3 �1WU�����ؾGpv��,�zz	%�� K��+��8��Ɂ� �Y�TXY�&��� r���C��4'ӿƙ�|S'� �_���y5����#"�s~^.�p�C�,��gr
�Ԉ�k���^A��aৎ�|Н[�혓˿�����i��K)�{�n�B�B��ȅ�|P�Yn���>I�w��ٺ�}Z�]h�Lzdw���·��܎&������+�;K����$nHߪ���ůgg��W��:s��ߪ����}��H%���նh��ϩJ����r ��1��1�襯|O��G^Y�h'^VNM<�;(>ycN��
3�_���eB-�KB�Չ	k]�ӆ=���.�J ��=U2f-����9�_6c�7���T��O��!0����K�X�=�kZ�e|� K��J��ڇP��s��H�Z i:9iqi���D�����{@�*o�}	C���^Y�Fo-�ф�̱�L������V9k!��|;I:��?�Z�sɞGȌTt�jW�Zx�,����-���v����l�o+�H^�����K\��,y�qa�Şkc�����C%�`���n�-���ꈽ��2���Gt{#e�_ڞm�*9��:F����0IDp
y�(n��jpF� �!5�l'���A�e�T���b=̍)FҰ��ň;���p-}(p����m\�����mj��"�D~��m�5��v�D�h;X!K�|�F��|��!�������R���i���(A���:x��B�vGC��b�\�|�4$D��h�D�����+���	�iъn�0���{�q��o��ٛk��w������Qg��Sp%F�)���K �0%�)��r!���E��m@D����r�f�Ne���5�w�$u�����sx]DU��i2�OSSN���~�Q��C[�:ts�;�� ��/�Q��h"?tR5da���'Cc-�U����:�L���ZMP�!a��>��� j�[5a�AК���YF3��j��Y�wd�7�V�D�/�([Zy܈��"ϣe��~�2^2�ɑE����6��R�EAY{�x�i>��咝w��V�?>���g���\W�C!Cֿg�&�.�j���h��" �nkb�v���GoF7mI�QMu��Ή�|����Tf1�/�#2�`��y�$#�3���Q*SG�\���$�m?�)��6)�
x|۳��w�6&U���L�1㊤�M3~l@����j}�e������gw�lH�]z��B��0ŊcC��0�o�� $�2kU��R������%��Ћ��G��h�!��9D�J�Q+J�l�\�/�U ka�2�R��.0fR�{�L�0���;=�3�]��5@�=�KY����5��ej���<YS�߄�
^�C�g�s������iy��ÊYYL-��]L�2K�b�P7�,��R�V�T������y*5�ϓU����r��!
�U���'�����4H�Tx栱���@���´�S"PFYXi�dw����v�D�P�R����V��7Jx�@��Dp�S:ม���UEU#�^��UT����s�9�l���34��Q]h�Bm���ߊwa��/�P�b5
�ɰ~��aN7���b���HDG4wfW��4g�-��!�
F�,Y���?'K/��י��0�%>��M�nI��d��$�2��AQ��
ˁT�w����Cqw@�: ��_~�!O8�jDd����.�����XՀdZF�pc���=O)��I9u)c����f(1}[s�����⁳3�=W��=����E�Q8UT{F*�Pl���q���r=�Dr�Å��2��e����<��NkPnSJ�OM�p3۸�87��t�%j�e����Y&�JtD�ӈN�,�A +�H$�Ə�߷t
���L���9�Am\�;�#,�n�Pja|��*�(�Wt�-Ϣ��[q�@���T$�ړ�,~朙��2�j��c��d�@�@x��_�8�.k�u�d��#ϰ�ֆO+�[?�,�c��4	��4O�8�ƛ�����Z��rn�{�580�-�Z�_^�mfw+�6�ފ�k��x�������꤃�ʀ�
�-yv7M�}����-�(d9�O�T���V7�c�.x�R;�,��`7l78��e+�xM��"���E�7g�j߲W��[)��_��J^��Ǯ{��#˞{Pp�a�Y�Y����y%v���T�O��V��&��#�e H����l��SQi���|f��5�};������4^�p�k1�Q���n��s`���|0�x�	d_px@q����5ݫ�3�>��q�M�>��˻ 
 s�=I�Q�흓�i���٣��}�T�Z�Y��vO�ȑ>"+�b