��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܫk�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�gߎ[�zZ$D�H�=���3�r�-�7�Y��B
6����I?�����k�'aQ=$ X[Mo�o�����o~��P>��]p�]�9��D���M�y�~I�ʘA��l%�T=���溟q|��iN�NL��zH\M�I���u��L
�{��D 0�w��h�g�>%����2��*u��ПmX��)����/�̑蟕�H�����6[_ �oY&�,P~�
�c��~#�	�5���6VCA�F�_/�c�o�9JW�c#�Et&�.�Zv+^l��!����NB��>��92�L�'mܰ^�,���EM�5(Q�x`^L����QR��P'��Y>[�|Q1Dʪ��\8�� #�đ�aB�l�ċ��!�:�G�ѹw�v��r9�3��S3 �靘}�E���~.�k܀1���
��sv��!(�IP5�}��LC�w@F�_��h��ޥ1w"�"A����U�D����7��y����%���kGj�U/� q����c
l+�^Z�@�����`۽_O���e.v��_c|����Gd��5��R���S�	��KƤo/j�re���iG���ح�r��Bi�HC[�m�&����K�������-�Xcy�{fjI�3q���������e2�*RJյr���I~�NN��(c1�"1���;"�;	q�ky�[���z�J~}�*��&�)�ҕ)l��-;�Yci��q��e�&�|t �I���&i�$�&��������e��+&00樂��d�K�^p�,QT=A��SK�rWW��E4���o�Z>2}R�P/h?TF��M߸�������b=��l��čKܺ�����xr���mq"�$�|cp����1�	��������l���P2�X��3�E	SFE4�w��T�K �(͟�X��.d1��+o��"/�A7��L�+~�����=L��ɱ硓d�y�/z��ɻ�º ����H?<,X	�LO%Jo�\�eh�@q �����+�Xp��77���>K��u%���P��񀛚u�S�Q�u��;���\��C;>
?��D��S ��]Nι������iDJ��<[�0��h����[����X��N����ѧѡ�(6���:G�"$��93M��E�E�!g �w.{�,�0��T�����yK�t��d�@�6��`��eAT�n�Q��B�TW�b����B�=�-�edo��0������sTnI�p񈎉"�wCS3.i�����W)(�8F��Ϗ1
�	����<��{��P�݆�S�;p��Cp�uq}r���V[��W*_�B��Ϙ]^�[�����-��M^�����rq�3+�d|�G��R5���/�c��>���g4�-P�Ld9m:�d�X�%q�\9@�>`-�ܻ��ׂ9���:���20�CP+�r,Vtn�. ��;ҿ��*&Jx飱	��"�*D4B�\�P�Gv��Y�p���Ǵ�������H��q���pW1u`���E
�E�ס� pr̵�vYarR��ڈ
;a�)U	ɑ� �";�n�N�ޭَ|���~:���t��x�H��q�sK�K�|��=c��
�]ʺ�4�G�����䠕Z|���́{P�*�";��;�5�xrb
S8�!%�����O{�Ǿ�.��|�&9�~�B���	$h%K�l�s�ۉ��f��k�7�����p[(
��5��_r7#m[�}�Q������B�fc��ne{�����r�|��@$��F%�a|��6�U���>�2ėX�s�HSŁ�u�w�㪢ͲK�W�;i�جu�2t�L[��p�S3�Ht��[wO�+�c�y�R���	���)Z�ɍ�/��i��u��F:$d"H
sǑ��$�\�+�Y�5�uB��X��Z�nU���D�{9y��l�]�ҫQ8��Ѯ�3(���m
J�;�zh�2���� ~�6���͜����3����sDA�s�f��|������K����v�G͙��Q��m���"bL8��{w��a����nn�D��d��W���M�֌��t�k}��!��Z��x&d�PFT�8L����d��U�TOw�_#ao\�Eef�9a�P,�2c��A��&F��T�b8:�e2%��)Z��9�W	;���!8)n���q��d�b�ku�"!��ŵK��&a������)����@�(H{���k2sP7N��D��Y)�KL[���A���e��*T����S��J����~_�:p��("9���!�Rh��"�c��n4|�v��DE
o��|�Hg�/���h-�˦�ws+�%�{ߢ��ߴ\��Jx���͔�ST����Z��qo���ތ5�1~UH�ۈɅ/����US�@ ���i4;�Ndw78�S�^��l6���]���!�f�.&~w2��a��m��n6�(���ȓ���"ȳF����Li�c�j��+a����h�P��Je���_�
k����D�oq��1�;�j�ŭi@��CVt(ȯge�c��w�������C1�YU�4�z�߬%-�QOg#�{0���yb�@�}�ڨ޺�G-���	<��_�गqLܗ���
**�t:L侏�|��
U���ִ���]Q�Z�L�ZҀj\N�yy��"
�-d�?!֌�=���<<���}���%=�vڠ"ɉK��ʎ�h�[?48*ة�D�j2ojoN��mŨ��4V~��C����y����r� K)�*g�6��8����umE�ޑ>��(�ՖA-�XU[�H���I�tY��{M�pک�4��G�̩��u�͌@�7�(��Mh]�*
_����M�EhꜾ�'%:�
��RRc̸��w>cﺶ��Zĥ�<��Sm���?��<�F����('����	���?nW�j�0V���1�ZRXՉ^��|���:����?����Ѽ��"�9i��v��7p�O##GВ_��r/�*g��D���{���(�,��@bp�DZ���>w�ۓ$�Y� w���^��A��_�A�� &�����E�Yk��М�Y��t+ǅht�-}��BK��MI��z}77�M�$�{�u�QrU�4a`9��N��l'����3�Z \�&}��=|pXX���=(x��*w���<y����1вq;EĊj2sqEf�'Η�~\�Lm�ɘ�����q��5� �,��_y��yo
մ9ge���̱䁪nۤ�Q�z4ی+�SǏi���*9�c�y���i2:0eP����C��-g
4�����7��n����h�ŹP��~�ץq]�M,��y��#��k�H/.��C�ٝ)j��Zj�����.x򵩚�<��9��Mh� s�@_�Z�t�12��%�9Ǟ
�.\��e*~BP,��6,�d�>(����o7�}�*���, ��vՔ �y>V������/�y�8�,���q^�ӫfnym��5a�l+t9<i鷱�X���A�d�,wH��YN׃�.y"�h�䜔i���͇?"���8�eɽ�7��Y�t!�XK+��3ۘ�a�C4Gr��d�3^�*���nz��uLg� ����&g}]w+���F��k�Eq,p��;ɷ̧�Ks�Ͼ��������3�!�~Ni4dc.m�%���<3�C�H�I��[ZA �4������$>����}��|^!K��[sk��׭�6��r�$�d� ;.ȏ��6傶�2`6����7/��ggZΗ^��dPz8��b`��)��_��R�xَ]S���u��hQ��4�!PO�u] @ kA�nk9d0��n�f��{Ǯ�oZr�^T��^������G\K��ºm���hYbJ٦0�͛��ņN���8�-/5K�_�J7�g��{��88������%�AE�1�]sKZ�j�J�τ�h�V�(g��9;��&�IVi�ٟ�e��@S:�?�O�VN�ރ��_w �ߖ$'���` p��δ�F���#���.���Hy��
�5D�&���LjI� )�:ƢE�U�N�cg�m�md��Op|=��'�^��,d���m�!�G_<X�����Ls�ţ���]��p�'D
�s�_,�?�[ǰw�;���k/��Z����R��&�|$B�~��� f����nH���=Y�Ǒ�T��)��tR{�H��
-<�4�=ϰ�'$Ē��@ȱe�ʳT2?@|ӭ�)�:|(Q��/�����c����W����F����y����b�D�(�դ2:8��Λ�����b��������D��Fu�t�qq���\�zQp���<�C7�G�i{�[<Xw/�6�C�0X�Qݑ3.�>!B�Xd��s�o�R]j����`rN��m���'�%�A�R/I���7�������1YB�����;}(��Fo�u�w�B�GyVPE��Jz'5H��E��2ԻPܵ�٣X�����༳��/i����b[t�t�cŐ�jE�xx:���ħ�%�6��Q��_#�ww�E���sƻ'F<K�w
7C��.�8�V�Ǖ�1�m�vF:c��>��ޙ�$�)h��Oı��+�		���ʧV?�l�~�!����O"���o��6������bB+-qH��a�c;KW�LOXԡ2�5Kew�a��x��z����'@G�OL}����Z�T��У���0y� �j��r�ۑ-&Bf��y|���E=G�Zĳ�e��PY-7�[��<�|.
鸫0��J��,�+�\>\~���!�M�(���\��A�y]��S�J�[6�{�
�
��Ts�������A�*N5d���+GRe�t0g����Eظ�����.Xa7}��d���!����*p(�5L�4ݲ!5ۚ�=�Xb㱳�q�/���^��-���4@��i_����:��O�O@7�����8��6�IcEQd�:���<�D႐�PW$�K{�u��B]e���U�Ţ�g��螜���O�iؤ�����y�+%܄�ɏ��9��|�q��&��^��f���������r�Z[h���GQ-�6ˏ�~N훢N����q��Z[#��mfn /�Dݳ�$�TӀқ�a��d� 4�	�-�U��>\|�[��I�r�K[�Of��9jFY|��Mپ]��`l�?�[>g�uI�$�4F�V4���m�^�%��KZ%�
#uɲ�����mf1E����,p�V�
��yϽ��R"}*���̪�Ia�Bu=R:aR1���f��4LЏ�<�t�!eM�Ҝ���P)��@8�'me�/Q����M�^&� ���n�"�KV�_�>��������	.��SkG8���A�S�>�mR�W��{6]u���T6Ƈ��x��P0��'6S���J�gf!@�U������������(c�L�U�n#'��=C�9��q�j�/�X�j�@����G���8�D�1E	���«_����͛�J�O��4=D��"m7���Z~���q�՘R:� B�D\ѽ֊�~�h$�p�4x�����Еd��� ߊ3sŞF���k)�����������$"9?`�y�;Ԗ�\����>���i���5�3�V�����,!,(�I�?�����V[���b�mrf�w��r� �6U�˧�i�Z �x#ْ�5¸��p�IC�`��|;A!��0�m*���D��5mv�a{�;E՘]� �#��Fk�m������ʔWd� �L��'�#u��8� 9yoF��Z��S�"��^�3��D�RW�������#�\i��6�Cf��p�CKݭ��*���>D�֖Ek��_@pu�&j�����ٽW�w�2u�6a\��:!^�e"P9$���Xk����>���2:���I�_�l���+8`��Lp�����L�9̦Ɍ�?����T�bH"{��TS�h:!���_�_g쀷���a��g_���+��[����P�:oHBƂ.D��t��|5-�|ᥕ��Sq�{��ŉ+
F� �`�2��
G˧�?V�f�S��G=.{,�%�\�eç�3k�#��"��I���2}kV�������"����GI%��"�yE�3Mmm������	˿I�pÆ��{��9���>^�:���?�#\p���Qg�q�`&��]���Y��:��ɍ�10�.?2Ŭ�D�9�Y.�H���Z۠��|���e�ث���� �^��N��^��:��H%E��{Rw;d�y�a��ؔQ'��p�{����)p�	���a��W�X^F (̒�h�(��
�=��g"�z�A+{K1w����x�H��Gw� f������Cc������9y4���$��n�+U��/?ℵ�gR_�����&=�PZ4�z�mH���B��5v9��e�9�R:D���&@Δ#%a�5��{S{1�w�>�`n����*�nkL!��2��r�c�L�Tߠ�`dv$lδV�2��t7+������K�
����doTίȍ�kb��+�~���I��z��{������o���>��'c��5ZmGݚ���Sm�D0H�.`�Y%��P;�/1�~������0��֯.�w~V+"�~E������l��!� t�g�X��a�����w�t���R��dOf f=�f]�Ճ)�/Q�K�v��ۆ�)q�J���
4vE��(я��,��gֳ��M�h ^���Vfmq/�FD�uj�oD���L��%Ol�;4�f��[N�Z4++�X��HN\FT�BZw��8�!懰-A�/	"*��A�_^�8��|�8Zo�>՟�`���<���>	ǔ7������;��f��i�9ݣ�<�M�}vk~6�e���pA�ـn*�R��2-GTνO�����)�tq�	�	���	 ����G�� H�qt
t��9�kP9�U�<�;����5���Շ'�����D�r���Δ
jw抃�5p��J!j�'�E�ʀ)��Z{�X�0����l4Vn���_]�~����()�6���@�t`��U`hS�"�~��B�Is��ޙ9h�W�%1��,����wH�O���| 0�i~��)d%��W�HU4[+E���<�h�	@��F�Ʊ�k�z�R0;}w%��.^V<#?�ݭTE�.e?ƹR�H���>]az��� ϕ�����!���aX�׎[�� �BMf��/��\0_N4���D6�:$6�"��sr�����%��&ظ.�o��í��U|�:�J95�0��S�<.���w�w���^2���*i���_-�9֜��*��f{��@�2�^��˜⢃��$��j��,H�j�l�� ����s�gj�c��(����ܡ���;[���a"$�~F:���ˢ}�&N}2s�|<M{�m�TX}&0��x^�s�R;�n����7(�y��Z��+ꔈH� A�i�򊪟xuv���M[� rv$�޴(zK��]cn8��ⅶƼ� u��k�������;�c5ܳAF9�[��e�.	���	˺�ưLt t�P��"��K#$� ��鼢�&Y��33G=FQQaj��/I�.�U���w�	��� >���������譖��[��<CqaO��Z��{�/!��=?��w�$满���5�Р����0�F�@�2R��O��`�$�>(����z)��
jBÏb	�(#?$�N��N��G��[+i� �L��4j%��Jm��xJ���
#|+�$�Dn=̏�b�� �r����Pp�����������F��	�F�0l��{�7
>]�,4J�!5ϼ�;�T[Y�ɄS�>/�M�_Ewg�i?���J�]��
+�ZB$��%��6F�.H1[Xo=�ܬ�<\`PUQ�~���X]�o�5�	̝�E�Ic�v�mQZ�+�2���}�ߙK��d�"3G�n�'5�m��1:���1�X&^�cF��c0��[�\�.W'�F<��1]��X-�w��:9������j��Ȣ���-%DqD�߉�upu *�nQ���n �)��Y%<J_���z72�Nki/���ߚ���7��rZ��֔����X$b�D���9J<lᏚ�X�F�!�/�CݬjBch|!a������쫃�ջP�u����rg����oɬ��@�?N.�� �$�	Hv;�-�!ȶ�$@/�&�KSx5B$��i�왝Vɒap��F��y���oD���ЗW���W|S����v�y^D�����x����Vh0WEՎ���.�]O�OZܫ�N����llo]9��
�-L���f}�9�G��^x뽠��+A=��[�Q����{<�����ʍ-��,�#ל�J��
�[�Њ���^�\_���N� rG���{j�P�[9�T�8���r���~�;s&a�="ϝ;/�~��(�mH�C�>��^��1�����s�7)w��Y;�<�Vkd�@Kz���b��/�/��t���po�PIe �\�����U'2�L���W�hgx�jd�PL1�1�k�(� ��k-sނ�1�ݗqq�6�� �����:�Y��7r0�"�UjQ�VP��x�6�R�'����AU���=`�D��pۿ)�2q���%e?�Q�-u.���V�"T�L)OݭN�G��6�"·����	���q�w<����D���Q�FmQQ��?���_��拁։�C��w�(y�mc��kG�ȗz�r�]������#a�:K�u]ܭ��G���Q�?�2�~���R��%٩���U^����9g�>��^��?QQϽ�\��ߺ��'c%�!���l�ø�lv�;9��a5%N���l2WHH�C܂�k��X�G�Y���mp�����Z�0WI����jod��'��`R_/f��ʯ�����
�i�s��b�q�%K�v�W[F�}P�_�d��?�q)��`[Q*&&���	��������LX}��$��<w��϶�������%]�k�n'��p����D�4��/jr�^�jc���5�lS���EL�FY��w�Dw&���D�	��uĦ�kUM<�?>����t��f��$��{tS�Ţ�B��q��9b:�^�;�A�>�9Z)��BE�R(���7ek�V�7����r�a��j�*^P�#NOTN{j�E3�!�PI�g%m9ɏ`B4+iǹci�ˑ?Z�q���D�����	�fg�do�(¿�T����.>������ӂ���|���8r{�%Ci�㾶�n�q���3B�s��*��}����k}���U��;��7�hrQau�[G��,�ۀB=�d�<i�[3wG2��T*UO�C�t/R/���G�wC4E��_�ַ�� P�,3��͡"����-�J{��.q��@Q�^�h>��%�I�L��n����;?_Hc��m�Q������j/�|��.���`߲��,%ޚ|"M��c�Sv0M+��J���Y���zR�z��U��}y@=����/��nn�8�R�EF�e�a�=-IcvW��%F��0�,+�"!�<�9�Pj3q�k�":H��]�7dϖ�uIS��	�rU��~[��C�Z�zHWV�Ќ ��ļ��1���
�룾�VM�W �m/�mu�yЋ�?�g�Y���q�L���Xп Y�G�$H	�f����rƜ2u��C����,*�YXϮ�S.R��D�)�P_�.�s����>w{�W[޾��v�EX�z�����W�?٪g�3����,�۽m�8x��"��c/�lP-ߒ|V3�u����lX���O��:$�[���"�F6��V�����5d2��7͇�CK�t�i�;�Pز�\�u%�C��E�����:�,8�4����R�c�2}(��{��RX�K�z��Q�jI��D9�:FQ �4.-U��e�͔Z-ˋ|_��<Apv�|c�m��*���'ϙ���1�<������v�x�s�$\�#?�)YY�:��:	o*�}�>(��K����E>�����R(>N���De��Jm�9b�_�����;��ޛ���W�=A� �$�����9�6������C�Μb�Er�B%mD������Ԣ@���'�� u)�4����4��H�ft���~�`H�@E���̓v;�r�lv�4?�����+�`��"���2��]<�zt8�������j�x����<��%�*y�R�q�Lb��C���@ʒ3Tgȋu�C���j�<w�9��-��[�N��7xCu��iZNk��/���_^6j)��[g)���Y@'������E�Zp�Z��|ڍÙc������!��&&'�|Qb����+P��XS,�&�/	�!U�k2Js���9K��~Z��vX���t4_�����#fk�l�C�O�l��L�'����t"뉔�׷���\�1�������q�7�.A)�]+��sՎk���U��a�T��{Օ�w� o�o�6��D�̇,�B�+�p�h\�qCMj��%��KP����M;v��R����Zu�L42F�}:�ي��@*Ю�h$�n��"�N/}��G��;�Z�|l�R�,D\�������hJ�×�hW�9�`Q�q���� =I#7.	I��Z���l(<a)��Ƹ�W�G4~��Ò�����C�v�>8Uצ���6���X� ��!et� �Eb�s!�X��?5�P�-a��c�g����B����p��V�k��ή�QS�.�ʩzk��YOB]�*!]�Vh���8�����ǆΔ��ØX�j~��G����oόx9��Z����G�8#Φf+�����O�v��6���c�h64�%<C�/������H:Q�׶��׷�p�D)-��V
��_���M�ìHU�W��e�O�4�.t�
is�����zpܔ����agA|)4� Iw=����#X�o��˼���PC�`��x�Y��=\�]���<JȄ���B%t6�u]ͅ�%D�Vt}��gq�e���D�lv4�c�0����:���z�>m��̭P�{�_΅|���s8O��{#���6�T�s�
p�O��ϙwf�4����pD�*4��>ep�}9@x�0�_�3zC�-��mI
<O��]{ZЊ}��$B�_�r
&�����M
`N؉+���{�j����!/ʎr�������rQ�V����A�K��0ͣ�}U�:�kR�M/!%˾��-`�T����T��4�C�<�6� o<}:32W?m�v�P,��z��U?O�t�m�܇>�r���n��A�����<r��fRV�=T��8���0��6Ԧ��~��ɫ��4�����2�~��M�3w'�7(�t��p�ff���e�����nO�h�]��gS�/Ll����ZB��_�#. S7��� �ʫO��%>.�3����2�T����C�QY�+��q͋m�6t�--�fr��C�
�`bu��xͤՅ������+�o�\�RQ]�no�,u?��	N&��h�Rzh�p��^wjz��ˇԛ�B7����YWZ�>�=��])V�k���aG�CH#�p�4c�T�vGJ0��VY�U�Tr��B
A�Aw̯��,ax�O*%��� Z�*jv�ΐ�.����
������8�b���X���z��q��s�A"��l�O:�oI�,�HنU�;�M��r#,��iRQ�kͬ������4`5��TI}�d=�_��H$��=������ǼL®K���:6H�#/����{��Y/p'(��;բ�؆yzslBt<�s-%�Q�? }�C>>A��-܁IѨ�X�Nb��\��iQ����b�y�R�[Ba8-\J�0m�Q�g����&N��\�k k��6�gY&������۸�?�~ӑ��=IV됬5Iė�o���l��3��"n���2���f��
͍V�]��U�LLU]P�{�4!�2�VR�����X���S����o��E/