��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2X~�*���O���k�<Ζ�?
J��I���iR��eϴ�J�Ij�Je�V�e��JB^ �9�E�|�h,����� �������c���k�zbr���A�5b���J�f�"UP��"� ^$wW�1�t�Ў��	�/G>�ڇ�[mȺ��j���K�_���)ϕ��4�����k-�mVs/��͆Cw�$U؇�/4dY���J�=������ ��e[M����
㌞c��|?vNqs	U�{)�i5�`�s�n�,쾄O�����h~�~ i�Yrx�"2�W�y~�V�S�w�P�*Zm��W�໖����~�or��6?��R�)>;\·���jY�i�M2��6 �[�6�G��]B8z�)s���^����)k]Ϗ�E<�`;sV1{�%d�æ�b�ȴ�����r��`����n}F#c�N���%�u��e��N/������,��s�,:'W+%��.=+!N���)q��~��^Q�0�%�i�GP�9�����w�D�o�[Q<^��q�Z�1��!��1b��*�^��8�h��Č�ɽ_�aeU�,��c�����[>`d� TcG�~�F���;l�QA������'ع(��)�C�N(]�O�on_�w�<4	��(='�HyN��H�x�6�+�̴�c{ڊ��a�MOq�<��K���E"�F�r�q�z��e�{9)�A��,���'M�M^�P� Z�Ig%Z��Y���=ԕ�1��4F��T�o��rW,w��v�b�'~u�������4��I9�"��Z�/��` Մ��.�e[ǃc(��Q�-X�MwP�9m��Bb�DV?�O��m�o���Oh��;�
���'�p��5�3����W���"��G����� �^J�l6���(I3ݧd��7%���0U������������t�!ٛ�[��b�V��m%c�_�s�U*ih�R�U�,4171#�\�f�����.��i7�s[S���Cr�q��!I7D��R�X���:p��讇�l�=��O���ׁ=�rp�s����Ld���=�vi��l�äZ���6����*�H\�P�y�6�uz��H-J�Ku9r��+�a�VN̥���ؠU���]Yd��(>PG7"y0G�7�6�zd�>�q�d��:Bw�'���ﶅi��#��+*��>�1�A63'qdv���2� �����TR��X�x<h�����p.Q"O����G��+Πke&������{��eVÅ���U�j'6����Iݨ���#�T������)A��QھX)���y�=R�У!@��+WV�4�7�4����[�LD1>��Q�C�w� �8��Bf�T��5��xi��mC�J�YFa�F��˓o�x�}�ɤ*� eaJ��>��>��7O�Ƙ�?G�j��'��u�S��D\���:������s�!m�L�x�|,���
b�[YwԀO�`S?��|{�	�@O�E�䍖��kǷ/����ra��R���j-��}����?̉�}}@� X
Ȟ�����D:�o7W���+/
\�Ӭh��6�ec�dh��,@H���ȯC{��.��~�xj�`���(&��In���ܦ�Ÿa��jS���*��'��8�?�(����@Ժ.���ڣ��2�ܺ�?�w�-i������2TG��ժ"F��B͎VOM�����K���Ub�E�?~�MD�/rԹ_��dgq����O��O�������6Nb�>��ª����<���+�)�!x(����
8�����	�M�)�\����h�ENϨ�\)����e����h��T_�x�M!�7mB�j��j:���=�&M(��Va�\vA�Aq�e�C�!=J��i�l��>��m�əJW�S5i��Ǘ�0��m?�#N~Đ�G�`��i�5G++���@k��Kk��'� ����`��������M����\��b�Ǩ�Qqf������z=��j��vz�]�/�S!�X��Ev�����]��,���N���V�h�
>/���;A�!�-��X�k�Qg�ce��H@�0����VS|Y��eX:G�s�)�µ#���`�IHQTQ��Ԝ�F��G)��[���МVƠlw`ٍ�H����uk��am�;��q���ᾮ�,�b�R���r�b�V��w�T%@��4W	]G�&�2ZukX����U����0�x� �3��.p����Q�%
��)��ҲC�P��*�^�Ļ�v��%\���|���c-������#u��!�����݋��I����m������|yU��d�a64�~PReL�j6zr�#�|�0V�1&�����z̹�����Q0�43�=�=�P�ܢY���`b!�!եjE!��0�8�Dћ��P���P,�����qR���J������d��z��(x������2�6�xzC��.�zt�-g?��W��ض'e����S�������Z�<��~e������Fb�q�Y�Cc�-������N�̲�ߒ���s�ə�i�m��	R0+J���ģ�	��� ^�I���uj�-v$���9�4��X�9��+
zXA8�o���W0\⫌f5��~�p�%�X7$�R�	.�t�`�J�����Wy=g�	��V���;��&��b�D>|�js ����a�֩�Q]#]�F�7��C�!���ꚥ���N���9��ڀ��8���(bFdM�(b�m��<��pn$��v6\T�
>�-ƾ�?�S�(k�Ek��+�O�(�����"��`�DU�66j�H���ӦZc�Br��wv9��_<^ ��X�M"=���0��?�!Jm�t�aYU����_|��qQ�QbS�R��˄\�� P"��X�WQ�˥YQC,0��I1������!�
Nُ�h+}  .�ӈ�E���\�'�n��I�E�p�$�W�
����1[�k}�h���A,��H���Εzsf]���g��&� ��У�L��Q:eR��	p�/:)?�N�u�L�����)��̜@�O��\~���/�!��?mZ�J���|�z�h�����,��J3=</�a��6���l�Fu���Z2]w!D�m&�?"��6���l��00�*�Q��^��o��+Iܛ}.t�e:D���+��7�bzj1���qTs�0���.��i=�(>�r7��;�k2��<Q��U@�q����卼,`�u���K�qB<�M�1}�����M��gh|_���T���ά>4��G/�l��}��įW<�@K�n5�hs�W�[0����������䨖�ɩ]%Af#b��(X�ᖆ��lH9\��V���r=���kj>�j���V����.[{�y�Q������o@O��֫W��̃���7��A+G��=�n�7^��ş�Z,PT�SI5�lJ�K�^�f��c�]�*�B��ݟ�Q��htguf�ZT�Ż�� �>���8YX��y��F�}M0�,��4�`�_�=�ўJr>Lm�Q�0�a���n��@ɀO׭scI
��gs"*�<x�qqyGZʢ�qQ���~�	�EڪǙ�ލT	3�ũ�&�W�g��Q�E�ɕ �_iP�Sck%��rD�U�W	o,M�Y��o��'<s@8'�y5Q�P��>%���4�۵ x����#PD�-�sk��^RR�U�!I����A|u�����Sk�V6XȪ���?�X/���>��ſ��ނ��m1��A�mUyr2�}g.r:|X�!5������8�p7��9I��i_�
C�n-������H���U(���T*v!2����GۣLܕk��	Ȁ_����J�h��W��0�@ 7|}�iAD�.�
���͸#z����aN�d�Ux���n��S�K\���߷�`��*R��<���B�����p�9��I[I����Rkݍ_���PNY�&-�l~�ⴖ���1�8
O� _�-ΏΌ�T&�ސ[lQ����H��[~T\�Jy/G2\<�����ņ���9c�8w�����2�wR�U�����A�2	��n�,P���0{ŷ�wᶇ"D� ���D��4���9�P���������j�'��m=o���\l��r��WSL���^g���ǧMo���G`%���W;�]�R���D�z�(��zm.T,��
TrW��l<�s�P.�DAG��A^J��SA�#��W�Ȕ>��rnp�:^a
��a�d�}��7�&�t��9,�vQgNqz�1H�nm�	��U��9���4���)Rni��u���+����b�e���^|,PI�OhN�"d��A�Uks�yI���\ E���Y&'��2��S�n��꠭{�V%�u$S\s�ly#�~;�OnoO�!e�B�A�Hh��碣<5-[��B�8�
H5o�)Пc�{��N{�����*��g�n�Z�S�f���C �s�y��=%�a���Ȃ� ��*��^��
H����J]R�sT� 7���}�-��a�̮㼊l6��f�f�$��0�9Kr�K�}��t�{�YZ�Iڊ$G(��aGS�ߒM<9l�����(|\@I�q���LH��Vt.�#��-l/��h7DAW�ܴʽ ��!�%�;�0���{��V��������ߎBu�,������PX�e?�x����~@����ޞ^`S`���ge�,O�Ϥ�K	�@�z���J�&*����u�m���U�����N��C����K"|(~�̑���KM�{��X9��g�jݨ��<�?�iV�	*�I��J$LyMV��@���6�o"�I�>D�������-�Ӳ���x����!�'2�4�[H�#ɾ6�:	�+&"L��!_�.~�of����5E�{�쳙��W��T�R����)��l�_/�T�w���8��>�t~�i��`0��گ�ok��48`�E���\��'��t�=�3����x<��12�P#a�d^p�!1`���'W	���uE���!7%�S��*�j�p�T˨�ݳ��P��U+��&JԬ���j��zW��֕���U�V��˱CMܗ�6	!/����J֣Z���Ro����p�9w���Vx�߭./��$���5�ΤQ�_r`R�����n�D��!K��&��-�� ��@F��U4_���V�����[3 �D�8V��#��&D�%֚��#�X�$�Ѱj��<�3�+]Ֆ���0����ۯ�oԗ2������)��_�%�\f>͏.d�18�ܥ�4f�2�� �*ֿG�,�#;K팫e���N���Yy��k����_d� :���JDm�\|����%��(m�B/���-����~Y�ཀ=Y���QF�D������]4}��f��R�SLg0�E�}J2�'Ϙh����Ҕ4y��p�<#Q��ǹ��N�@ |jV��##�m�G�����.	�G)��H��6�u{��*���*��I����g#�i����P���S�A_���,�2%�x+v��C��i�֓�
xh�ˍ�4���a�8�L}8����l����v���Ap1��cz���w��R?���?�Uf��:�������l�Ԅ�QB�nV������;��P]���z"By�G���1�wL�)� 9�u����<婖
Ώ_�|�ዘ)K�
� d�u/�D>��յ"O�o���s?N� )��zr�rGw�v��lH��';����!�aC���¯D�Ӑ�soŗMF��V��Ұ�vt@�r85��Fs:��qNm�=���"/���N_RM�xH#-�Xxx�'XH�\X�A���b��؜��q�g���t���}M��
L���y�J_�H����"��s藕8�����MK��ִ���c��6<�S �2s�N���X���f_R�ԧ�b�԰=��sdnق�+	^��'�]Cx�Ǻqc�F$kqS^��3������qg�VH��ڻI��`��fg��/u̝�`��\��!�+�$��x���nŘ�4Q�՗���p��A(Q����]=�z|#��ʼ�z����E���k��Q�ND�Ӹi�䲧����J��!�������k����ÌD(�H���3�E���/��	�$��?�}�c>�(�A����I�fq�$`MQ�@��?�6'��{d�ʎ����3��C'�t�RǦ!>�aM����%O1�/4��|N:F�ʨ�3Vx�!�7�9U�y#v<��pϳÃ)$���ч�aV��"��u9�R_φ�5񫚕�)�C�̇�Re����f僺�({���m�Ƞ�����3��9L�+�����/
k�|�]��Yf����(�,� ���T�$�!���N�d��hc�����̲g4�-,k�q2>d���\8�u��:xσ��|lŇ#�`	B����GL�>5z�+�٪	�cD[PK���s����0���G�2�pFw��]e�����?:\M=�{<�:��`a�PZ4���+Z5�_k�ч�X$��!�{�k����X�����t@���.Z�D��U�v1�"C���kNJ�S���!��2�*�o�ΉDQ���%�dӯ�J(�;�v�'��k�E¾w���7ɍs��W��AE��}��=��JRu��ٛ����V��b�m��e
N���J,�eZ4f�x�����i�f��Ϩ���ڀ3;�����tq��K0���K��Θ��&�
�e,ύ\r������Y̲#�k�l�8�6���7�7�s�wdW��f/�7�p�?z6�U֧E�OV����亭�%��!��'#��l��z���(�gj�Bo�����-.ZA�&E���ݫ|��|��q::&6�Vɳ�Ӟ�Ϡ%~?�'�}ae�����E�@�X}G; 8���l��c��P��{�e�~fA�LA��w�.(i�$%����l��T��|�9}��"3���Q����|���c"��~�G���Og���	�[E;�}]���퟈7�c��nbl~�����p(z�	�!x{�W���"D�=Fl�ť���h���^e�����V�|Ǯ%fえW.az�On�Xo1CW��$=9AM�9K73K���{w��-�ޱ���(�#���x���U�gV^5�`r$j�v|����p��!�*���׮�A��(,Bfl�=��Wqn�9� `������USM�קKM.� ,��E0Z~n���T=#�<mK/:ْ��p~j�|
DΫ�(��r��H ���>�:�5��C�B�;�G��U&��
��F;ai"�S+�� 0��}9����������y���Z�eO��O:�%kD(��\�FC*�:��7����_i3����F��^�D�����c$t�v\��Ҏ&�aа9�W��)��NQ��>@"�����+~'�h皢�Ҽ��pA<�����o��-]R���ۖ6�>��0���؈8ʹ�Ib��/�tj:f���������m(<k��1k[Kb.���აfa�*w~��C���K�88�ȩCTO<�����F�]|����F���5����J��v�3V�x�'1��v���h��f�y ���y����<j_���A��L.3���n��qԛ�Qh�w�$�)�p����O�^$n��)^�Z:ϑ�A�9��eI��I1n<��B��p����6E�$_<�$�'�4.9��}?�+ߢLWQn�ذ�<�O���i���s��⇇�C%BA�3_�����$ͦ�b� ��'[��p�}!/7p��4V'���t���5"��+�d��g�<�H�U�K��0-�rf�`�P�a�	��*M� ��:xd���j����Q���}�[��,O�b=��������.�g��'^����z�p��uD�l��I5���:;�T[B�&���+����P�Y�O�_s�z�8�4��n�(r��l��#$_��>#rs�_�v���r;C��a]�P��a<gq���~ŭ�_O�>U�fEH��d-��O��U 	m�H��K7�4������]Ѫ쿥u�,���da�/k�� X^�����̻��u���Q���D���p�g���ޝӱ�*�m
�s�mXZ[V��t��-3��J� �G���c�9�9Tӯ�M�k8 *=�����Dײ�ejT����k,oA:b-�v�����7�{����
FE1m�ʭ��">��n>�k5^���^�����_����f���"Q�W֏s�r�����/��%虴l[��q1�q,ښ�V|�\�F>�W����~#s)�t�-5�f��S����F��}zp��m��&~��Zz4�޵|��'��^�̔�����L1t�^ ���3F����o����{jxWم�vp[��qQf/�t7?t�q"~i*Ƽ�ٶ:����/�ᯖbd-p�q<	�X0�s�*Ma �Yr<@���H�0� �F-���lc�R���v/��P�{��鐊O], ?'s���L��婧�Bǔ�s �)�&���q�Tr>$���j�����RZ�L�1�^Y���$���ਆ���?"��`塅ܬ%q����tQ?%`��ɕ�6�z�mYA2瘥����:����K��,ewwg+%����l?s��9�Eq|*�h��*z�ii�@��GgMYy���bN��Q_�$f"�)^[Y]B����E
by�>*�W	WbO:A�_�(�-�ѡ��ޘp<�Ihjt��d�� ���}b�lvJB,����U��-������t�	wM�05�~�Q��&�n�f��S�h���T�m���c�:�OA�$��N!鯯w	���MA��q�����.$��j��y^�
�Y�au�5e��b�Ӗ&4�B�gC]~i��_�<m&��֒r�����~��G����+��F���;�7�Z	bLת2�K�'�P�1#�};?ߤ��O��Κ�_��ޤ3!��w���̶@�Nǒ�!{s��C�b������"+�`��x�u���kf��w�:j��!��>�*-��|��^��̏��z�0l�i�
�B�AJ<�e�H�ow�����@'�Y�����Q�7�+�kv�=/_��6�+�������_$;cf0�D����	p�3^;M� 4{���-��5�7�Th�~������ճ��:#=�4X��[,�r\L�����No˺�G�*�#���è��Z��Y[?U�%�~��6��m9k)j_6:{��i�P	E˳��_\$�ݨ� 9����b6#����M��LW[��m��� �j��$�KA��H�����oLIm<鄅+P)�V����e��Ag�� iC��g%�:P�DђR�3��C�#'Rⴢ��0y
ȵ��@�Ĩ��������r��b9P�i?R5��I�QF�>#ge���zy�>+��Ԁ\ _%��?���x҄�
�zYU�4-|���3B�B�cB^����&�m*��>��w/'�Le9�����gn� ǐ:��*�VHv�(MPe����94eh<���hoV�1���U�ʥ5V�"��Х�=v�yb��Ć�����'u��r	��i�5Q֙"*����x�5ƿ�`YtƟ��m%f0�	������Є3�;�s�<4tM!��%ŉ=��y���i,�$�LW���wVv4��y1�aELJ�l��$�A�5����]��}q���!��{�;�����wr��ȘVx�x�t�jM����]O865��ΓQ�E0�xH2�uSfMv�/8�+dA����o�o��/�>�<FFy�ϜE�А�X�ڽ���GCouS�؍<P�2���1�0DY=��˩��4�U~ů|��[��M1|]����ɻ��E�>�-Od���I�8�o5n���a[���N@;�#��NA�M�5��?(�!g�`�G� ��$� 8]�/�r���)*���6 �[G���Y}ٹ���n���R����W[F|ot|%�� o��o��TT�pq�{���4�4�7q�V�(;��o�E����|�ٛL���f�K�y@��{ճ�t�GC����@�����ɺ�؛3�0���Sa��b]�Բ��TǨ�o������0`����6g@�&i�5{�����WI���K���h9�ȷ�,�-��_��*G�s�����6�/�Ǟv����[,9c����2��:qs����ә���*���>}�������: F]�(A��L��"���� ��3w�y3�l�d��&B�z���������@2��I�.�7���nߐ�'\��?���Q�#3��[O��v0*�^u�s�<��;�5�$#8�����2-������ڸQ�/�"���v-��*�^�?����*�oϯq
 XF}�
��7J�O�_R���ܑ}��y.��y4��)	p#�9̍��
��A�3�����o�Q(�
qW�`��W݃PwU,}�t��]�z��Z����6}�y��g����aIx��{�A�t\+6���n=J��P=��(����ʙ���� �EGv!�0:��L���=�Li���g������Tr�%9'D��Q*~%H�����������dSq��$���e4/��;��}ڂ7�쐈�f�tw�� ����U��S^�F�5�';:�6�9|OI�F��qSI%��jʀ1~�v&(� ��p[�	�g� �q7�)}/�L	��'�|oH���O݅�ụ,Q��jf՞\�E��QRE���DIIV���e�?�#�9}�c!&70,B:Ɠ.#���*W�̆c33�r�.�(��Jٗ���\����Z6����X��pU'��j�������A��X��&|�S���>VafB2�Frw�y�0��������w��|�$"�|G����� �dE=��<�U��|
zج��l�s?V�;f���ƨ~��ë���g���'ղ�A�����.�)�RLa�I|�x��Ŕ��vFީ����1 (X�t��mMy�D�*�؛�@�@6A[	����00�7M��6)��9����}�L��4�������	�Z�R���;a�[���:���۠{C6�3mr����&��7�<D�_��9@�+�����I��%�g����C�wC�.�}�ۡf�	O�����o�TC� L�Dp�[Vȱy
C����	 ��L���ǂ�#jH�)�qof#�-�O���>Hּ�X��a�����f����EZ�!����L�.��ⱉ��5~7�t���?�k8����ƚ��p��&�*E�n��c����F2��yL�3�9I��97����:p��Qm��=��+��X����2L8��5P���XEHd���=���OLplqM�WM����z)��_+�޸b�ic6��?2�C�H�Sw�	r�\�~N�i�]5���s�ӘM��j��(�~����S����D~ơ��Н��+ qq�<����㆟���ct�sH	�?3{�w�ٿ5�%K��#��|?�3AЊ�zfA빇>��F_��$`}"�G��)|��\p��¦�/צ�ԗ�+f�F}Q�G(����wL)�A��b�p�u��A����7�p	��1���dc\��{v��F'��d�bi��"��Utp{�[Z�<�=>�Z��8��ǒt��!�N��9��M\�m�F��Y��=)U�O(�T`�� ���8��
���_M��A�Ͷ߄<d�j3���Ł�xRI��ֻL��Ϣr�$�:͛
�d�jY�M�(N~o4`n�VÇ�'��G�"�G�G��Vh����.p����	$[5��#�{�<b��j����I%m{| U>F��}�Z��dA�~uv��C�Ypcu�F��];Q�0���X��s�jC	��0[�u�/z�Vڿ?�I�2=eMF1�^�$�?�
�}'��7A��Ε�p�%;
���������8�E�[/����m^3Ύ8��LD���s�B������$~�+��A8�L5�u� ��h��]&آ"h����`�U��[���l�e�6�����/��}ȋ��E�D����Β�� %
⃽�.�1m�����u��c�*��i�5���C����D6ٰQ'/>�E;�*vZhŭ���¼e�5\~�ƋU(Ot���.E�Ϟ'���k��N�JOT�O%o����i�<�|X�����:)ޮ� m>U�l��#����.�\�߮*�E����X$�����,������O�����������5B�A'�7��p���&f����)�8��V��֧�Ղ;�
�6��}YzH�+'����Xgn��BٽJ̦�ga��$0�m�mEݗP��Y��d�{ �m&���	�������̯dT;�Z��ݛ�A�U*�W�h�'�V{ ,M�\_��PJwݣ%t)��m��Ņ���	���)����p����c3[�+�$q��m��t}�k�A����:Z>��o�B��9 #&GnX�f�pmd�t��������&<�V������) 3	(�� ������O�ۧ�Y�,�U��H''��p��1���'����`�*�N�����Vf�4��N�n�P����D��I ��x�g��W��!|�2#�*7$�"�9��6�5��q2Ak��]�l�9��*yT��� ��4�C��, 9R4�S���HW��[f�s��iC8lxkY/����x`�Hl�P�-?����C�a��Ц{M�\����
�Y����}��1QS�m>K�!xU�lL�)p(���f��+�a�VE�p;����`:0�/��`�<'���C���#|*�,�+|ᗟ�D��9���,��lrl��9ۚ�	*` ��;,��><T]״�E���t�������d�r��������s�!�	~зefN�92A֢�2#u6��&�m�>l�T,��8B?���$��a[ܝ�� �iZ�x�w�#?&⻱�X�T?ᎀ6顮���X�'�v5jn�e����B�I��k���5���
	�Bl4�W�騼����i%��A�\5�r�y�x�}Ǳ��&6��蔓�O/�V�]�N�R�o]Ƴ^���+�UVn��K�d��iV�b���g�R0�V<ł�e����̬p�+��$v���ǥ�vM����T1 �oڦ0.�BG��Nm3��Wi���>Wl>Cd��漗B��^�S�s�X�-Y�h�#Wٍ�S$��,�!��@�ꅳ�=�Wwq>�\Y0��!}DK�I�@�\
"����m��e�u���s�L��]-���W�+�{Q\��K�?��Z1���8P@�~�^#=4\�� ?�`�{nS��3W60."W�����{M�xXj#[N�Stc��R�2���F.���ܝd��q�)5���Q�s!ZF]����R"��\�
���%g�g3�eFJ�-Ȫɼ;T<d�vp�Κ�~��io�[���f�A+�[R��8��y�2���fw�B��+��֕���&q�t��Ǩ�����<�F���zFԚ�eP�����!d=�4�� Cj9A

c������oP���Mf0�A��Lw+��=_(�pe��S����s�K�Y$�:�B%�*��7��=U��s���H\-��!�c��?�]�. �W��L��s��U3�dS? m@k�&^�O�AI,CJ� �{Md�~$�)%4�u�0���un+,� ̖x8Hp���1�m�q�6�QR� iv������g�zO�@2�vs�w���)N�hx���<՜��]�c]�eVM�&YE�i9iD��:$�x@���W\�=�b�*�>����j	�d��b�駿�Z�q�����	��C���%ꓮ숗-����:��sg;�ǋ�x#��KhW-4��
{���
��p�e��_�S��b�}֊@j��ʔ���r�_X*�#�$�?��ڸ&q���o����,,Wp��+:�}��v�l����c2ؾpA����_�Ϙ�����GU�79Fpi�I�a[Hk;���ȍ�Ư|���X��i}����	j�Ջ��B܇)'����EV��i�ꭤg��� �
>>�������W���Y�e3g@�0�0�qH�{���Z�d!ʌcĜ�w����d��1L9w;�n8{�~:���Û���˞���4�X8&�G$(�z��O�P � a��^��#RN6e?��˗S<-��OK+�=�I�{jD��~��l8ဲ�CCk���$iڳ��&Sڦ�gR�T���gƽb�M�q��g�`�O�N��>�O&�4�S��oڥ��ݲ�H�؂�S�x�M� ��ߣ�y��2k������;�;M����ac�Z�)���Œ�S̭uO��|�c�g�Z�7z�����
T,�o_���-.�L�*ZK#|Y��g�-e���A�Dj��YZQV���� E�/����]��*����b]Cڵhbs8F��IҮ��=R ���v	��iף���ES��媪�g?���/�邍,$ќ���BO�%���H���9�3t��)�B����`�[Ͽv+��߁���������BSlWr'��C�0�*���-���V>Y�g�C7�	�;��%z��,M�7�^�i���OB��Y�5�P`m�4���,e���$�<+BB�$����B�[��_�$��6ӥb�B ��U/�1ȉB���e�l҄.8�Ņ��qIh_D��*z���R�,de���!��#�i;#"Rŧa�> ��R�`�1�ܦ��'r��p8���㊮}��@h%䏛Q�=G!	a�ء)����T��9�5Ic'}�_�i�ʨF�&!�ǲ�ZK��K��o��5��B�1[[���yR��v���ڧY涼��8�������+���J�uD/�uBԬ� �0��:�2�"�M��l��NNOld��U��Q�s_�Ԑ��fao�g�<>!�Aj����)\���A�����Z$Q09Jн�EXhi��/��%�.�l���n�`:柤�����nYL�J�ؚ$��p���6�7o�*`���Sp�G��^M9ɂ�L_7��ʕE��f�o��:b�[b^3�&���(y4���6P�*��/�q��a�&���m�1,���	���:i�ފ!�3�Pg$�Y�_9�j@~��ue��
L�3K��|W=0)��فY`#|tL߸�[���M�Q���O��6W�[[#"�!�s�e�f�+dc��V�{��n�����q�-��;�)>�<�0�c�����=^���}v������`���w��������'�?�R�j%��Kp���2$��`b�^�"�a��#ď��Q	�3�[��ռ����pEv:t ��R��}�rЯ34������ʋ�NI��iV"G�Tx{Z����Z�6���0�%�8���x�y�z�Wʼ��
�J��ic�$՛���)���>&"��6��9�o����u��9��Ow�$v6���i.s�
�mC�!�ݼ-~m �+	�~իɝ�ڜlO�p��ՕH׷Z��,����>�v���3��� u>S<�F���Tm��w;^�r�Â֥�i=!�<r�X�"�&'�a�ⱚ�ifM3bZc��x#�B&�I@�'� ۸��dza���F���nH<j�l7N�x}�6�Ijդ��NnM�s��b ��n�wc?��]���Ŕ����A��	q��3���)L&�lš�E�&��8�V�&�| �fN�Lݏ\K����ZZ���Y�f��ִ����P�'+�Ʈt��F$p:n����w2ǫAuGA���XhPWK��Kv��&j��O���r���a�+�!4��Dn{#1��!�f,
�F6�v�D�I,�ķK�� �T��N@�恹��zQ�J<����ܵ��:��~��JT�s��˽�>ٰ��D�=O��z�h�I�=�&����p<|�O`�y�v��l�*���i��c�\�Z����+r<Fh�D���a��q��VТ��̆n�/KbeP�z�hh�_Z� ��x**=���b#�E����k�� �9$��/���Sȹ�xg.E��,�1�B��k�gh��&N�����E�(SH���$�}t}f(��,����~�(}1�/82/��W��s�0�dqM�X;�D���gc��mf�� B����ݰJ
j�0H�ߛ%(�a��[O3,��hT���'�s�ޣ�ߑ���I58�òć3�|}�^�1�L������,?z��d�,*lx�QC�E�nń�'�_陷�L��b�yv��o[��Nr�|�U�ܲ���)��_)�޷�`B�ba����	4?CZ�b��!�#7C�
4(!)���1����[R���"�0�Wx��o�wQq�����n��>MS��	0_��U���ѯ����y|ӛ�|���3��w@T�o}����n-�6��T�oag��c�\��5u���"����}��CQ��գ^}���� �7����܀����,	���[)��3*�,���BdG]`W���I�]y*�c5bթ'��\���͚��<Sx"s> M2[G(�~�̇�;�\}��H�����r 0��J�&��R�@KF�0����=]:��E�E�u� ����{o��n�i�ظ��X������_�Q�"D���*{lyB�.AG ����Լ�y��g 	Q���c�H��q1����~���-�������Q��d�qC\h�8����F�$ ��G�
݊�X����<�G7F�QZx7l�%̽�?BZ� !4q��{yvxA�տ��Y��jn	���c�B~-vm��*U>�kקQ�3�:%�q�ID�?��u�lHF�N�hIQ�e�#���j���+6�+�4#�T3\N��#�&96�p�D��d�y�lG��ID��oXQ۾�;�}N�	ZZ��;w��m0�	{�:xPZ,_��=f���r��l�l���]H��kg}YҬ(A��1��)�z�Z.��������^_z��������H`��S!q�V>�m�(/ʺaJr�=�.h��ڌ�ƪY�x����!x��8[�ƒ|�Z��<���� f���Q�,|�����Kvn��@�`�m5�QX��A�05̍��p	N$R�nϪ7��O~��Y�X�w�6yoo��G��s��R��M�ˡ�U�3�0(�@�bE�Z�K�/������:���I�-{ˆa$�v/��cJp�Oex�W�������m�q���q��f�>��d!X��q�1��c_͞P�A�7T��1���ےAz.z�+�^	���722i���mKIL��4��UM�B�k�Y�����ӓ�Aq���H�!+e9��Ϯ�:�D�s��`O�).A�m���L�1./oFD�ybR�t���}�p�t5(M��P]���&�ov�Cu~�1&s���{���\@#J�'W�%+�҂ۤ�jM��D����� �#�E���2�[�T H+��M�mV�%��t���R*m�X���`�-�Zl���f��wG�r�ȵΔۂ؀oHP^�?ղF&��\������3u��X�=���+���M�=�Ъ��������8R�PR���h���1c��3�G"H|!-=G�cJ0Z��xfJ���մ�Bv�蔱�Eي|[(B��e;O<B�@��3��A+�X���${K�e�)��(�0��������ѵ�L���# /�kF��T�VG6�F����3�f��/sckd��d�ϒ�NF�2�~�ک���h�����5P��;�N�R쾃���/6���U���\�%4m	8�B�Rni~a����bUF괲�c���-Ҋӎ�6�j���5{!�g�ͯX?/��"Q&�>��"eF��2[z*���\��ZG�Y�����{�xI�k��b�!d�yD�!*!��9N:f��Lx����{.����e�;}��Y&�J�3�>3��D$�����"� KxAb1
'kb{|�0�Li�ut|"	�n�RT5/���,{+s����ν
I��)�CR޿�0XC�tTb��'�i��c�š����&�O����L�?T�,��θ�K4�.��?�{߰��!��$�."�#oJ:��c�z�Y�q�Er�����m6�:��#�^�����{*��tK���M����N-��ݐ�}��i%��Ymhi���K[��w�ذkn�r���%#��WQ���!�J5P�\[�E��.�~�4�4�����Ҍ��]g���N�B Y��J\}}����6�=��N|��M�S�k��?M�F}m*�gx�O+��j�*�͋�e���D�� aʜ�.\?u'��f�n�b;��m��S�Nd�ℂ���7�#C7q�����@����G�i��R����N7�b������Ç�����E��c�fS4�?T�e���^��c@��;�W��|<۠;mh���d��ɮ�>��A����;
�m�ck߽�wR��W6�qKM�I��-��X܃a�g���JW�h�j��z����(�Fɘ�^ե�[uM����`h0�6���t�1Ӷ���j�۠�_P �)�]�P�D3�M�;'����H��Y�Af�С�[��Xhg���np[v,��\0��ߓ�u�a�-�l9#��j�6�H,���l�?��ec͓�K�K}7"-�r*|je�O���TMGx�=$o�j��3�h?-����gw��B2 �:����uWe�4���f�\����_��Z���[�P>sǖ�$v}�$>�b:f=�d�G��"�̹#A�wn1�1��(Q��$�N�/����� �>o-�ff�9|y.
?��#�[y=���q5�U���{�JUo���-ؔ��ը�#�R�\i��,4^��D6����7���:Z��(�J�C�g�U�4+�!�&�u|Ee�j\��8A�	R����?9T,�����'*y�׋ #gHe��սas�

��@Nux���sW2�<g�_`)_V�t�Qe������6����W$���;ErY��	c;;g��)U�:�6�V)��$<�67�v""��e�(�U���V/�ܙ��}2_D�(J���tl9����va�}q�TW���[�DX����c Ø�U9��N�t�\���@�o����ݔ����`^=�6���.�����zoj�[z�h������ROJ����4�V��xR�|"����uo�a�P��Ѳx#�1?u2Y̵�$�>������k8К�^w�|�����!IE6wS��2o�Ў���ȳ�c�VM+���g�*)qy~�ߚ5�h��OBԉ���H�'���N����oYs��^��I����rxD/�i���J/q�#��[6�m)��}��S������z<v?�G����-�6����ۡ>k��řb�jb?�U���I�]���"I��˺��㠌��,E�R[�>C.�f\�p��?B�&��Խ��M���|����{
xf �6��&LdNeNw_�Q8g��눥p.�Eo(#d��H�5��ݸWk,+)��D���爄�wԋa#>��0r�A܇�WB��=KLɔ�;��a�gyL��{y��b?��I2�s_�Ώ,�Fh���n텡�r"E�u��e�pdC{��a�ƚ<���C�y�7h�*(TyJ���kZ�Z�Tڽ-$�ȧ{��ۋU��°��t�RE)�:.�Uj_\�]z<�Xq>��é����mѬ�gD��/�� �����>~���.\l�K!���[C���Ͷ�"�ۣWMV�JƺMe-59S��f�S�h��tC����v�?ό5��x��҇؁��r7#���U|vyy�]����m��=kM�=����)r�n���LΎ�	e	��<����^��)�1�Q��w:%�'��c�%USC�qv)|n�	�K5^j��x
��;�}A�`���.�����Ꚋ���<�u���F��[L�թ3�"��0��+0��Bω>�H5FҷIj���]�d������}�����Yr"���>Aߺ�/�8����C���+��c<��6��3��S��),�ĒǕ2+���^���r��*�=�PƤ=�1F����>�m��vV?���� ],��=V뇊V;��w-lfFv2e�N�k��iHe:*��f1ӓ�WEP���"���^-|�~׋������b���$�p�`��G��bk}[�9\LJ7��)w���d_��x����e�Ųt-G�4�����^����=��N|�H��(�zXy�2@U+B>�ӸV��������ɹ����|�x.�߮juo8]\sA^)���M��9���6(����dG@$I��l�� ���� �_�\_�'�0�bB?mA5v!i �*6��%B?RU��"?�ms�RX��W���,�4�Z/��z����İ�̂�`^|��K��/��i�2b-?P��4U�m������/eZ�H���dY��D���E�]�x�6.�iYJM�8-`=�;{1E,$���K��4�Zr���.�e߈��s�ne�:pf<��W��bѿX!՛}%*4�B���A!��p��oӗ��"��4ʖO�b�k��MZ%bS�ko��<��%��t�4(b���&,�'8�;�k_vjV~�Y�ܼ�yjպ9]$�Sp���\Ԍ���>wX3j*�4�,b���|��3������ j�\߮|�X(��jhB$L��I�nq>�L����r�$�b�Yr
��5���S;�K��o�*�m���� g�G�ak4�G[��%�}�ib{���ߣ��T&���ED��D���<��AP����R�O�����m3<��>�?�C�@Y{��Z����v�3�$Ї���P�#y���D�xfq�Y1�HH�즨Of���Z�@��Ӟ�n��\�L-? �3K��HArcHe�5�{{�o΁�23�mW��	ѷ�u��[�͚?i>x�w����)��ܽr"[+��	����5�c�� �T���X�
����䖓�!�$������\�[E�A�sAJ� R�k<�0(�0���ݞFHkgV�ok���>��dA��B���F>ڈF����!���@Ӕ�A��0��B���5���Ƭ�W?��׫L�hˊ� bAeh�ɡ�����^���鱨3%��6x(�j�9���f����A��іsߓڍ����V߆p�c+<�w�������B�t��H�O1��}OV+�J70V�;�hW=��z��++S��g�Cd��T������Q�|�1N^	ͱ�#��e��<��l�4���Q`I��*p�$�������o@_SC�i��&��&��$b�/`���&M]�)Z:����:���4K�(�0�&�M��K���ƑC��6gr*ּ,݆Օ��:�<���ɱ��EQ�c9�'���CR���f�ܦ ���0mhf�*q�e�7��h����2�kz�tǣ�{����P��s�ߦ*eޘB�f��$�����������d�"AE�3���N����_�mK�øΦ ����2��h�iC���@(4x�a��"A��&��m?Z�����/e��`%>-�AtD��$a=��s�3*�Eݖ~�鎼�Wz�N����s9Y�O����E|aƣo� {C6&1�V�%A��Ѻ�Sl��r��w����UO�X.�
���\&�g���5WV6���}6�&j��<mʓ+G׍�^y�nB�f<�Y���bB�%= x�&R�Yn��D%��z� ��KͩM���߻��sO�e
�E�$Q�|��#bGj����J�S������g`�M�����f���x+A1��O��	*�E����
��
#:��4g	P�>7׵Fc��7���9�!��)��$j�$gTC��'�� �/���B���?�B��{[�n�YL2\>�)�A��VBMP���Q��{iG�28R������E�!�L��X:��W�32�K1taV�%o�<��Xm't$w*�{{���<��X�{�/��1w�=�qr��'�2+�:��tOO��	"�w�R��~�\o_4i�l�0���J��'�>�	�����W�J�6�@v�}��U>�x�"�#����`�@�+^W��>�F�P���K�~�r�v��4���v-�����7Pj��:dc�N�o�EvGA>��%¾��Q���0�K{�ϒvQVʫ�W� ;g{���{I4%��p�B̙呬��d��b��xW0����j�����0bQ@	�&]�R�#�ڎ�%(+�*ҏ���a�I���nF>��U���h	�����	�0,!������F�5u�x �|n	�7�[1ym!�y�=�)�E�Z���3$����;�u��������G0��0�y��x���6����%��ܭ%`O�F=�y��T�ܠK��C���3���uN��0�/��FY�T�(��K�s�ἱэ�ݞ�@���ڤ��H9"�2	�v-F�uϠ����O���>$8�Y��)�����V�h��i�;�6�ӯ5�����v=�dr��}�b(��k�����)���b,~�*�����$���1���l
�k*c1�_K��R6r ���}��t�� ��s�A%][���N�M��(�G*�}��/;Š:�Vw_#M͔a�;�|HfD��[��#'Ε��W�t��s����_ȸ���Y(帗�}��͖$dTb\%��THn�� j`+  qֳ7�nb�J(�������*FR����Pg!�$�L�9wdJ*~�Zg8ڽDJ��E����r��1�~!ߠ6�ұ�H�ګţļ/��V���n(u!:���y��^53��0�}H�9��.�×NA�P��
p�5�yC�C 
����({[�a��*��
2ie���: `A�%vMZ?G��iUQ�pض0+X{�����gu�D����V7���Ԭ��Tc�aa`�$� j�:�[[5��f��R̨�Zj'L�a�q���v�'�_~ݷ����ȀQ��1b���p��`߃p���hR,�.��Ǿ"�X��h5U��Ì���Y���Poh�� �{3״'!̴��`��#h�*~0�D9��G�|j�ҋJ`���w�����m��<����
��Y�!���~O��F$�]�b�;� _BAQ�U�"K�r��&��%��i�/d{{�,�rU2�ޭ��c� ����u��D`�����lQ2`�C!��{�TLDШ\s'�(���!�����	���5� I/��'B��l����������U%�L&�~��-
�n8.e�h'�n�&%����������IK^Y��(+g���E{5�p+�[�_#�8�2�(��:νk)W�����T�_^)��8�Ì�`h[P�c��]�-�4���;�k�5��5^�%$�_,(�	��t
�&
�N+��zFy�� �t��(^�(�r?���.�V�0�0{#"*�F�~�x��AI�Z�?)n�_O��[}1RXPec�_٤;��o-��<���0i���}��Hx�Hhmޱk�hD�	��]�ۛ��8`]=v�8 *���sy��hɓYR~ ����e�VO��ט�J�Ip�2+<�;���.�)�=x��^�)��)?T�9I�N?�M\_B���Õ��5���K/�T�d��m���N.��Ѡ�Ab�o�v�`�綴\�<H�P~���E�c�Z�0_��p��N��(���C��WA�l_g7� �[��;�x l��;w8[���1q���-WQ8p���/$+2�O^>����w9q������Fl���Z�p<H$�Y�:���r�	��t/)q�Y�5z<�Og�Y�X��z��������L ���r�/�w�k�i��x#����Y3%r� |�o��4b��T��	�{�S��2O���T1�j��� �oٓ.����q={�r�E4��X�������9��p�t�b�����>�m�j�xl�b{�V�A��Hm���t�?�F[|���w��0�

���3omB����3��'$h|au��h�ԇv5�j��rQ�Ze9�[�Z�s�ũ���m8I�˦y����<Mz#9^t'#)���xx������X5��[Y�I�F��)����/7���l�.�M�fW�lδ�DY<�i ��q K+���Lc�h���_�o���)K6�y~W�H(k�/�z��aq��1)%����o���c���F���2 z�nL������q\��LoC/�J�z�t>�X.��`|2��ڔe m�h,�g��t4�*Z�4I]P8ɴ��2v����q�=��@���{����" ����?��$�v���-[�4 ��%
ٺ�-�igPһZ���������*JG�P���O�+#R�fI�4��%OZ�梂��&LAЫ3,�F����U���wC�I׊�� �B6�˚�|8�x�d�MR���9}�L�gT���"�<�y7��T�J=X�K�I)	~B^k�
:�9���O�襊�j���73=o�%��0�2��ϫÅ�v�t��oR�9�J�&j�HM����L��<�۸PP~3�����&��@��#uq�-g�ϸ4�$�$΅*��`pW
��7����P<u�#��)��W�bh�:�do�{���������\����6	����7(���,2�oG��M"~����,d�[3%�%#ҹ��k�G/-��Fw�������,9GJk�M�*L��[��oh�k.�t��9�kj��Di9�R�eSR��F�g$��ݽ;Zz!�ir�i'�M�0{ַۜn�-������!t���X�Y\5)9����k)�J���{L���eE�e���~�]�_��b^���]"��
�E�{e)�EV����ޑ�}=�mA�.ϕ�xx�	�^$-f,9��'�C�^��}����� ��ɻ}z~1��4����$ ���B~�Ț�(].�]��ӔoJ�!C��j���ڵ�!���U"�����a��a�Ģ7���eؐ؋8�u���pI��La�GP.1������d"u��~�� }�i�fL��l���b�>�T馆N#�)��f\�� op2x`	W��mU�d�0��L]���#0�m�˹-ׇGD��bs8M7��(Z�h�^�B?
�;�)	�		w���v�_v�;��ôv�3M��LDV�ӑM��:��,9v��2�������C�y���qk�]fO?N���{�g
�I�{�I,��<�5�?�:7O�n�O�y� �(�b���e�y��!�G"]�����MڶkuSB�NF��<>o	;s��,7�gR8;�X`.�}=��b~a�V�b5e�����q ��=}t�=�/씝��^��-�$�޽����k��P+�U�M���.�dkh�'���M��!�Eک���`�i����
>�H���_�^�{_!(P������م�p.`�-����v�Ys��:�����ܞ�4^�Nf�����L�u%�8����']��1����	و�2^Y�11�U��9���~��>����7�n8{������5s1��	�̋�o�ܦ�j�.��ֆ�? �Ch״��e�آ����Bl�>t�UH�������Pwki:���f��-�<T���,��f��W�m�T�1c�8�]�J�qﳑ=�&��q�MC��բ5�R�jX�8X���kǰ��Ճ"(8a�"1ׂ/%�:�.�>'z�t�&w�Fn8���OR&R�ͤ@諄�
)a2��j�uDd�,n�2h4��Y� �_w(�A ��A��?'�-[�E_q��F�1�Ի�O)j̀�a�Ǎ�7���e��g�xT�7$�DP���=����|�xH9���� JX�FZfF����;ǁ�!�-F��ֹ�E��+�����{@�ȣ淾_���>ɾݣ-CV��V�qWG���}�F��4Z� u��캠و[]�ֶ�3�Ήg422g���4�U߹�hN'�AQН?�k!��Xi={�ܗD����a%R1����}6�p�W���/�h�d`[�ڏUwd���{��(����n�8���Ή���:�n�<��5�)iū�s#���ߩ�⨫ǴB/��[�8$!^Ł��94���f�Pi"�]��²;6�ځ�&�C�J֐�B�f�����g߽���Md�k��m-h؝ָ��̋�����`*�\ŋ�a�	 ���aҐ��%ۋ5^�"�)Y_gU��/�^/,5Z�}+?/�/t��cz[��j����C��k��u7xmΗ�Gh�>��c����o<���]]W�}��ɷ��lu<i�+ݪ�<��Pˀ�HC�w��i����څ�!�bc?����U��u�M�*ky�Jk�7-_���k���b����0��:xm�Cx� �W�aJrk�ІO���ezJ��}���	�䓭�ʠ�Li��o���R$�n�톣�x|c�(7P0�B��҅?�7���v���2�����4pd���,w��rm��j���{�i�.a*����>��p���B�$�	F�����2���	1�P	���崀x����&�[��ȕ1%'|m>�z�k"%�/,��S���k�B�b�Yk5����h�"�A�ѿlXc��yCD�������k�H�����{�"�9V�4{��g������>Ǫ~�*-'�A<,��z�p����}�b�����9�8�@�Ν/��[i%||�>م�@��	^�^o��[x��t���X=w״Qm˵C��nxV�'���Ú�"����+J���岖�h�Z/J� ��Va7]��>�a����|�X��!�T^kRTӦ ��5c�)�8��GFx��Z�.zq��p�d��f�8� r��>���Ǯ�����v{(���A�Ց��`o���OP�/�V`��X��E͵* J����\X�W�~�=��S!���#ow�ѽj�+�ôpj'k� ���1}J{]�e\���PVT6����Q[&�ֳ^,cA��@���P����l()L|�/��G��M�G$�}{x��Rg��nUAΖ�+�j|ssĆ��ߚ��ˬ�櫰+0T$�5��ٲ���e#N��Vuަ�Mc߹�&L;#�{_Xr���Y}�E�L=!y8�I��ՠ�\V����n�6�ʤ�]ua���8���E5TmG۱���c���wlYn6�n�w��T�b�����8�M=6�K�m��i-*�|�X�������	V�]:?��N��!G�c	�{���Lv�͞����N)v���r��ǫ?��7���g"�A=���c������\���Mm�Y6ղ�ʿB}���i�CN�8��f�?$��R��=�8P�U�c ������:ڸ<iݬ�5ˈ����}����kP���OҊ,2�[u��3g�DC�R���l�4�lsyR~ղۦOS:���LV��z7��ݎ8�SQVt��,�\2%<;N���͍>Wp�'�
���o8F�]�g��}�n��vT��*�Oz7�XQl���.T�3�N�1�8�:M"�8Bb�/3�%4�;����D���!�Us���^ᣆF��3�����O��*�F;|��"�^ �q$w�vw�9,��~!}�q�*1�Pp�A^bXّ��is���B�h���[4Չ �nŎ�K4��F %K�x(�[)t4�8+��y�b3��1I�a�`�6}8�)�䎬&
?  %B�7����_�*������ُ�8U�7sQD�e��"}؈E��C7hm��}��R���j���i��rG2����p�t|j��K�80&u -}�aҪ4�#G���l�b5�,���:�u�?n(��:��¶�Vګ���&Sɋ~� ��ѱ+�A�ۣ�t<�����S�+�ڄ �
��$�ĚCo+�E�d���۟a�2�2m���%�u�7F�/�������vo��^t�͜Хo�̻4~�)�)�^����)��Q����]Y�RSܠk$y�'v~7道"�4�z��V�7S�L�Z���a8�%�Z<Q|))�L�	o���������ܽ3�o���e���9g���+�����������z�˱ �*	҈u�cj�dg��-��N��gI����J���
�#.������eC>L|z�Ziw��d�z����͗��v�y>�Y<�4�4/a�� Ы�F� .�ݛ�6n%��"��92N�I��@�h��C�[�%Ӟ5D	f
�j��G����b��x3�%a/89����cܩF��;?9�/�����S�!�wf���;�Ā�0�ܘd�]^aב֋B�&�
$�9�ێ\>)�s���i;��C�pO8H�@�E�nZ$��l(>�,��G�gB�|Icp�ӫ!�tS-��g#1d�Sٖ3Y��K�ܨΒ�mw�ޓ*R�����&��ف����>�^����{[T�T�*�Fyn�r荨�:��ߴj�/ϗ��������D�~���^�1�!x���1A��X}	��rx��؍���ڊ�8v�����lT��q�m?u	�GQ(���;Y��T��m��4Q���鹬��J�{;97E&�i(���<��r!�M���2���m�0>��"7O�8��h�~��)��ДL�n���=§: ohp�yػ���sxC��԰����8DƯGF�B��ū������ʝ���X;��|�{7/�O	&�b��3����#�g�0�Tmܘ礜���`���i�E�l�$� ux@�D>3��X��U��e\� �q?c,V�¼����S��!C�&�P�%��O���%�c��=f[�� Q�$nQ����g8\�|�y��"�m�QETx%�A�ю�s	�ԣo����*��>��гA��9�jw�%�j�:����X����,�'
����&���F���S~�
�+���b@_��E2��y����ɪ,��9�n֨���}��k[Oί�Zخ�Jc}�p[�}���O���7!L�X;�A+"G7R���q�(�k|a���O�E./��e2�Y�!�NE?B��I����(PE|wٞ�z�tf,5����YˈGʽ�����}����]^&��hǛ�%ϐ	��+�Gu�ɏ�/D8���b��J���-���Cm�׀�k{����?G�[0B�OA�N���)�F���2�b�����e�>,��.q�Bސ�݊LԨ�.棎����'UT��	�G%�;��l�&�F��܆+�/G��H�pւ�����AѶ�2x����u�\���3�8@7 �����:3���A���(����񌬞[`�2.8^�5ܐ��#"Խ3�+��娰ߊ������m���f��^\��=~e���u0;�}��� h��P���æ���� ������`OE�Gjg�!j'��_�mh��|���e�w;1B��_b�<4(M�[��z�9�O��I�m�t�&ub�@j��w�3�,�5u>`D�E7��ĩT����V�O�/��R��M�^���Z��1?�ylS��_�4��.��Ԅav����zy�K�
жY��M�눕I���ɢ��z���\)R�g0-��w�ր�!P%_+�����sh�A��B���7k�&�©,H�?t�b�����-Ԅ����4��n�U@�ۜ/��S���ѐ����BY�Nx�3�]��'.�!g�x=̚�8'��"�8�G3;%mx�a|����R<��p�rp�M�8�E��i.�&�=×�o3�50�4U������P�G� Zص�J��c!�a�f,������5T�\�J�vP�d���Βh��/<��4���s���0��K���I�`��~���y����sUܸF��`�"�u" ���I�t:�bZ�-�)�i�v�t�!�e�e��u]c��� (c���t/�C�Є:4/�����zۯjpL��	�4Z�՞�[=8�������_�a�����?��W�;9:a���V��1�7�7��/B#�JBu'1�u5��
l�������Qes�cT�⪭G�^̞P���������/w�2�4lJ�`�.X����qX]�����4&���62�y0��{7۳:��4��w	���J��߼K��xQ���ke���M K؈�!K��>����R����0T�p�f�1�O��<<�2~�}�r�DA�u�D���[6�!]�`�c4*ٯ��XPe�m�<��̎k��X'��7T,,怳O��U5;>�jA� �Q��9_9��nO��T�{zAAmZ�-K�}ȐC:$M�`�z���U��غ�l�D������9F��~�g7Nf���>�J_! �gD��'A;0�+QC��^m��$г�[;��5�84f`F^�V�;H���H1� �N5���'������Pl��C�����d{����o�����	�.a�Ud�t�5W�]E���͋��B����ۜv��=����ir����u�����þǊ+�������J�F7��K����#��^ �����>V����U��R2Ėa^�w���H:��Ҽ\�������{8aJ���}��Z��w��g�Y[�r�J�{�~�q=��;�T�v� .x��-wq���іmY@�1�[���yr{P*��
d�Puܑ�������� 	�� �۽���dn������<nz��[g��z�����l���~m��W �N�
 �� (�-�����?��TJ��U�rQ4��qf��f�:g�%w�`�L�W����cq��j�ů��G0�j����:#g�¸�����Ws�?K��]V��<m��6:�C�G�a3�s����.'#�����%����7�����ǚ.�I��un����{x_�8*�U%QQa�DQ�@?#\�P��U���<�y����PB]�5GHJ?��d1�s�~�*\�fI-h��jEbƁ�C��i�Ձ��T���^�F_Ҭ�6��9�������oX{���!��i����0��(^�gq���ԝ�/-�0\����[��wz)��C���qp7xk�
vm������s�8�]��{	�%���ր2�q�:UZ/�V'K������i�]ǘj'�^)mK�6!p=@��%����c�l=�X�&m}�$LjU9��P��ن:@�������9��i����	d설joiQ���d`���N*�α�B�	��.�[�}K�̅��Y;p��q�<�$�]�[,�ϗS���i��E�.�f��OopO5%��l��~U�;|ػ���IP�m���u����@��4�<Mf��@�#`۫m��RCg�}�h�
'۸{���=Ԥ�mx��ݭ4����fUU���bL�V�����CA�*o#̑B���n(��Џ0`�=��^t�=n�ߩ���\Q�k�Ugv(�fS6C>�ɥ�t�!j����=Rպ�#~c;��\������]{�[�b4��j!ǂ0*�	1���K��}a��JZ`�N>�K�|^]YN�U{uE�?vPF��̈́Iu�1YY�����_��h������GӖ{�?���a#��=��F��"'�y���\�osW|OY�P�_5�uV(��[]+�'Ɓ®���~/�4j�ٯ[%�#��3��@xqJ�B���3{]��$�VH�Q����R��b�]�����7u�&"4�M�"I�F)�S;.15��|L-�!��5s^*��L���t�!$��HJ��A����U�N��}(��£�H28��Y7,jLd9d
�DX�wd�&�w1� F-L��mNX��?`C��J{^����sd4�Ν3�Bn]�Aj2��J�Ϙx�.�إV4ſ�1�Ή�Iݶ��Bo�N����l^����Em���M�l�J�h���d��H��Ĝx�9F����^���јLC�h�s��0��M�ņ��HI����$u�/a�?A-�����~w
Q�4 �W������*����<_�3QGY��{!</�%�ı1SB�P4e���7�B�_��)#�#��@�]��%`cMSD��A5*��L�C�7���m��c�r.���Aa_n�����5H��OJA3�?��}���~���q�qD�#���q.�,���Ȱ<AW�H:��	Τnu�0�uA���WPMa����0���rv�?��x�;�YD�B{$9[;�J�,{���B-����������1Al���m
f�B�p�`����e�k���̓����S��S�����8��c>��nz���!�N<��Ha	�ˆ�������w�4�e����i�q��4\�nx_�//�|����I��zP�e|aw d6q�-�ʗS$�[��A��.1X=�I����5}���:j{Ǔg&���7����٨�?�7�B�lŤs�����kI�Kɠ��/'N�֕�q��a�Ӂ����`!��&s�H��'z�m~�D7K�=���S��C^��+:�Jr��ڢ�/%��� �g(�A�|�*4Sbv5S"=�e_��K�q�NL�����.�w�^Жo�3&�P�g�2|�/*���.[�늦H�W�V���|h�96E�-Vm✫b��������J\�cN�rs��70ЙۍY�C����3Kq�F�H�'���@$)@φ���k���r����U�E�c���>T���U��l��Wˋ"=�^:�h�U'~��P�ܺ����!�m!ѣ����^<W�w�ቡ�t����W^0'���eLq�v���|@��8sئ��C�Շ9� �U��b�������C�~m�l������g��믅��m�o#-so6k��]����IЏN��j^��H�r����^qy�`�����&�[��X��>�Q���G��d!���+����}�Gd��JTY�°t�o�M��y�Ze ��&�|�4�*>3.�ۻ�j�a�� e�K:���5��=A�n����9�+��ahK���7��[��>�����r4;�mI���YK�q�E��Q^2��e	��8�c�� �:���88E�0�_Fc��	7]�[��ʥr��XuV8���"�f�J�>�� �����΋���
 �_��f�
^���3��Ws��K�K'�H���/GY��_�/W<�-M��Ӂ��s�d8!=`@_F��&c3�F�^�����t���Nj*Q���BD�L�\mH�Aj��P�>�Nz�R��t`M��)���hc&�Y������޽��ٰ�lb�O��f4
���i���A���$j>?G��aC�(���y͈�{��t�m�;��{"l�̯I��'`����=�s�O�`
2K�}7~�|�
Ϣ���"^|��/`X�E<���Fi1E-��{��\3jëd��HT��CDJu3��GyN����"6�2WL���q�u��#��t<��$d^�V���8  �;]��x�����+����6e,x�߬�i����c�eS5 �Bd�c�H��:;�7�)񹗸��}Р<]�ۇ#�a�_`h�T�[k|�'�B�u(���G��L�d��JD��`���r�mu����uW���:�8B���>��t�EqY�b#�� �}�W#j����P�1K@s,�*N�5h?�G7p �S/K�p�"A6�*!<����5:���:x��Ye����8��y/4�<��?��~�����z���%
�q��}�a�x� ą|Ѹ�/�x�#�ME��{3���4P���c3�BaS��]}�LH�Л�ph��;O�{���#A��cB(^��.�γjeH���I����'#�8�4��U�l���3Ah��.t�eNn|HƂ�a^�Y���x
��n�P$�|̛'/>�AΎ�tz6�z����_dy��e�����A��% ��
^���UNaU2�V� �-J���Ze���VPeY��9�!M�*���Z�����/
jOr�g�����-��/�K8�B��4� |�x�]�&�oȰ�-����� /������ΧV��C ��wz.�Ŷ��96]kql*�l`����Q&C׊#��4VШ[r����a��N`�dE,,=(-L/� ��2cF�1"��@��M*�j��$�݅�Թ2��f�H��(���y�\��Yh��e��F ��CH�o�)��Bٵ���۽A� �:w�e�.����#�m$�I�$����C����Y�/̐�	!���Yh4�Ӌ���M���N�����y������LT>�6%���5�BA�B�W^rk��0f
:��13~B��)J��$	��k9
$e;�z#Yt{T�������?O_b�g��P9�/�N|]ƅ~�`Gu� �ϴ8o��T0lt�� G{`v�8��gޕ��;�m� �1�򡦇{`���:���)8�>ѡ!kq
V
�&&e�'VLXi�\���g�љ���7@@R���2`�ә	s���=�)��p�zQ0��4w�0cȸ��̽ء�w� �2�s�@������9G�1�����~���e�UQ:��	'��(꾱��vJ���2ލv�5�8��JU��	d�y�ՙ�CM�,pO�Y�� X#8$��`���AҔ�e��l�BT�`;��a�����<��Sю�RD����\R����U�0�j��ߥOG�H�+�&�yn�]���� r"�@	���Q=� "�o}G5򝫎���� <��ω�6�׀�g��ɹ���f{ y���%�N�Ei*���J>^�_&�xQ?�f�`����#ǎ�r�	��m��1/��eV}����,��_!��D�w�Qؕ��P����'�y�n����EN(�ɱ��/�`�Z��W��N
������q,0w�X�#��m���΂��y�y�B��K�@|_������?6���	0wܖi?('��/�R\K0$����̔���� ӉM�O�u��(R`å���U�0�nbs�s�?;�C��	7��R�R9���m�iK�U��/�(UX�����L��p��zwO`�@��G�ȸ.��z�����AHpi��$�^-�ꗨ$��go��i�<��Q�E�]����N�ŝt�s*����w��R�UN�qK��U��K(�f��6�S
��!��8�CƄ N4�'��;���g�� �#/z�LM��ˇL?m�{�����՘Դ{(UO��If���q:	��1Ji6#�w�/����H���r����2p$Dy��D{��B���'o�i�����+plD�<"1IǗ�dn
cG��Zm��i?ϟ%} �d�Q�<պ��T" hzp(dq�c��Hm����'���
b��a�n;���qN���A���C���SD4�F
�r4�EF+}~gr����?C@�-:5*�f�aEr~B���sDSqt@1cx��ԍ<��'i�]�����^9E�ne4��4���'Q��ɹ���]��t��
����%<Y�0*�>����P�:�n��)����E�ȉG\s;���g9QlpC5�^֊���2�2�.(�sg����� ��~j�?C�^��ס$�?�&L����_�'Tl�y�R6D�b���vx�F�[�$����v�a|�4��*��H"+^Ey'm�XtA�����tmS'�{�6p�<��U�6�oM��?�LQS\<�-K|���0�E���KÄ���L ��؟����g.8Lb�H}�~C+o`q���DCfv��*�|5~ɍ37��&vb^�w���u`��FD�b?b������k�C�?�^섶b�$�^�UK2��R&����`�õ�c0�F���I>�	��֨��=K�Nc�g���_)rb������ ��*��@�zY"��C�}�V`_%���وzuIQO��޼G��^]1��h�g��e9g�s~f�ޣ�JzV>�N��*j�c���v��Ea;o!�����6,ı�IL�H����H�~{��E��hSG�Z xѢNK[u�qf���,�h^�[IM�1��<�J�o��D��awd:|�x�x�z���{C
���p�7mIJ�a��;~���*��.�D3�s�aI8��X���^g��]˽����*����?�}�C�����V�C��t�����S�?ֵK�Ƭb����� �vPM�F(`�50	���>�c2�s�������R�NP�D�Uݿ+'+�>��K�BA^�3�O�{":9I���a��E橇
Bꘔ���#'��im�D(@��֝���療X�p�/����hʅt)�?�a6�0s�jg+�D�
���d�N�����m����E(iu��⪜I>���+�鞰P���X�&�ޖ��J��R�azVԶ. �8���rvr�ͱ탄{ON�n/���3��꧷�")Ӵ�,L�n���@P)�Y�H|q�ܦ�H�?'8�	M��FZ>�Gd�(yC�M��7�sO�ۛgĸ0*Ta `}�ǂ c!�m0N���~���Z���>pC!���:N`���J�$����<O���</1�U������N��C?A���n��olzd_�-��󚓙�'�ƨ�?��0�v"y���z��K/�>߷j�B�h�ya;=�.�k(��QL`�4#ê9~L�AW��;��>��[�D	�g �z��*mTp�;��ݕ���WS�*��-�,���\|���F4���R�P��xuϮ8MK��#;�Ɩ�_�QYViXN��&��uFZee������<
q�.��@�\��*���>3!�c����S��.��o��-��\+�p� ^��p�1:����G��ZK��/��)�����#z�g�֫U͖k**_��}v3 ����N�FԦ#�^�:�]E%�:� �����ya%1urM�Q�Ç)He)#{��t�[���]��eU����}����Ћ�m��qj�,�ӕ[t��8���������o�?X}8H)NU+m��C&�>�e6����;�A�1rǬ����H�"Xf1o`����Q?����nQ�^=o�Y\����(���N}N����\��l���U�"��¥�}@��9��N�L�7>�U�<�=S7��p���(}�{�p8K�j��
0|@�����p�k�8{V\ɸ��2��h{��<5l>s�ꌈ�����l��1kg�C��Y�ZB|��o���t~mӈ�An*~�!����_ߘ��l+-����Z7�؝�����_Bj�V��w�y�o���Ll��w���P���M�F��֩r��@���m�XZ&tN�
3I���9{��[����ӏ���h���3]b��J�@��+�!�`	��m-/wdh̖7 {t�e�#̒�if���5
Q�M���f��h���i˂_�NB
�ڑ�ZA�/u(/���8��߭%�TY����6)��|�|����r��<�L�x����uח�aG{�D!�X|�׏����#�'>�/�~�L����3�em6�vq9[��NR��р�~`5�'�� �J�,q�0���` ��,�3 ���9�%�7�Z�5}J�$gص;��=c��,��"�˚�'A����"ծ�YoI���骶��&6����@��/��{��(�bk��#���9�l®q�,>�OW�s��U'����K�-���Q&c�T5
�18���su����|���[1�'���Ɨ쉙�-�zX�?Qf�MEs���U!��݉fЁ\�1���$"g�O��&�k�Gr��*�Q�˫@�M�{#��v��8�ypa@F���y�~��K��a��x>�sH��/�[c޺D)�4�!�`�1�~H�"c��ֲ-�/��V��AQ��n�,�ɦ>�k:�ύu��g<��m��c�I��"$��C/t���l;���UHO�_]�m���	� _�������QP�>b�1�r�������sA`�W�tC��-��m��9.��I�A~�}I�����W
hl$��􅽙����k���4�d�Q�H	����}�C(h�sOB(��}tF�c��O}#��,f5�Z�#_ҘJ��:��hr�o��4�ދ����>�%X)�Qp����v��eY������<�]�5}M�O� ��vk��F1:����ȫvU��ӴG�����Ǒ}n�R�@ȃ�����_��qRI񖐱�V��A�����`x�M9m�g���u�b:<�X�����)K<����B(����K�H�Z�i��"��(mB �ǖ������#�4E��&��<z�Y��)dr� ���F��*;Ik�c�47&Om�U�9�;�5�5�>P�#��F7@�b�+2�U���TFfW� ޿�"2x8���z2©E�ɔ��C�Z�?U�XQ���X(�P�îрD�#T�'9��YCJ��'8��0Q4��g�?��´�δw��Ʌ3�����y@Ȳ_�M���}��o$�$SlsK��9R:���[u6�i��ZΜ�pB��|)�S�9��qQ�z��/�%{�e��⟋�6R��́a�s�;�,Y�)F�iU<�7��L����,���0��\臧�^d��7�EoA��xvROj^�/�(Dm�{��Y]O�q��ꘑ���[�9B6�kJ�#?N`�s	 셑��2��E�Y?���%���-C'@ 5���Y���"�>�%�!���d:��`kWI�|
�Z���6?d��#X�vg�ा �9j��":k�����,3��i���`~{���%�0����s�N�+;���a�Kf��j"i���=K��pT�2��!���I�z��Yi�����uk,�ql�9B!�ΐ�0X�,ء�>H��44w!^�F��d�+�I�<�!Lc��{^�#�昊�JR j����I��5|<L��]=8ώm��G�Ճ�Ο��7�������X���p�V;O�.�s��k)L�$$]$��V��/�X1Wk&�S����%+��$xR��D_��G��8���ڵ$T�e	�䶫�G�!�)E�o�l#�t�������Zs���̽�p���W��&��1�헾��Q �}k��;ή��d���G�o?G�r�����v���뛚���-����0�� ����3}~i��	M�5ؿ�+��1����D8M)���Y����fk[p��j��I�[��U�C�� i����T^~�[&���:g{��T�0�@%W�͕�����ȝߙ9l�2���s\G��jyz���X���9B�v�h̠
�6�$�ۃNn6�ca���i �D��;�����z���$��E�Ax�5���{f��.�����b�W.���y�:F����d�j+��u�%��D��M͊}��r��c>�4�:��)O�rھ8q�Kt�l�s�Q�/��P�7ܿ�+��f)��U;!)������J~�DR�x�����T�L֔�g��g���:l�]r}�y}(�:�~k�'&��й9���kYQ�?��|Z1�Xyw�Sg��������Y�����I����,�A���T3T�� �>��x��s�m�7�Z �"�!�iD5�W�TQ���и~�<t�L�]���Ul�0��;\�S��E����.b�����$F�I�3�;f�F���_�/��^
\l(S��"ͳ����(�y��"�?!͙7�n� q���DG#QŮZၠ
-5{0�:�M� (�۷�R��o�|�#!WehI�mvu�z�d������ķe�3��D�˔E��G�:�L���3<�۶���4;�y��K��o�P�b�4�)�08L��0�u
��C_������1��s�7�=r��t�)�����CZj���t�䤦�b��>�>̫+aV>���|0�x܄\vT�d��Ct�;�T�
���D�
e��rA�ܕ;���5�^{����g��_p�1�� cf��+�,�G~K�c{J2\�����fF}$S���c�K�1��rIl~	�����Ϩ��P@�*�5H��K��9���td���w��ޫ�{�- �YB��Z�E&pԌ��6����h!�A��s7Q?)@���3�3�C�yg��)MBj�j��M:p��pʆz���_�Z��T�eg��^���kx�˙"�YN���n��Dr]�@�[���Ԃ���9�K?�j��ɩo�,|�b�+7��U�T�8!������r��O�f`������� ��0|O��P�.ua/����aW0=.	=�~�X^2 p|jC���c� �}<S
�f�_��~@l9ӏ�����J��nK�J!��pJ���3+�;#��h���iE8������B�⨇b��llo��S��_�>�h�<�x��Z��������؁6�g���Ք�ݷ��_mr��/TQ�B-�'Pd@���$aa�I�lBG{Wp�;�e`���F'��j1�h/�ƀkn)*.�=��ܜ3�(�vw�*���j�r<0��L�	