��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��r��U8'��e?�l�^gd?�����Ժ��9�f��=�Q����[�Dx�$���wM����=ߧ�+Q��b�V�.9��]��I���%������D��cI�1�#�h�Ir̐ξ����$>���*� U��6����Ǒ��U��}}������N��vL��C�(`	��~L3h&]��o¤�f��=ԈW)%�5�q�x <^J�X�V�>��OM�>�<Rd�������`	�/7��r�"����,��0���ݹz�!)��69�G��¸e~�b��)��(�cr訛��£���XN�u�]��n��b l0E�?�2�fv����6&�T��4j�Ҫq5S$LY:D%�m�-"�e�X]ݛ P�h7r�)�a]l�ɼ���7)M@�ղG&�X���&�J��������ب����8V�c��t�^�+�A�
�'�N��=�h��x��O����R�XY[:�d�Gb�X�L$8P��0H�����1-���=W�kGXc�;-�A���%��溮MF���-�hL�������U�B�����l�˧�`B��Mͷ��B`'���D\�v��=I�z��eaƾ���=L!�u�tE��c�jiu0(ۢ�ƔH��L|IM�FR����3b�tZ��	��I���	!���-����,���7*qTl�Y�_�����ER3�8w6�WӚb?���)�%5C���M�O��Պ%�:�>���`���Em� �-	�C�����/y���	�F�Ey�֞����;6q��+��-�l�ೆE:�yz�S�	RL�Ь�(u�ɯ����C?s!L��V&a$IUI_�|;kO�w[�>��ʭ<@@98\ ������fFћ�K��M+(�U�L}%f�	 �2��(�w"���wSP������oՋ��"��=@9K��W��z�䨊��:�I��wxlp���U��%t5mG. f���@_=��L�CJ�A���tR�%�rr��]|�}���HVX����q��\L�')���}ѝ�|���,���')��J�dv&�l\I�?�\ ��g�tnƢ�`�c��37j^3��j��H�@곡n�Fnt�X��#�^[��݅Np����~���VS�A΅̽��H~������� go�2g�����BTv
�Ӑ����#�i#�q�_~��*�y���l�R�[��B쿉N�/��A�~���c�ޮT���Y!>�b��Q��>�>rmOGl4c���LF��
�Wu�k7*[�Ђ��f���Z]�{&���!߭���C\�r͂e�6�����c�[���n��Āv�UU��v����q����Z���26̆�����N{):O{ѯ���S��6��@��K��"x�SvԚ�hۼ3��]w���`�G*���C��92t�#��7�T�܅�Zy�:��C$�,΃�uz�u��gm�DT�:�qNO�i��nb�n7�`��cH���:o��)q��4�X�9�b~�7u���T�}�B�QL�ح@�L�0J,ˤ%��������TP��K�r5�k�r�W������K��$�S�8^�*��d�T?WہN�Z E���X�!���ݩ�Y5��/t�$vz��R��W���b���q���[ԗE�+I�3�96�����L�֑l��G�"��7���H0�Md�ݶ4��6T���qXO(�՜W�	3Mp���;�+Rх��	R���f ��re����1�WZ�3p���R�	��k�=�%KX��^�9��G%�;[?���0�9�Tq "� �z麳}3���j�b$#�p�K�&O{W�{ŕ@�Z�@{�V���ԓN��a��������QIʤCo�&�Օ��e�ZA�8��J+�M�gٹ7x�KeO�3Mr�0¯��.����ձu�N��b\�����!�r������~�s��B�@�84�ܧ��v:?��ߨťMrJ3M&�'��Z��&k�,�Kݤ��3S-'���'��e8��@{�s�V�5>4�@υqL|�M
�|w�]���?�;�vyx'
'�Ŗ��A�S[��3��M�c���xA�{����6$i�k:q��'qY�"bm�yG;z���Ӱ��i5^���\Z\ީ�I,����]U}�����h;�Δ�1�������#-��q'�}����`k���g5�i��eVVY��߼l%|�� #�vq�+�-�e�U*���%>�ai�ژ�E���H��!�if�$X���Ň���u�����/�CY ���o#P����
�!�BUVq%;�F�}��\Cf9�s�6�<��,��M��	��=g�ux���8��bU�����v����k-��¹�7:�8�o�,����{�O&�M��6�����]�^�qP;"�d�P@*T��õ�E����
�^�3nM��d��R<Z��	�z,��γ�D�\0A���5�U�$����0c���� �?�۝�?��Z����\o��[�	�����K_�D���m�lGP��Q��bK�==����_l����/����!�vIJ0������Ӽ��rɨ�����Z ���']@'���12�L�MI��\�\�ߵ�]�3x~�����_����sQ�i���ЈnӅZ��EM��ɦy��*E�7��������dQ���t��<x�:Do�+iU�O)��$${_4��#��+X�e6[}� ,��d��\)ꎄ��)3���r����uI������{�+�j�-L����
`��b-���l ��� �X���%Њ�L�:z����F�
����8�`e���W&4�l�G��*%to��z`�-�ʙ,��R.&|�Q�c��iѭ��k�]t[-�Wz�{ɫ�"�Pj>�.�S/�y��;�3}ۡS�F�0b=�h ���*v?�}pR���qs�,קKY�c�7���I9"c��ռ�J}a��8IQ��ԻA4���V����7éָ
��H���4�Ҳz�\������u�cbr�{���5ꟶZP}`��ܡ��<��q��;4)W�I�_Ol�{����9�\J�Ɵ���g憣�k�u��nl�L�Y���I���20����ӡ��ly�
R�M?�A��pW���G.���y�Ro�
�[TϪB���FU�H����xh�xp+@�M�4�]�1�O�濡��� �N��7֙�$���oC�`[�<��U��t;�����b��H��Q�=�^��/si>{�f�k��.��.0�哯�-$S��*gj;�og��Ԏ�G�%'ω㺭��.�A�BU���V��c�vm�I�3��tӀ�5M�z�S<P��|��)�?^�JJ;����H�W�;Y���,�kP�_@�zn�v����/��uꠠ)�Mrb�^a��2aR�{Ϳm��M��P��*h.������,#��<����bR���o��`�S%D�c#ps����Z���b��Ҥ�,~`m��gP=���e$}3+��߆x���!W��ˬ�vp��lpU���f������ �,,	;q�暛�����%l%��pL��`+41d�nׅ@9�K,я��Z��	#�I�)-�)���^vo�&l7��?G�	ne��x$��CA��Zꜭ��;A��1�l��^ƜY}�b���~9h7���Y�TD�jА�;d�aw%�V�g~���u�R��k�M�ם��9����J^�bm�#�ZFJv59��0�^�V��y<L����<|����qCY4a�"�S��K�[dڥz�������hW	�L������Tu�Խ�4 �Mz�b�(���~���E��E.:)�+I������H�ħ(���:�i������ ��I|�j��E�����=%y<�苸�Spu�� T5�ԝ$d�
+��ݴ�)�d�遹K�k�?;��\s�DZI�Ȧ�!%v���l^aO��+"�{��,|O�
AfN��f��'�U�)��޻�������~�}��p����α��ݼ�:���Xx�;���7t�q�<�ŭƾ���M�V�<����7�����g��-�:������r���+�I��7�^�� ؎��R��S"�M	]�swOZ��G����^�F]�"��`h�����&�K��|>�Y>����c����-guC����Z�Hq���M����`�{*Zr���1�%V�#��^e6����K���\�XG���3ވ`+����Aj�@���W���ګ�Ӡ$���s�<-�`�6�um*�s:�2��Il�Hu̶GҀS��K�(Q�F�fc�X�s
�#��=+�B�j�D����a�e�l��������I�@��pn�m������Z�S��'r�vd%�j{D���Ŗ�����+�뫂���)%7Jw��'�?dʷJ��1�9�=,�� �K�{�T����F�DW&V �4E�φ�����NH�-�����t͊]���6�X�D^ԕ;7H}}�<��ph A}&�a]��(�T�37��⎠�C���;�X���g���V=�>�S~��q�F�㾯×D���2�k�QH�PS*ךܶi,7��91�;!��z䆽D�4�B��Ԡ�A]W$���C, s*
*�$Q�+'^B��O�:��
��B.�C�����v��w*���2�1c55p���1Mє��HKq�.3`/�}eqx��.J!�>+?A�Á� 5��}ÒNR?�@�+]b#D��7����3��ʾ��0^`���E��E�+������v�4msU�Vcu�0d���z*ٗ�-~� ּN��0J��C��%�U1vD�7�;#;LJV�Y�V��{�hf]��}�pS�A���>�y;�DN=����0;��%p)�m`x���GkßJ�~�r���ʛ�^����E�F}�zz�$Z���<����x�;�?�-T{�\�|�j���UL\Jv��a�7�����e�������e�~�Y�$��H����O���!��O��Aj}I�	/29���>�kt���[)�j��b_��z�#�%��)���j��zӈ���MS�MS�M!��Z�+���H�Ht�!y�ُ��EI���c䶩b["E��T��$��Ѕx�7 i}�wjw�8,�G�Y�:��@_*��М�B0e�Y0<$�Jňቮ�?a\{}a��bsz]ߑ֧|�',S*W,�-L��?��yv��g���rSu\��2V�;�f�-��TePU]:,�vzR�n�'󞉺wĔMݤ�$���8�]ԃ�
�p��/u�W����YkG�YED��a���YF���O�s�5�t������;_-Z��˩*0���Z�*p���x�:=R�P:�:�ZQW�i�^���EҞTn������FQS�X#U�R�j�M��I��+C��2 vu<��	t�N�5{V#"���p91 Ś� 
�ƱFv��s��̚��t	��?�}�й �_�V��"ED]+G�|uy�bdG��bV�5�8�D	�v�4w�Ȗv)�^�{7��t�����\o���A�
��!��w������`b3iߦ^���}S�|�},qm�ٱ#�X Y�E�X�vT-��wo:͌ҁ�-�����Gm�A�,� ?!��"�N�]W�\)����1dr�~�t�@x�+kO5�2�*;��Oг��Q��$J�g�"A�E��E@��bWm&�Ogu/������3%�'���ހF60�CV�>�	��> e�"��]+���Ɣ?M,���n䃳�]LI���=���7�d�yإ,vx}�¬�A��Lz��|D� ��|�%ՠ�<�g�$`潫� 汮����Km�A(�m�3nyvq���Js�W��Kw����'�
�>>S��S��HBfJ�8K�0D�~�m�3jC�Ar�,�62��.�'3Z����
e�����ǣ�)w
����N9�!v<���n���slCA�����?�H�yn�UnH2����C�{`�g��#$��"�0]���x��l��}�	�`Y�)�L��0�9FT�)#0[���ӡ(�o]=�:��#�n�Ì΢)lP�!��a��6�\S����������≣Hy�S%�F�����X�zF�q6�.�CR��xU�O<=u�/Ao!' ���桽����r�q(a L���:v�AH�Y6=*�	eRO$�5Q�kL���/�I
�x!���z׼��#��`���:��&�ҜEL�Y�}��Վ������HE܍Źz����bǄHi��?�}���?�8����L�rg��,��ơ�\��g�=�>ƣ�����`!R�kOj����ڛ�J�k3��
�/5���r�
D��\V;Ð-���M9��dqN��I�\��}o�ﳄ}��ꎩ9���H8��ĎZgB�5m3�Vg�j�N���%`��H9�J��qLk�߲�l�L�1�w ��o.d�uUu����y���Ǔ���z�\%6ɡ*� sZč��N�1��0��
���6s��ռ%���w "{�G/�2X��os�Z���1�D@$�#R��ZA�Y�V���߂�e3a�s /$���q��Dh�n3L�*�h�:i|mG��A�V��u�'��������&sͧ-k�l��*����im6�mx��=wj�/Ԡ�q�0��2���Lƀ�P��e����	;����)^�1�#�ˡ�&����.�$
���q��6.������l�ξ��;����4R3?[9����Ω7ֲo���J��j%����C��TrD
����$�.z�.q����X(N��Ʋ[R{l|�o�`xJ�Е���O�1c��!����q%I��W�迾G-�_���Q|���L
CÆ�ܯ�J�Н�?��Iqu�1=h?�$��X3.M�~�YS���F^��]�'���R�_ ��@,�����`@T�J_]��zOK�D��/^�s�F�HK��i R�o��e?�=[�V��b��M��x�p>��[��$���oFFM����(M�������ey�
�A"yO@)����r\krpi�0t�*���u6 f��$�c��/S�z����inO��Q=3�����y��)wʱ�pN�8[���el�(�M���@݁t�)�U/�!��l�b��-U�V*,��ɻߵ��^0������@x�H�����t�Y�w_G�N��Y0�g�ym����)�d�6�s�I���L
TۋHEnC/�Qa&S����#��-��{���{Na��S�\ݞ�	�E���ln��xR��[�r�PL���:���L�x�Ư�.sއ=��Q�,)��^FP�P$P�ilq�O������{H� ���k��
��=��e��� Kԩcv\3�H(��1YV��,3�4M~7�@���k���ǡ�h]2�Q��~{
0/+2���>�K�\�����1_��Y3�aChr���k!�{a��I7�p�)��lX������D���or�y���,�&{E�3�ŕZ���I U�;z�֌��K��ԝ��YP�Ӳ
�Ѡ���2����wp��+)�����{������o�^Q��u����J���mؠ��1!���2v���ƸgK���G\��S�,c��������������3Z� +{3%fμGJ|��%��Эq���L��]���͙�w-�U�pEN�0Q��q"�ӧ��я�E���V{/o[�k�ǀ��Un�.אR��=����ΐ_A�֏=�ږ�{{�ے��OZ|O�}����[GI�?��B��$�W�In�2�CK�&�p�����i����&%/S��7�߹��������I/�j?kOt�ks,֟
��-1�V}�����������Ezj+H��`  p�t�ޕ���T�x;o[_@��K�� �F�?���9.V�0�� ��b��˛���#���"��(*�ķ�/M=���ZE���kPC��d�uy�{�#u_�
�Ɵ�2�ă.�^�X ��ת�F4����1��Rۛ���u?O���K85;b��R��'�� :d�>���Z{�C;��l4�׏���񙆱��U���̫�d.Y=�~)��V�nuE�WF���������]���j]��_<+C�W��@�DI���%�ƾO��\�3�iL�T�Dp��B���;/�1j�ƾ�RY��Ft����/\&��k2�	{�Й�Mu��9��a�}�~����6��ź���� �4�6���\�q�&ԫ�b)/�k��X� 	_{(eU.J�T�罬���2s��V�4�7�|S����=�� ͥy��Ze.������������HR=|�!�����G�TY�}��HN�����x,�U}>�眒��� a�ZH�� ���O�C���񁙿��*�
Oc���� ��%��aJd}����.h�S�'`�MM�[:G�QQ��D�Y�2(�~C��
&�D�tx>�����Uȓ=�gN�nlH�:r��v9Lid��3q�3%Ͽ���L�t{�s�f�-�q�������#W*W�Y�<��#��1u u���[�:_8Hs�gJV��}��	����.�[��t��]���ߥg���"�E��~�"�Ϋ�Î��}���Qv�[�(�
���m��x�2���yj�m�ˏ�_��/����s����*\&Y�[ӆԩi锋,�� 
��,�"x3j� �AV\
Z^U���m�^�ٔ���]�R�Ώ�%�f�3�Z�ڬ�f@	fNY��2���u#�U�w�K?����G��W*^D�'�%@l40�l��u��9�a>{�yI��:�r׼�,D.���,���|D����.� �Յ�ȑ�R�!��-�//�8�0R4t(���"?�ʒ��w�aŪ��M��Oj�d�2��=�܆��!k