��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>hs�*�U��Q���qh%ws����dު�����j�"�^!P!�P�<�?��_�x��4#��hb�teSV܆�=� ��(�kSx^~�^�eyL�iTP�Y[M2�;Jqɡ��2 ��f���s�����c)���\�)�Y=vScXNt1$6���X�S���qmTy�-����	�F���w[���2��g���,��Q �:޳j�Μ��؞�OM�J�ЉV�������ZH(��$�K� g��DM-�C����7���N�(��R�uF�����C*������H5N>n����������Ù��Ya�a�C�-�1��W��ia$�����d�E;���Y�:�$�tΚ�&�}3ӱ"�i;�P"�M���)#C
EeԹ�<p�B;�p/��+���jՖ9�����k3������W}i.�t����[!��ߪf��k������8�����%���A�u���
Իw�P̜06�'K��>r�U���iV��
q�����7��F4K3�/�+\�e��aCp'@��~����c��OM�sM�O��M�aR#�����s��=����I����_k2��TD���S� S����ud�/�������:�� �J!��r��J�5(I��/�/CU��b���ǷF�4ѷ�>$��pժA���8�.���z3��ԇ���=:B�ԪK��Sw��n�\�V69$��	s����]Aۙ�Z|6�A6`�^�5S�@�e��_�	�ȍ�s�o�xWu�汁)MWe�RI��_A
�>��:��J��U�"�c�_KfW��*�JZ����~(�������W!��.!�b����{��O*�b��k����B�=	h�*D����ܔ:7�׹y�T�A�!�H���W�j��Z�+mx>ÿ�����܂�
��}"�tnL�H,5�������O�J����uHBa��΂�>_*�yH�
�Ķ�t�h�؎���˸� :@^�J��_J0/K�l�SJ�sC�`�^���D)D�ӵY�?���o�L���k/����~�{2���x�q^����FW����p�LI��μ�M�Ъ�u�F_a]�@f���9��ۓ6:��S��y{L���y3Ħ��
�áJs�` ��3��q���ҩó�QM���#;߳m�#���1��h�P�e"��PT�+=>��k�C�еͤ��ط��(}��݆)V�Y	�Ba��W�U�Q8��#�	��!�*͕��j,��/�X��擿��o7e��Hm��g�=���ҟ����aeu�[:�V�a5�R&�-�A�'�hl����G��n���_-� I�.0��6�AU"�fC횤h|"�x��2�]N
s>��֬>��叩u��+���)�E�9SF���ܐ`6F[��I�|��ku�VV�i\��Х�#f���m�,�۱��8�v�f1�A�dl�.�}�#b%VX�G�}����|1��D;$�M�쀾�)�:̽�з=#a�G7�)�;�qv�� A۬�� H��{Yۥ�X��K�����X�m��/�!]<�P�c�9���Q���᯴#������Hd&����Ğ�W[�yÜ D����~�9R7 	U�x��A��..�I����YTZT��Z�l��k/`�Z�#e�\]��S=Rlz$[]�.�$�G:�0��1�Ԋ�#�w��h9�s��Uח�{ŏ������	�4'V�5�<p���8]���U 	R��kiH�MW�K��	�Z�m�syf4�8��@���P�̚q�S֫�F���� �X!Y=��0j�����d"	�xCn=
Q>(���h��!������l�J
g�8�_eZ�"�^�ɦxt����0�#:7�^q�X<z������aY���2#�g�60�m��ݮv�_��7Xk*PC��ڋ*j�2m������y�*d)8���꼞�?���T�Y��D-N��`�/�]��8��[ʡl�fo�ԕ�=a����p��9��[��wֱ�X~�r��y_R��d ?���D�����?GE9�ir\q�[-�K@i8�fUF��-��ώ4"�ފY�!�3lYOI�>[����Rgv��~��TRy��?�m��tx<T�*x0�30˷p/��<�a^�h ���d�h�¨7���W���֘���©m��9��Q��J���sRY���SS
fn�4O��� o9�k�l����2����T�Np�m�fʜz�Ufm���߂�S˾�%�	�o���g-���5H-ZV@�Z4N/[�d�=���K���&,�0��U��!��!�^<�z��#�m�T�nj߰;Yw�kV�s�	"����8.B�\o�v��E��j<3�&d0g�_��߶�4��or��gb�s�SU񶈖�j��~�w�����s1����p5t����Oʴw�Lymn�>h����"�)�&:؆#�����j��\���-P� L.�or��H'�X��mq�E���S\ڪ����kB�%�04��ĳ��{���FYЉQ�E'�����oe���Tw�)y��%?GBmw]Φ�n����^�C�/Ґ�U%���l�@���u�߅Ν�!�0�_��`�[�q��;v� ��$�cB������W�ܦZO�M��,�'a��$fn���&ZI�'�<��r�H��Kc�D�=V�� ����Nj�/"��ɳ�e�_]eR�I щ�)����c<��)d^�E�u��&`S�8���	4�4�S����	�X��O�t+����X�i�)P�$D\�"sYL�@6�[��d �줃Z�NH��F:�?���w:��0�S�ȆSt6��h�Q@�6 O��&o@I��kQ#���q�a�2�m� �d�������Y����5�n�}$=�����Ød���}� �('����r\��j�)��`C_�{n�d��)������k+N�/x�58�ߴӈ�a��l��E�n���]
MT���Ln����]�i�4Z��l*}w�Z�7�D/x�| k_�������2��+��y�d����N�o�jw��1����})���Ω���(u.���`���B�����R�Ӣ�X( �\HI_[YC�J�6$5���̓�g]*x$?��K��	�+���ta�o�j���\�$�Dд�Ƚϳi׬?�6B��Q1��7߼<�������R��a��@�S ���s��7m
t<郛O5 y�d�{�U/,�P^�,9zPKw��5��9��G<���Fe�4!w��<�;��/]3�<�q�ti�R�ѕ�k�r=c�Ѡ��@w+Z�:�d�eaA�����	��@[`����:Z�Ș�{�ƥ?��9[��I�B���m}�Ƽ����R&���h�1(�f�tK�82%*z��-|"rρ��{�{��5�ѝ�%1I?���96{m��:�:��Av�T��Q��;��$��uk�͒�����4�����'����c�&G��������˅��P��?�i#$ԇ%s�t� |p�CI�/d߆������F�ˢk2�""���rp����B%d�$�`����}+a���f�f�����j0��J0�ΰtc�O�
Ht2���� �p��x<��mLrթc�h�t��/wQ�����2�T	'뺦0������(���P��}�noбLi�J����6�E��Ϊ��b�Eً�P��k=��@mUu�0zn�m����Q�pb� i�/�t��}߽.�z�W���LH9ͬ/l�/�S���"O��馸�!��\-61�E�3n����I�� �k�|ث��h���	� ���@�a@�nT:9�2��9ֳI5��N�,����|��G�au`;�*�]_��A5��[�?�	��4D�rxr!r�b���a2<��i�-
?%���[�m�e�B�~?L�'��'����(�@�����Nt�E�_A
�P$*m�Gy&$Ơ�]��C�ddCӓ)��[��
�>`����������vh_-��f~w-�Q��,.�Ҙ(x����DK�/���b��zʈE��p-Ń��/O-�E�U~V�ϡ\k��d@�ļ���F��*�3����K$P�C����'?��A����|r���%a�?��im�/�u:��*�h�J���t}�E�r �ν�+9�t}��U�f`�l!ޔb�f�6>�5�Z�8%}�3��q쌁\aq��A(�6ƅD�1����)߷��P��U�ѷg��U�oJ���$ɢ��w6��,Kf~��h>�̊r�T��4v5m�k�V԰�ip�lѮ~Lp�]�m��U��[ݸ���N��<�C5~jTt�fsxކ�*�Q;��>�(U2�g.��u�w\��
u�?�*�W��t��]o�R��93�b���N��#l�Z^�S_�w�~�}��}aG�8�����Vc��;ԲK'-rt9o�� p�<te���R��9� �u�/C[��l�1~�����́Z;��Y(�d�)ޜr0����My��m��r̔;�� �1�������ގ'pQ*T?�|� ����6^��C_���?)P�o��N�TNp��b2��D�`��� �[����#��������Y�j�3¡�s�P���t)�`���[5�1��C-}�1��V��"�f����=��E��-�\���"=-�����!��i�'x_y:�`ƻJEe����Y@1�߹�#��:�N��F"'�wo�����8/8~On������8�k!��# �A2�[x&WJ�4>�n��VXV��vMA���4�Q��,��kY>����N.�Y���t|���Ӧ��4/���L��&���Y�oξ�L�"��,ӌ�:5��|�^k�/�J�.��ƚ�Ơ�~��j.5�{[��p�����.e�����N��}M��V8���e1H`���QUm�uP�q�����S [�45�FRz8�!ǞD��8��ɱK�܆�Ú�_���AI�׏y*�a� ^��Bt�2@-�nUHm�초��DH'�[(#�Mw���W�gn]e�i\%E�Q�1Z�R�??��ܣŘ�'��#�W�2X8��V����{0{N��t�|�E8�(�+����P��#5 Ư��D�wg�d�-y�x6�S���;�<䏢f_�ia!�=��R懟�w�3��������,8&�R�Bc���^�Mw���z1/���|/��u6��^f� 
&3�+!��h�R�� �K��J`<mlkFq��ϵ��Y�s��	��N�a4�5���fDg���	�3z������s��XG���ý��Jѹ�����sG�4�d��X�4�����ts���m|�����i*�i�RB��3*ƾc�����H�xry��yz$By��eg�w���0�BO�T0&�(��XJ�R���+C��Y����.�g�VA2�+��"�;�"/�>�!��~���&p�GD�қ�b�̷�V�M-��RN��SD��r�UzU�-^���9���7"�Tdi+�Tc�Һ�_�L�$ʃD2n-H|�����Ķ����tn�U���ko� �o�g(JC��6��H�aMe�'	��N���5��A��d�"e��ɑ�F`�����tS/Y��4o�z��g8���3s�^�Z(E�X�G��&6⤫��[�~�o���u��a��x�.x�����$_Z�Z��k��ss�u��VHAD��� *�̣�U��1p��o���(�t[ޢ�|�d}���)�/�tN��dW1���I�p��Uin��U���PH������=i?�33;�ǎ؏<�!��T:�	zҤ��J�|���޸�eX[��Ĩ�3mOX�)kZ9�˺ߍ��&��1ָ[��Z���������T����׈k���U���N	�x�}��X�W���#L�kNm���A�-9w0�M>���ww�B5�m����Bm�v\!�x������<�Ex�ʑ�r�ʬy�c!�����P��݁$���d{��W� �����4~-F�����CA�����F����*�5X;3���G��T�q��V��a��7�SV��e���ൢ:�.���C�����U�!�.�yD��.��ѧsMN��h�5����T֙�����������8eN���e(�Ss;�;D�!ļ�[�c���{+�N���{��OB��׋��ɊX�p;p]x��.��g��#�e	r}!�^��w�V��[�*qW�[�B��X��t+��`��DDmE�B��=���4�g{�F*:��x���g>�jV�U<K�k��y$ǀV;��Э����MlB�*1/�F� ��Q7��;����b��������
.6�h"��~[~���6�JN7CzO���_�O��k:{���X��}d'/C����� <�ZEh�CN;��O��d%���`��������A��I�²�Zr��B�����譯,IG8���fO�|iץ��/RoV��|��h��9�1HTl�__�T��n滬a@4�E��^�K�� ��e����:*��;�I��E6��p c1���
�@�Ap];lM6&7�dX�A��q<ʛ�����D�3��#�k�%���1E�BQ�[�9�z� ��uSW�z�O4Te.����p����f/���v�=���;y	��a��mu��?T,J��dk����e��eú!w ���
|J� �C�d(�~ވ�|x9���aN(�G��#�C�ܰ�Tʰ{��:�8_��OGb�{���PD��è%!�g��A�Љ���E�P$}yO6˸S��ޟNP�"XD/�\�Oϛ����q����"
�8�I��-]���/)q�6����l�ҫ�[�Jd�J��/�!���[�I12��P!f��WDy�ꕌ���2�#���7ڈi�/����C�g�LS��6��r+����fu"�� �s�*�#b),��*��ʐ�
l`
�Ul�9=���l������~* ��ZI��m�?�G'=1�������5�2
�Z���u���Mg�	�`V�����7�����02�=?4��8���Vܟ9A~���}vB뼺T�o�;
{�v���Ϋ3p8't��Qۨ�z�������z�������3�A�zW31X���̪,D����q�n�ǀ�.p�5�rm���M6�l1�	�B���|�JO��+
�6i��s����<1��!qg�c��b�n�[Z��1�b��'��/���s0��+q��F��s�Na)R��2_�h�l�T���iU�p�4m�ȰYj�ܣ�)(�#
f(|�� ��[ϛ؎��
�Pۗ�HY��9}��J͹Y�~���>�/����v<�Ka��y&��L})U�f�~O��Jm	����:"��.sv�R(1��{-x	 u�L5v;���(��GR�]�溒dB���J�$��c ���m�� �&ưu��]	��+�{�[7��7 �,��:�¸V��A/�-0K�~H��>#��u���{F����[) ~�����9�=A�p���1�� $�t
G۾I�����/<��?�SY�Ш�'�
��(c{�i{DyH�Ջ��LĴ�R�W�Q�ٯ�ta�����V����4�V�OLU�����1�$�ʡ[��6� ?0�aj��.�uZ.��q�9Z���𠗄Gp^(`W؏�*���V�ڦ���@A �"�ҨdshB�