��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��XMXl�M�x��ֈ�$ɜ�A�_�4%�Y0uȈڄ�(��_�f4�f�!w��>��z�
��B4�]^�"����	]������xp9��Hyem��k�¿�ջ�U�#�}��[E��4�?w��N�#�H���5�0�j" 2����9�ϺE�n�!\��*�wo}�\�輜��n#l�'��6HKìԀ� ��҆�*y�O���������¸d-���KAh��~	I�����*B�%��W��(�ZX��"Z��M���2�5傠���,�&�dhD3J���]رq�$
�\�6��ڳA����$Hdgż���6l��X�Q�7��lP�!C�P��cx�,^���=��ָ[zJO� H $�
9f�zP���.��^-��ɝ�NM�'J�kJ���~�=Bb~ӎ���W������Y&_P�Ē����GC������I�N�6/91 o�x��G�
Wr<0�?��T�2��Ef��^���J��:{����!B��C
AW{iJ�g4Ѯ$���-�2���X`%�W�h���T�?�M����m��̱�
��iކF�~E^�TV;��D���<�6n�Y�㞝��6�T��Ξ�Op�S������lil�<u]����pC`�pkr�6�݆gNw1��cW^W�(X����C���%Qw��-M	q�z2g` �"���'�n���ŀ,��5G.�&9�W��<��Y�c��焔�ѺN[֥��I5b�@��\v]B�!�L�\���^��Ne�]9�?Қ��3��d�\*\g[�^ �%V!���z��&�{�5%��
��� S{�E0���5y*i�����!�8}�(�݇a���Ս^�A^�]��>����L���y�TMJ	M$ڔ��� y��Ȓ���Si��D+�?�4�r+,3��9�����������qq�ub8j�i�	h Қ��XH^��Ͱ۫Iٓ��d�C/�#-�\仩g@Y`�	���3�#�;4��-?�a��gW����!47AE�-��c9�<�F��Ze툂�k(<�i�����%\��G�S>y�v`.k[�QO'CN������Y��G�PF�-`ݡ��>e{�d�I��W����us���hp.��ҁm_y ����G�����u:D�RR �{t�4�ڷ0�.6�c}�o\�ğ��čZj��k&�se��d]sQ^mE�R��V8�s1%��WErw6�y�t�d�����7�[0��ϋۨ��9�D�9�ѝ9��B�����f׷4��.]�;sV�%MT�R��o2����O�����r�>%eC�S��j�=1����ԙ���?L↡�x�ŋ�L&Qě+̓��~��@� ]P����!�'��y���򝅓|��N�~j!؎dhv6��P&���ۨ`���Yj�uP��-�K4҆Lr�gPP���o�%^��Kѿ(�BD���0MF�u��w��$� ��8W�f�Wa^UNMl	Tk�4%,O,�o���UA��q�kb�Ûn����8�?QlՐJ	'M�Ӯ�Eòj��'�%A_fޯ��̼�������3>l�@��Y����_U����x$q3V��I���P
������I�[��:H�AX�j^ij��a��2At�:��+}B����:�k��L��rv�qs�o��Vd��0G*���退����y���YQIgu�~�)�uL%�C�3E�~��ϴf��V=+z�C��d�1��t�.&�����ӧ9����j�"�4=k�ق�;r���*)�'T�
�1Ŕ2&b����g��ƆGdNT�:�����A�]�}.&�!�$��A�8��[��OG���p��`��i	������^k��8K�_�fΑ h����m#ao)�Š$ Jn<��iޓ��ŞGY;��nw�tH�sWC��q�8i[��Q���%�� �::�lGs|�M�:��*�E<wNN^��iBf�{��9����)3%��]8���o[�e�"����3��:�_0$����y:��I�N���:k��	�1)���I�̕+�`5��k
��K�=�6_ ���0��]h֊�=�C3J��)�*�#|������r5T� �j��/�D5b3�|�<��J����ʷ�c1����tc?�3dB]e��u`_b֛�ť%���Y�6��uK�}8-|�8^��D"�>LW���4��I�^2LSا�Z��p9Q�F:�xȼ.�w��Bѱ�vxN�=���]��ُ���=�\�:�F�v�Oe��& Y.�+ؘ$��a�`�`p�Vgmk���Ө�Z!r�V��L�JMxp��C_p��B�$7[�'\&�)�Ոv�q!�Wݿ����s_�X��@' b�c>���,�o�b\N�cA����ޚ�"Y_��F�u�~(:�&�P���D|�/"�i}���KR�n�������aF���Ya!J0�U:V^�cirj�!P��$}}�"vt�0�x!p؁�(���a]u%A�~����yQ��I�)�8�k����K_�;5Eq��U�	���ga�n��{o$�]�O	u��Sg	�ǳ��`	���_��N��ڜ��+�;�b��#�;*��Q<-a�B�;��"�iI��[U9}�Pv�5V?�̦8�F�J���о-i?d��>�(��CoY�8�ׯ��-�ui96#�����v�4�ծ�h���L�\�0����^%/ԯP��)U�� y�ɝR{X����̈́VyH�����:໦שK�Q�����kI$�"��g�)Q<��R�IG���ɃOT=�GI������h9�֘��r��������D�(�Ce�P�
��	X��qㄊ�-h��X����D*ZS��Xok��H)?��ck��H���x�u�5.��œ6p������pr4:6�<����u�T$k���/o��2�'�.���PRoJ�4�������쭗Q���D�N-���ng'�����xS��Fh�%�������d4V!.Q*�~�����;�����' D������PGD���Oǯ�Nb�k9�s�������5��,C_��#ծ�����.���M�#��y���E'�rN�.r�B�0�B�b\ha��U2�H�]	�]z��Y'�7O�鲀nI� ��`���K�{P��5��n,���{�D��W��Uڕ����d�W����[�e ��d��Z�p�U��.4	@Cj}a� �*��v8�|=�x��ʼ�X���Ǿ8��H}e���E���>��K��χ��Z;B�ȸ�Mc�oZ����nG_��=�/|uK}QB����.0e|._�Ae�S��F�a���eF2�L5��/�F%Q����*�-�!�����CJŝ-�s��نq�U��$�VS_�
&�Ja�Tt� {�	���Nu�k�,�b4��ﶲYb�Ѥ�0/���W�����A�)]�w��4��a��$��5t��b���q��Q�� �s��&UH�-�G�9f��m�����Ľ����|�@\��c���;�1�Yh«�H�M�L���4���HǕ��gj
�x�+,��𼎾���i(�r�Z9�0=.�V%��a/)Q�Sa�8s[
�ͷ6v9?�[v.N�=wc�#��H�E|%��6�TVj���hTy�i	8g�]�_���LxJL_-y��Kp����T�����ރ������2g;�WA��k�")�G�Bn;�߀���B��𩹂�oA��c�O�b���>�ڡ�"	#
��0x�j���0�aӅ�i����lJ{���k�&��2x��"�ڭ�Yo�ۢ_���Ni�h���9��_��U��ɦ��ˣ�1H���7D ������-�Y&Ga���g��B��+�5u�}�މ�Q�R�V�����ĕ�إ��T~;c7�Q��-��GfY���4g���j�8�-(�軗O쐡��y"�3"�@^[�=Zf�va@Q��A�4��jƯHt��Q��/F��6��Nb���Z^�I�Mɭ����=L�J=���Wq�_��0J����͎�9�p�f-z��W�k����f���n��{k���>���G���<ox����l�D� �̊���E�ۑ���ײ<��^d�3*[�2Z��AR�]E�M�O	?�,�N��<a���"��b~ӣ7�Ƥ�U�MeF|�������A(I�2��7��a��a�conu��o�R�kK�lk�ڝ�P(�Gv����Z���U֣�e�T�(��ƬBn��I�x���3zȣg���̀s�cC�0Ȇ+-��u�����h����0���a[�������H>A��G��h��+�'�`���ZeV�E�x�x�����x-�=��w��#z?/�C<�};A��������a[���~�q<cs���۞"��$ S�Ү��I��8��jwЈ�H���£ĢH�Ϸʊg��繉����E
���.�����PAH��]B~.q>�	8�3A��P�Y�ׂ��*^ɠ�~z݈2��~�������F����E*�d�����2����ϕ8;�ZFU0��z�Rdq�CȊ�a��W���:�c�̯K�ީ�8k���_���~�;�z��ɮ%�aZ��ք�q�8��� ��~/&PR��Z�޽b-=W��;�TK�z�)+�^�E�]4?8�t��!~~��޴�^�H�+�>k1��N+�G���!�u�[v�Ss�7��.����_-9������-�^���=�8}#��J�]B�C��j�Q��d-�|8,��=�k��-5xǢހI0z�yʞSb���P�%�>��H�|���!ĺ��D�t�É��4/^�\p<��8-�/��;;�1Ƚj�}���T�2�r*�ۢ�@&a�o���"I���Z������B��.u�웡�~S��Ϥ�6F�b4?!�}3��|N����n��5����c�K:���Z3.�:G�7����=�@r���{�P�>�����z�u�P2�À�<V��l�~�Q��E��?Ј�R��MU@�.ny�cx�	�;��#�� �P!�*XBpt� �p�w{���D0��G���=���`!}Y���Cm�6#ž��?�+u2`����3�8G<> ���5��Πv�ڧ3�7�X��|@f|�u�v7���^߳U��}���.�h������-��3U_���K%g@��阜i�&	����`y\J?� ���y`��d)(7��HHA��"K������kylg<Z:�������4�?� 9�7��:%�Wp3&ƽ���-��]μ�m$��X#4l��˸{!
��,��S%E�����G��e�:`��`�����9V���0�E�,�3�O��k.(�w�?�n*�ob��'��ۙ64`,�V����N�z-�G�6j#q�YO	����0	�\]��)3.~0*͠�D�l��Z'�p͘*d�S�����)�߅7���ǭ�R�R��\��L�e�#��%��l�Q
��ݜ3�C�|X�DU���V�9*�����a�e�j������x#���-�̗29���?wF����8bFB]��.�3W�6d0�hpgd[��7�ǋ�s������� �s$��r)�S8�jt�#5�H�X��GM�œ*m�vQ��쾖w�(bk/_`��5[rR�t�׳�`�덶;�r�fY�ֶ&�Zo)����D˧�UsD����DsB�n��xRXî�W�>1-��'�5�'��F����<h�4�����-��/neT�M�����X֪J���j�^۫?�ua���m2��� }D���d3/����M�Q���S���ުϫ����%�W��TtǸ<qG��)o�@�ǁ� O/dV���"�=�5�������ژY°�.
��Ev�;�������`L#��>��i�~ח�r5�|{�s*%�U�ҙo�#4�Ъa��5p��t�߸��f�se[���
~�S��qmҠ�?�o��}`oǊs��ͅF8h��/SZ������-��mԸ� �Q��y��|qO�%����(lՁ]�R}Hz�>�.�F�"Yr���Yg5���� !3�aªaMSE_����EJїE݊���!"p��u����5X�Q?�Q��[eD��\:����G���1��f�5�`�-*]�M,X�0Y���"�r�,k��J���� x��	{�.�Zc�F���j=��3jۯ[��X�?0�+!��5�쓢�����w��6",٫+� :5��ߊ�)��7���'�?&W<#;�n��+;Q0^'?���&�"���f��3�I���5�w��XIN�-�_4b�1s+h��#�3���XB�.��2k�(Iw���If#[�4*���X���]1�ˊ�~���"K�%V<�n��S�n���ru���=P;rR�PP[=Ahu*<�~�_�ߩ��z�C2Y��g��Љk�6�	�#K�NY����&��NY���3�c.�8���ϔ����` ��'�g%�Rc?�_���N�����-��=�rXN�"2�v���	�yT[�P�ъh Wˑ��9��y��=���J2"���o�8��.<�zy �ұ�rI����8�-�>½*Bb\+tp�Pn�ц�v�('�k�T�w���>R�Y���"�c��	0S�ek�����p5-q
�+d����*v��N͕�7�r�ک_L&)`aG"���лA$�mwg�ag꽫i�l�c�+���`�"e\�"x���»7H�7�'u��<r����Ppv�?i��ݴ'[C=����|�`TwDe]Wx7��u#�l�lo��#����^"���GO�.�6��*��]�P�o�PwDЫZ�W��tB�`�%ܣ5Z�"UR!�TOȂ���c������e���;�Ѡ���&������\��Rqf��.uvun����윒�DӨ{0\~��鑭��xs/�=c��yF_%�p�n��0,0��e�{E̾��@���]}�XaU��F���K:�\���	T�A�bp�2��#�I*Y����t�GxbK ��si��ZK�Vj5\5��]�4ֵ��$�t����@3���A�MW�e~b�����1W�����)
�~���^�� �>�#�
*���KE������A[��вŝ��������3��������}^X�X�m.쌵�.,#��<;5�L'*q$��N��U������S�3��u(��gx�j1AX�NCҦ:瞗��U��^lD�o��X0'��� =K�$�>�� ^� `Yn)<I��U~�����Ӛ�tI.���7L�S�G7��ep	/|����C�� Mk���}w�yLM�Yg���e�b�P�V�]r���Qg�R2Ey0��J�;]��'(���������yBɂq:�a��.�5֟��e�}?��N|�"8�^����j.zK�/ə�����/T����w.��~6�!�/����>��C,��>M҅G���,N�z_��o+@I:��N���HJ��]�Vg��`��Ehw7g���.86�-0�0�����|��ϵ��; ����#� JP�?1��ۖ���е����?D`׸��7�no���/l<���Ø.��y��5<e�@tw8�R.�z��u/�#f�(��!aZ� I}����.��F& ��ญS9M�N�� ��	�9�)3Q�:�o�����V�(ur�Ft7��$�"'�H�2F���-RM�m�o�,mhA'��㨽����!���=�rV=�W�p>U��:7sWIGb���l��| �z/���;�$i-W������'��~i���趑x�2�=����Y>���K��W�	����ˈQ;9���>m�s�bv�.A��f�� ����,�����<�g���DΑx`	ӭ����@��9�2�1&�ٖ�&jx� �P���
a���w�P�^�jY�	&oO�o�:C��c�u�f��ך�mf#�6�x�?d�0�����a�&�zx��B����Wr�"^�ㆁ@�� �@�x���+�bQ����3e꫷�Tq��vY�=p��03?B+R,���;���G�;���Ǥ�@���k�4u�y�8d჻�$~W!��i����%�]H]�MB����h����y���HB���"m/�,�ybe�(���)��X��{hE�ԉ�7? $�/�}Hŗ�ł�� r���=T
�O��4�3L_�?]�y\�y^��Z��;.�����}S}�jE��w@��%F?@D��,�cvZ���[QG���Cq�W�W6O��F2���}�gE��uy�?�-'a�XWM�k���s/��Yh(�\���߆���|7��!m������p̚KvM����;�Y�O�#�����"�Ѯ����w�@���$1��!2��9槷ۃ�q�����jW'{i��o�!;>�L�2-�U�H��eGJ�R.D��cN��'�p=���R7��'T�DA'�m������:H	�
��H�x��[:�A�`r�m2�_HuD��c��l���SW��Gt��Mk$����d��}�-��7�b�^?#b��\A����sIs���%¬�cLL`�}A׶�6�:
�t<�V��Ӡ(�ڼW��u6۠����ԛ�>S�J����&���3�k^Am5t��L�߿4����C�?��!�yP����o��p �$�g���N�'ֶ����ԊM��L�Rݤ~Y3�k��^꩝��l>�`�0�'ʆ0t.�<���-�ӎ��E���v߁��ցAR_�oӅ Ŭ��7
��t���D!ŀ*b#�졎A1����	WNܗ�S#�2�'Fd���/��/J}���rH*!����i�(��o��E��z�s�ƅ𧦿�w��I�o�� �6Іǵ�J��C���2
h+k4l��H�`�.�kTAi�|����j�"&T���I���j[�Rϑ9�{Q�	�iI f �V�)�tbL���C]����b8���i=��̏O�FY���LbbIK�n�gMn���@��� � 8�	*�w$�RZ���ք�'��Os�I���K�6�ڟ5���y��T�7C	���X��%ks��.�x�6?M�,Ю;ߩOW�����@Q9�f}�̫,��[9�k+�@\--��N�if�D?&��J����i�ɣ��;j����^�a�r�T@	E�Ķ����r3Z��u<e�dD�y<���
� *�EƔ���Oů�hQ���P�<vكb9�acOe��ǔ`c�k�9Fidc���f)���!ۋz7 )�~�}����[oY�9)z�2Z�+6��L�4�6�}dx�eb#��l�F;��{T7���Z�I��=1��/}�ć�r8̶��<Zv���L� �FU�<eyI�HHw��"#��e�\��[:Y7��MӛJL�G8H�i3�=��"�*��͉���������"
��M�r���"�A�j9(�/3L�����͹s����+��q�(���0��]i��w�-I�U6`��-���Ŏ��R�ы@��wI�w.;:n�#�t$�@.^<�\�� ވX���'>-�H{"T��Nx�z��DaC��������)����f�_���g��.KU`9Bk�?�V��q��P�����ם��noO[�QH�e��yyl�
���|n ͢�l�\Om'�C!f$���@���i+G��Z0���N�p����[!��{⧷$~r�t��k��$[rg9�����B��U�@N9Tϲ�Q��ר&����m�K}_ɧvL|��B�/�_*-���Ր� e0h�e 뀅������a퀛w0�z�]ȼ/��$�S����썅��eR���!�!>�H��Ⱥ�ڱ�e��'Ϭ*B4�3B�d��P�B�%6�=�?����wrT�UE8�3MC�-�����t3T���R'��G��ú�~�m�@l��I:��F=��t�v|�7��z��P1�~HW�uP�Vĸ�L���U��}���]��u@h��g�SZ��C3���A�l�)9�-8G�
�P�՟�9S�����qs���.�)fHW�>��`��@��p�ê;Gp��A�=�����P���Oe�xiXj�K���������Ŧ��'�L����r`g3�bṨ�F+s/B�ۥVD����|��������	';a�ӎ%�������
�:��\�k��L�����Ŧ�]?Il��C�eB��؎C7����i�&>c��G��1�;8��"�\a��^�h��
ZK�|H^ln���[_q���"����cp�نj�.�d��1W�g��A�O��ܱ�aY�xD�6N��)sT�r�힢��I��������q�ߢ"�.)�P�A�YKgj@r|��ׅi ?y4����\�"Bz�{��^d8p��[=�<���%�d.�/g�;!hs`�� ����S�B�FQ�g��_�b�k��	⪊@(�p>� I�����l��'�����C~�guW��� �{�_�h@�2e�����.�B4y<dK���h�A[� ��R#�uv�U�����<vaǅ�L���V;�~�f
p<Ԛ,꛵���BZ�/����0g����0+oDW
�R8�.����1�T]Η�Q�mi��k��1�AG=�����r`7tFPo��q<C}�i�Tg8U �m�ƴ�Q+�����޲�OiS�X��nZ&�B��}j�wW燶���̕��\&L%�%�R��u����B����+��5;�P�@�]+x��h�C���r��A3��1X�}nq�g�� � ��9J/^!J����4J��k�у�ݜk���t�Nj_b�8����KΣ>`j	�C��6�� ��׽��i~�>�����X#>+g�^7BB+y��M[*��E�έNg�֍{�����ҩu��L|o�=��ɬ��6�S��R#��|n���۴��ܞ�Md��i�|��V��5�ENE���7'��^'����?%�CS�����:0�RDa��-}��v�0K��t4P�1�`�$Z�C�E�Tn��m�o�����+{@u�����e �F`��I��N�T��(�nɆQ�^���ɟ\�9���q%�3U2�����7gV<2m�&/��X����/�о������O�/������'��6ؕAv;��D�3��uTԹ �@��wr6���
�uo0�o��!�Y���U ݘ���K� -?��ʈ_�U&�Wm�CQ�> �Ԍe8���R�O���A�U�����b��2R�۱��z�u��;�H�����i��_�cc_u͝)�	T��u43������uF=9y����~��*E�)wS�]��8x��׋n��6�L(g����r��Vt�)j|�e��y:N 5OSA�u��UqH�b��S�	��m?�V�� ���TFŧW����_i��\����[�,�,թ����J%~����+I����N�&���9�����Q?A�hW�i�=��F����d�9-�S���Q2�|��s���R�#���i\��h�V�Hv��`�ܼL�8��-�M>�<�@�U�G���u���9ʹ!��<���cDF	 _�"X9w��^��w_T�.)��!X�S� y�OǱ&4H���"��a~:��|�l�V�`�����l��)58�`x}�-X�K�lh�J�ߪD6�T�Q���yY#j�w�����3�6��z4�������0N��Ca����T��sB�k�|���l{'[u�=�B7�N� �i�)��F����>k��wZ��Z�#$5ob�9�&�]����G����CQcp2B�L8a~��� �|v�U�YW��
��v!5��t��(��n	ӣ��^�
���˞ .�Vr<o�@�]T~�$��1KA*���I{\̜�?�:�l��O�o]���7�j��0�"23��1���7qIf(t�@�g��V�����F�ur#1K|�Bz�� \9o���{��wDq1r�'���Op�	�ԣS9;u+`'\��d���� �����(�ۏ�i@�u�Z<���p��4�|V�	S��&��6�OIu��z�{�d��뺄��ݣ$u]�P�<
ƹ��d�pUԃٮ�Paq�nX��J��� ��K�9lMn�����0���zC������Y� ��O����5����"+l�6�N���>��Lz�[�b�^a@0�lyd�Fo'_�r >�{B+G����WI0����;�f�>���NdiL��a�c��:	T$���Dr� C�U��1���tI�闽�Jء�'�ț��x#"zb� �R2�U�{
���ڬ���������I~�碊6�$�9
�P��r^�����B�ɾ���82ܖ��;�%�as���ҧ]ѕZ�#OO[c�"R_nn��dtw���Q��ߎ5,Z|�n�0�#4BO�C{���Bt�(���Z��J"�8��<��r>!�wڜ��s��ǚnT;w!m�|��f^�Z�$i*!-��i��}�kЌ��7١�[�R��	���Lؙ�O�o�$���h�[Z	���\?߼)c���$}����.s$n�`��|�i�m�3r�	$Y����G:~���_6��P�V́���2��6m�o{qg�D=���G*�g�+?~���C��'�;-�"b�@��hq���=OKun�*p�C
� {�A�	{���d�ARp��Y�ן]$��y`P�4�6 �I��4�m@j�𲫉&&��ד�3�)T+��Q�E$���P�C����Ҳ��|)�i�STi�T�&D[�[.@���)�y�L���73�h=t���8�&�e#���:�""�W$\�9y����0�C�#���;uY.]������