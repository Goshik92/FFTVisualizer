��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>�� �F9!�/_g�T@_hm/a3^��(#z�dZ�E�����v�h��|���-�>����w,.��N����9Z�S�p�ւr�p^������[�G�C-�Dʩ/�Pm��[���h�L��,����>�&�_��ĴN��E?�IC����z�kxC�e�$rC�H0>o���_�?�����i�Ŧ�.�"��?b^��=��[ԋ1���&��	��,2��s�M�L3���Oӏh-|�Κͧ��#a���v(0U����l~!��G����}��؞��tY��һ/S4���>�~�ʊ� x0�L(,�,���jp�^�)�Z��C��r�G�&cn��
5�뙢�#��Q���ؖ"M6���M%G(N��q܊��8�*7}��y_�J���!�&ȷʗ_N�J2�I:!����OzD:�f�,��!�<�4 6�!l�(C�]���=�+1�E>0�κ�1��=�oW��ӓ�V��$�&I���z��a���>s�t�m�X��������TX}8��o���.l���G0�Re�:|a+&�f��Ѡ���م�vѠ%&]d,^�Ú�[��x$ %e�ݒr򑻫N<�-���yO*u�ѻ�qr����p�y�"�Y����OF��ĭ
�_��.8^����a���M�q#
�����F�g��GA�\C���H�Q��ߎ3{�WC�0J��z�]�ጒZڬx�RωSE[�f&�����}�Y 	Ł�E{J��!��x�\�J��ɩ}�nL��,�|����Q��!,���C��n�W8u�Թ6�^����b�7tfյ�GS�Yj������;���u>�<s�%���]S�?\W�ZFDK�����:�����D����w���0�j�v������9�ނ[�H�d'a��@k!���Q�}v�I�uмs@SY� OP���}�>Rw���p�A��[4wR��?r��B�&$8�@)�=$���Ez¯�Z�y	����y�8��st��D����UtǰXϋ쏫9#J�2�B'���dV�S�Èy�G����QU�W���"a��w'�l�]�R��g��.�TMT�#n��C�
̞0H��'�^��`Q�"�{7�}���bZ��s�
�I_X|�g�~R���C���_��.cp�ہ;��wɷ�hQ���m����	u� ��}؜۱S�ʵUbU�ܭ��'�������^�gᶡ�Rb�G�2=�� "Bm-�ؒ%����v ���JG�؈4�Ў��D;ƴw`�������S�&�B�-<���/�ԗ�]/@�h�䯔��� �yO��d�0e�E�����N������g�jwU�7�q��]0����O8�i��$\�(� 
%\�Z�%��S�Q�m�!#x ��vio@�5�9����B�B�[�YN��������u:d�pw��R�S���`FS�?%cf΋�X���;B/��*�z��9�� A� 5��*U"�z�ȗ��ai7�0��ٚ�);�$?��mh�ۯSZ�����;���&�xr�����:�vF�%ш��/��S��jML�K�0���~���۝���J�+Aq|�9{ Kk�;)F�$y"�d��r��z}���
����\G~���t7ԓ�t[qN�j�8Q��D#Α�H�3LO�L�V~�6f�T��SP�����Ic���ONqjO#��/dܣ-�g�bN`��D�	)*╱J����Hqf�{��Ұ����2����WLPZ� =M���d������@�B�� ���є�Y<M�̂&��T ӮBA��F2
���c$��3�u ��+�$��Uy!����y���"zD*��������`�Nl�P�ݜ)��R�	�� r�'��Gk�d0H��E&���U�O+��vtO�����994CH�$�oe�Р ��>�7f���N��6j��e�'�&�5���w��БQ���^m&�<(P����z��&�f}�� # �]#�3+���`�$By]c��qLO_�`�p�_���$�e9qJ�zD�����h�$T|�#���A�k����N�4��d���AlR!`;�t��ۧ��93���@M�/xWk��J��I9(�5��a�m�=�}�B�IXQ��h���cݍ�a��y�m�2㲅��qo����2V}��}������BJ=�$;�(��0��}LL{@���] �x�Xp�9��x��C���h;��PUr�n{����y�d�?y�E47Chai��(��PD=��O?�czY1{Ye�K�����A�n�J�T̔	Q�[d5k� k�*('�0�#Vk�x,ME���)t�5k*�A-L�,髙�q���ْ�Ƙ�cJI-T��a�I�������4O�JZH"�8I���=�P����:`��yF� q(��8��O�-�2 �M��y�FM�Mr�/P�y�����X�5�v���4VgH�jhga��1���Αkz���S����9oRM��v��G�6UR���{��i���BV(�$+Ȉ[�g��$������ �Z+CP��˧�E?8�݀��C)�8�@�!�r2;�6�RmR�`#�u� ��¨�"�a�Jl�o�lq�h0�\�=�jr�0�*�I	��IĆ�4��ѕ�/���yO��X�BI�MUj������o��Ԁao�*�N��{Xr�%�ٸ�p�=�Ѝ-�s3�1������K�h�*C>�T�����rI�Q�Ri�[(�
Ėl��th���T��C�U]'"���#�����{70e�Z5������6w�1����Q�D�uw�bF6)Қ}�J������Mг{�=EK���m�6]���bY�Q�*���[~qǈG���,瑴pn���vw\T�Q�;��������ٟI�w7,�)�Er�3uM���?_��g��~MJ<�x�������aҦ�~%!���:3f]��c�����٭n��<7I�k�}$�1�v�tU%.W���1 9�]`]/�S��%8Vx	T��VBK�|03�-mwu���a���`��Ɔ�iƅ'C���e�"o�~����[�1�ǰ�J1u��s��膎��8�{����� ��cbJ���k����R��l��-�T��W�f2����7���)�M��X���C
I0���+�@�	�lP�*f�?�7�E%�T/����ԇ�Z��\[��z�i�����l����Ӳw>	����(��;\qQ�L`Q���ß��	?ϐ*R��hy=K�� ^+0|I�Co�S��hpT�v����N�y�����1�0R3�~�R)�<�{�^�ٷ�#I���m�� �5�D'!�2�VREgB�0��tj�!�}=��)2H�r�E�EzKe^�Y��`����q�45g�T1���xӵ%F��PU;�E;�굤�f��� ��4�cXV��h ���C���'�&����r�	�E9�Y�e�(c���}�:
����a��MX�2'9���̀*4o���k�恏v}O�E�#k��]�cO*K�pJ�[�k��.�۶���9�x�>�~�r�$�ù�� ,X�l�w��n��^�5U�>�'!i�o�T�nF�����IK��^���Q ���Sy�l ���
z�ȞUе���Z:Wrv�[e�JXo��ՆCZu��\��t���4B��Yn˨�u����?F����e���Tͺs�EdZ_����<}_��6GZ�@=r5+U�P�o(��0����>D��
}��*|�Mʼ�?t#���}�����z�^Ɇ[���j/uG�+���xv��.�gP�2�cLS32�#5��"[��>u%&I�&��u���yKi�Q���߁����.>�V��f��X���%7�"����(�#�������[X�N��0��|�_:}O�R�Y(�y{���7~:C��>�~��!XD�>��}���d��Ȋ�2,è.������`֛a6#��
ͮ�c�
�B���� ����idy�yZ���ucG=�K��]_99)�
Ki;c�m�{��{f;����ݺ�y�隺4�ҏW}rZy��7˿�%��)'<�G�3�H�/h��⤘��=c�=qn���8���=����d�5�$)e�������{I��HA:�ineo����=�Wh#~6M�0|�
zK�I�yv6�
R�4�nD�0MZ�DV�x�ץ�.9`$[�^�ax�u���az�	< g_y8�tE�V�E�Y��J�`���1^��D� �����K	���N/�aJaKdϺTJ!۾!`���N?�qPU4B��՟�vd�6�5�,xT���ؽC����cH