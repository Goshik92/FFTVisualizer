��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ��nͳ�R[�ظ�_����Qq���G�]~��\�^�W.Z��ke��X�?�I\�zA@���Y"���a`MBl��$���X���/~%�cg��OU#,��;o�w�F�~�wy�0�Sa��qC�$�_됲��ݗ� ���D��.����v��C��k���<�$J��3��I
����<[�P�}&ʁ_m3�P{�
A���-X'�H4Eml�}-���i���[�f�c�:Z��� �B�O�P���c�Z���S����[_F�|=�����{1��ƴ�;���0]N]!a�OIr��"�p\�b�'�YQ�e���&3^��H˜���|��
��t��]�^��ΘM�7r��֗�?miH!nSA(���3e���'�+:AJ�N�al��B;������+֍b���+�ݑ���=ɮ��"�.c�%�zpM��{D �p��Ӥ�������!A(W�����]���AA8D� ~�F���S�� N�e��~󂢚v?̓�H�@EM� ��ݦ�c�Lc���v�������N ȸ�iP|�M�	0�����L����J)�0ɽ����X7IL����"c�'�m� O��ݘ �V�T�bӮ����Qx���2۩ⅺtH��*g�ڼ0�S�~���C4��+=�ke�ŋ��3�g�����7f�;$���t�ث�8��*Y�Ӥ��b�\�>%&;=��"|���i� �x� ɹ֒�f����ʺ~2Rs��kмK��V� 𲕨`�oX!�PEv�����L����Qfٙ��6���뼆TB���D����lŢ�㦏R���TJBl84]a���\p��+�L"�8���+\�:���z^�5]�_�^���6�Q!S�p\	� L��ӯ�w(e~��)!w���7�����¬�R���u��w��>B.�mfrN���};Ɵ�ן��D���[C"�Ϧ�k>��g�����0=�w��ӉgԬ�3�5�x���*�{Pg(�Z'���(|ߕ�&�P��Ie.g��̋,;�'����*��]�%�ZW:H�W61�_jN�T��T_>>�|��ˡ�l
��jX��t�{Y�#�]v����h��|{v}ų������Y!�����jb��۳��\>(�K8�%$n�&�V��s��BrN�q����ԪY�t��n�F�ޑ�T>e<���H��,���)�7�����I�ۡ���3t�1T��h����G)9d�c��1t�C����4?>��J�[G����p��쇑�f����~��=#vf�VXk��ܺ�P5�|T�� PS�[�-�:�i���>��3��R�{G�Й�ZOR��#`�h҆�A('*E���~�xA�Jo��M���=�J�����u
�����?�q.�[e�{e~߆�,E�4@\��Z�ӿ|U&@��}7K&.����Ć�]����ʀع��>Z��Jɫ�-j׹���d����Ǻ��V%)|j������U�җ)��
#HվU�
 ���5�r@��d��M�W�yJ[^씥F∇��SH|\��}��>��YM�EdlҥЕ�)�a�&�@U�v��~�r�P��;�>�=�d��I��~�d	)��\�P)�`F�g:� ��
�24�d?����Գdܯ�����5��st���RD;C�R��^��s�C�y�\��* �Q8&�'Pl�\�C�kD]Èu�����#v�c���)�<Zt��zJ�c��������W�	�)<]8�q�y8��>O��J�,9�ݞ}p���,>Rlkf��(:bq#O��ض�ۭDn��x��n�/����cG�9��d���D��yӉ#�=]�
�3+*�H�G�]�����~��#5z�u��:*S�{Ҩ�h�ѧ�㍜l���i��,��&��	�/$��pf-��۩i|i�A�h.u >������5b0�m6b���Z�! /�6����}�\�����ў�@n���
&�Q�\�f�W謁inc:
��}*����[�)Me9�����?{�%4�6Lp�v#p.N�P
͉��E7C���]@���9-�"x��@t��#�P;���VV3:H�}�-#P�|se6��O=����F���t�G��c�Q�>���ڵ?�:1�2��˚&�;�QӰ��3Q*"y��Ꜩ\Q�c��?6E�߷n�؉ b�ZΑ�5��kZ�y����x�!�	J�a�W��$�u|�ֲ������.<li}Uu�� >%#������'~��G���8�(��^:�UDq��1O��"��?�'x���\��b'�[au"�i!@=���b
	/:�`�V�:���vx��s�)Hwl�I��?�x�;�a���,	�3� [���O9�D�e�&]J����j6�֘���)����Ao^���Wÿ�Q��u|�Ɨx��!z}�d�ܥ���}��c�\|F��?:�}Յ���#�9�D�J�h��?c�.��Xj��b��*3T����@��ۿ��9�8'�`}��À����h�RT�����䔈�okzzj��'0�	�����L�@~:�B�6ÀWIA�ˠ�ᖷ��!E0���iMʒ뭑�Y�_l.JLv���j7�hgg���Ń�5N��8~���d�Cە��e�ht$�i���j"IB�2N��Ƨ��`R������X�u�7�?���Ƈ'A�@Z���NY�s{��������7D���@q@OLK����U�Q%h6��-�F��zumcL��6&U�[X�uH��n.�\�3.���
�.�i>M؛.V�IIm�=H�CECKh���>����ׁ��jج��F��6TX��ʲ1f�������"m-XB��+���	UL��7�5*��.���aF|�L97�J�E����#�����g��A�ģGu�T`���^����>��B�K3�HC�@Lñ�;�����hǹr��0�M���C��\OR�۞�ޔ�%��i�zudFz���~�h�Xw�}�K��u����.�jW>=�,�\����e˶U�8�2Y���u�*1�K��Q=�t�-�k$x�����������,���eJÂ�5-������z���\�I�)ک�ٶ�G~d�3C�d���b�3	z�Y,z��'6���੄�B�q�A����P�$�CR)�3x�e$�PM����y|?P"�*u ���[��f2����x���� �=��p�%߿���h
�raMY�/g2N!�	��c��x�k�V
����N�F��.A#�1<]E��Ĺ'���T���ɡ�rfx��9���<�7�ԺB�t��uݙ��.Y>�6<�ʡ)N�3ys
�g�~�Hqڿ����_�w(�r���nZ��	�� ��Z>�d�?
�
�k�M_,����a���˫�׎�mɾ22������:l��`�NyJ]r�)`��j/`M��1�c@�z�$��ᚓ��������*��"��}�n	]4�D�@�F�u��~QF,���D���q�;>WZ��̍�	��\���|�����`�wp��C�F���Δ1t�'1\��f�8�S�=�x�xwĘ����]�<ө��e�����; �ry��Y��XH��jf�c���*L�Se���u?�;��a`�c����q걀�\��Z8�Y�i���C���2"G�e=�T�õM�?jf[39@F�)�e��:�`	18	�N��B���\��c|M��9�)�i�g���Z.�|�b�8|GW>�Ё�Tbs��Ӷi�6`���ٟbeo�a�a�SgG��^g$�*}{���&��ƣ����AY0�x�s=��Y�0���)�s�wL����y��@�R4R�|v�V�̼,�0z�)#��,�I� 6�2�/�%�d�������?_�
�[%�t��L��<�#�Eȅ�F��R�s�=+-,hln�NҾ3�����u1}e�l6�h���B�c��Z��p�[}��yt�{$��Q̈�q7�"���*�Į>~G��'�|��Z�R�3�_�^B�J����t���M�,h#�n�Z��1Vg�k��c�G @o)�0(�M���(�ױ�����H(�s�hb�VϘ�&\k8my�5�5�|��)9�û���@\6!\J$u��-�,*�V�kx>%�-6I�E��<n)��a� ��M��n���z�gfeDW�#��*A�;l͌^�atVJ�5���=����P�Ckʈ~v�|E�gM�[͇9�����G�1J�f�>l��X��X��X�|��\�c���z�D<"�w�C