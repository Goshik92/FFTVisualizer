��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�*�yo���(�}�ͷ���m��~�D�L�sݚ$&�����s�%��j�t��h��x�mؼ����eF٭���kud�/RMѸcdb�>�{�)@�x��ĎDrŝD�
���q݌�Hm1����L.J�;��%�,ʊ͝$P2#�{Q�(K�F.�48��u�4(`2D�6~�[)�7�e	�3A%V�Zy�����;mj~}x>q�j����� ˉ�����ޡx�QTY��%z�ɤ�E&�\Ʒ����7�f��Ƽ�ہT��?B���|_+:���:�Ua��S�L��T5%���'�3��0[�>!o.����3��i	4��㱨)T��.�e[UTE!�a�,%�5���5ZE����Yw/w���[��?D�Y'�!�}�|����+)�ui8:�N[s�<qXɒ��F��`ׇ��Pi�#� x��S��mK�q��z����]����bw�̬"��b�d)�6�B����N g\Sw����d7D�d��� �RG@-]��� �T!ѷ _��WX�$��EZ��3ܐQ�H���-�SJ�~��iљ;4̝��cB؇�������O��WXO+'�3,ԶA���āzC{A:�.����Y���U�ߧV�L�-;!�{&���*�gi�b�^z�@��6���3}D�But�������e��)������L`~�l�O�����G%I��F��fW�|�J�^�΢*?��m�t1��$�侷�����-��+%�zP��C�"(!�%%����K]�=��8^1����]2��[r����w��焰���W�}]���.�h��2��t�/~p��s��Sgؙ��� �TS�0���l[�ddlFHu��΄Jz�c��U��#��&?���FC �|��d3 3����7dȍ������b�A�`2��E?�^�y���,&�8��A0"�����%�;�$���d����EkJ�F ����U{dK�����bM rVFF�DҒ���˹�P�KWO�4�2�М���M����qg�i��v-�+��Q3xV.��}OGr���ݱ|��~����J�~��%���D6�<����I��H�IFR����>+2/vT���nSD�bi��b�+�60H���L�p���'(�8�VX0죸u����߱��HS�^���>r�76#B����T#��%*����;n��C���h���Emi1���M�c�R�N̡�1aZV0io��B�J}���s�z�O���j�٦�2"9ztci���;.R~����V���C8(�n���9\��Z��_J��+��x2 ,�&��lS������@+���p��d��6��}���?@�f�U!�H��9�W��-�V�K�](k�|�(��3!x�ʹ����6|5��_lf)���t��������u��?h{nuN?N������#�Y�q�=BU�@�x)Ԝ-�/�2ŉq{D��^�g��}��|ߥ{d|��ƌ�Ο��