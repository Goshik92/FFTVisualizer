��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn�5ZD�l[E�ܶy�uri�hn.�-�q���;i%���:�n�ɪˍ�e����.�6UTmB;Y�K$B+1�� դF� �#b�B�;��h�w��i�6PP����<�o:3� p۪&چ꿪Mʱ�0YaLě��I��-��h�.�!Gh�w�x�bYBm���	�2��/����/Ϧ�c��r��t����}�9��>iACU�`���m3��r��p���4�����S ��CļN�P@b������KU��dd6o�pPQV�E��n�5=.-m<��5۝V��9��m���J��fB�E���A��O�q5��H���>�@%mH4A�f8��!_�i-�`��ƬRZ���.�pCe���IVjg.}�8BT.'3��5UW�⽽���]	g���B-��:E�K��V�-N�T/��N�l����e��cyx&�asY�+��t��~����tz`�-�~���4z���9��jjp���q
��]�ubzt��wy�ʷ��%쏀ʡ@ܭu�_�A��%���C�!��$g����5����e�+ت.��K��1���3����ۯ��=�$���)�O7������-肢6:*�>����ri�'�#��X
.i��T6�� �V���� <d22�'N�Mpe^��ㇰg��:ۓ☐msHQt��&]S�D��3�簹��`�� ����Q�<�EI����$g�h����ذ�z�e���=�5��P��	k��+�����u���9�F���:�E%_Ip�k�nc_�eo��s����k�RMh�� ރ�/:B�x];_��f>P:����3O2�Û�ֈ ��	�1Z���>G0�y�� |�%�'���,F�R��,�ݓ�Bb���{�}�^�{UdKa?y���C�����e�TB����}c�=����N��/_$�i�v�ב�A�H�mz�G�*J��Ð��,T֠��T�n�'���-k�^�4E�l'j��B�����+�L�X$�����+�Qci�D5�.s�|�!0V��^,qU�7>�o��Շ+| ��.\毐�8w�H��4?�$�pJ�gqAB4�:V#����c[�xv�Z�w������5�j���N���g���� j�/� :�����Ȼ"48�9���]�����0x���M����A�/�H����B�6�/I�uo�]�N��lNʂm�+�%(���#S����\��5T�ep���~��T�<��lѓ�u�cϽ����䗳~p�-?fJϠn��3�۽��aAI�K�1��|ϻ������W�&���b�|���$/����*�Vot�](*_�ɣ���zJ&�l�\��#P��n�C<Ҹ�<>@Tz��+1����4!r@{��O�[wӼ�O���k��o��D���f�b"�d��;�3�N(Fy���C�8��b��49�?V���s��l,�/섊�3�v�,�q��?�
#F����@�b�`#q�L��4A����_��C�$� �l�����j���  �iu��9���ؾ��L}B}��惬&�q���W�����"q-�Ȏ�8CnUÂ��6�99���CQ���p��7?t8-�œ&����x^)a�V0\�!t��eR�ҿ�Sf<�?�xs�2X�ۙqY�빌�OPW��g����5X�U�G��<,�n�}����_��Ǿ��<	4�zc�sJYax?ʲ����<iE��H���c�v�8h��9��=c��s��y���־�JBB�:^��/�ʰ H�X�[�8֒|[*����_��T9_p�a�?��k��i~��^X�9���U��р��~Ȏ֫����u���&9(nW���~��H�c�B��즹�?�����8k8M+ ����A��;��A욭�D�7Qb�G�q��Bn�9�L��=�ls-RB�p����V&	h�ύ����2��s^}����,�yH���|����ЦQ�����^ŒH���M6��2e-#�����\�u,\/n���eg8W�Z��-�*��+ =^1��!݊u����=|@���B��t�GV�Ҍ7k۵��\j���8��1�H���6�"_,����p���?Hm��Q��c�3��Y]c��_P*Xэ��&z���C�yV�I��Lp٥@l_!%+����A��j�NL���^��<�R);L��lɊ�G�$��l�a�����b�PMkQV��ѬEq&T�����Q����C��[v;���+u����RmU�~7O����}ioA�ZL]�-G6M�¼��
�W}����n��7(NF�	`n�^�\��2@y
��J��Q��۫+�ܑ+y`�E:�u���wKL�-OTa���ڪܟf�,�d��X�G��62sa�\]�����(_�n-��eQ�3'���}2T<o�y^׎� Utcҝ�*��y_&�A��$����e�()8����E��޴t�y1�K<7�1��3�]�+|�)�Lj2�\0!;�t���&�F��� N����e�;U^B	ֶ_8s��b�	����Sk�,�@�� �<2xs�]z�1jY��[g�n�&�_����h�J8ц�|�"�b�mۺ���@^iA�"g��
pB:X�.�q�� �j�&�_k�e!U]ѧ]��x䒟��W���
�����T�=XR�ķ���C+���0�i����l�t���sj���5Zs������(7����҉P�o��J���Vp|�5U�(G(*2櫖y9Lw	=A$l%��8*��H��1u��W��vi�-~�ޏ�Ȑ\h1k�A���n�k��r��V�* �tڮB�@F�(��!멵�*2��q�^I�A=�V�<Pl���r���u���_ �3 b?�Рuc�$��.���}w��n��ɹG���f�W&o*H,�.
�+)�}׸��R�i�V���>�����������{�P��\�m�*�H��j�7ZG�l�<���O�U4��`���M�!
/������^K��^�(���oc���JZ}��䪇��~_�d���?���Wv��a���\�ݏ����!�z�^W�I�	N���/����ε���d��4��P���nU�ۖ�-f#1[d/�"�~|X� � $��~c��-�Ex�M���+b̬�ލ@.H���)�~;�5(DD����wq�R��gG)"�i�*.�ǚ�(%X8�����&@΂Eыy���$a�<�?����Y���5[3^�R�xA�����J�&�P������^�k^�~���	�7w��r�̒Y���5i���	�܎7s�r�S5:���H c͹峟�i�{@m�2%|6Ѣ�c'q#���"b胦�q��k/l3*=��jփ�ǌ��a���uJ%L4z�q�#�Bi�8�h���09"a��������1{��C�'r�dk��J��s��/!J��LB>Ϳ��h�<LD��5���8b���C���R�Z��*�w#K�oTG<�D��i�c1��Ў�sv�Qh�
��f+��zS���=���Ѽ�q�D��T.5��i����ce*���\�H���P�;6�G9�56���ZuĤ�k�4]E�����,��O�|7���xk1��R1�W��E��p�.��OU�>�Sd�
�98��r�\Ei3�4ڱx�p��dzI_�� ������ȢÈ�3Ё�+}���P�Q�
����C��-<S��VW����vu��&��-����jP��g���ک�.\w��d��4��8"�`E��o0��\�I��g�BR0�Μ��21pI��b9U~���{��^�L�	aC;@e�)iM;]���2�EUzV��뱁�@fڱʉ4O�y�R��n0@��n�Fw���d�9��h�E�l�sR�~t�ŢGx*�T���&m��]h\v+#�����*eǅ���h�>��q��"[`�c���Sf�1�<�T��VbS_�v��E/V��Z�4Dh��z�����R�"V�<[Bɺ��OQ�v�m�ӿ}�=��f��ya��)B���74�q�b��R��J��z�L��0x�dL�,Hd�1�i�L����si�rk���l���y�*��ؔj�[c����^�˦�v���������j1 �@^��o�5ҁ9\��P��<����ˠX���yU3ok� �����R�֜��P�"�Ζ�-�(�0*�9�� V�}� %U$�B5bp<,��E�𧸈�d�.�*��ʁjC���w���!���|aC����O/�`lA5ч#�k��o��p"@K�S����AK'{|N&h�T��!+�3�Ӂ��H�OP5�d!:��UM���!q\���4"�lE���M���'��U�F����SN��N� ��}��*[L4zXx�/
b۷yV k�M}����o�_���D��9&����^�,�-XS��l����R�E�<2��%�y�Q�%���OC�x��ɬ��O�<�C�z^J�/�I��[[�^�@(i0�ϩ�QP*Ud`}Gq[`�B��t����$�]���H���(�(Hg�O�x��5p���К�����-�ޞ#��<��'A�q
I��ZP��扸lbSX�x ɾV��\��S"?0��$��DGC�Ek&�8TRs�
Y�OH}#��#V��פl(@��X�ɳ��b��/���=7G(&V�V1���s�C4!�,�{��e_<�u��K_ǎpkx�о��[!���]^�ze8<�VS��4_��7H�X�ӫ���?��N����{C��2������kT�����[�r���[:��Թ�K��x�w�ѹ��ȳ�I���1oF�!�G��>5<�npyS��ӝ�n��gK�.���`�&���ގ4�?(�@�BG:-��1ۑ��B�2�O�-^���p.����@i�u���x}P-D�<��-#G�)Q�mJ�ˑ�� �|^T͑͢u���� A�c�8��km�_���RL�Ѧ���qy�4V��J��O>��f-v4�5eC�i�J�y�ǚ�E�`���5!��E�"�vT�گ#Qܼ�7}���U9+N��d��A�Ƃ����I��|��[ፃ�t������6�Jd ֦��k����{�>1	zP��=с�Idn~�3Q(5?]b�O�B{�@y(� E��kO�.S��*p�#m�{i�a>q^�aI��M]̑K���mT�0�b��2����NՕy��#��w�#\�H72>N�L"�����ɇI��v���P�zK��A2�ޞ��2���<?���[_�a����β�T��g 7ƹ�NOh,Ɯ�Z�8I�߱�������5̆M��.�Xi;��� �k����r3K���n�����%-k����v��u����Ys�u�����
�E;��ҳ� �e����n�M%oѱp��^x}��z����K+ɵ��+[:��nt��	�5r��7��Zp@8���j���%,֟O<&�T��w�fJ�O �����V��6��T�@M�3���,�Ay�-�
'~]��$����]I_ץ����q�.����'-��,e~�Zo�5�6{��D�YU���[7_u�����xa"�s܊��9��(C�u^z*�n�,�.��)n6W���
�|-�fu�Y�`�E��3�LJ�u�3]��bf�\� �p�:l_\�nr ��--�>vvs23l_z���S�1�Wh�ŚSpM��@��+����W�ǒ8^S{K<h*@��NI�P�;Y�6La3�DsR�>��+zz��+���I�R�"ϰB�4ű�)۾�����L� �RE��;7�3m P̾/ Ս�Ң�'*�e~=l_G�M�L�P�|]��Fѻ�cgt�x�,5��~�����f���/�9�Lg�V�Dr�B�B�~�*:.��}���,S����y7n'�+����q>����2�bi� ���L��A;^����97�"���%��e�&��*{B��-;��t����6U�G������n�>ɐ줎V$" N~���g��G��bS��٘O��&�2�n�[5��}�J+J34�QN����(C�d�y�z�`��W9�Wcs���>��0ɾߑ����%����H-rX�G�g�