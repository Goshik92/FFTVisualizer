��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn�(���)T
O(l<�9g�)�\��ԋ�B�B�=e���X�[Rg7{��6(��@=6ggi��mi�4�Y�t)�%�2��DA��K�j�gu���I+X� � }��Dg�N��}ܻ�����~<�։���`�k|�*�	�;�b%K��,��O���M�R)W�x+��J��찄[��y����L�<�Fo[\'�Z{f�X�*�"�h��(�i���p1D�P�.��\e`�};:g[��G�T2�����䶺џ�׊��T|�6!�t���2�n^"�ŵ�I\�9H����G��!��I��z�ƀ�qA��l�3��mM��[�=����`D �J+h,�8��T�Vl�M�G������'Wy�+�3{������9��✝�ӯ!�A�6^;���w���Ja ��g��4������"*)<�e� � �S�ti��|���;i���x�Mp��ILL��}���n����cـ ԅt>s�S�7I�t[�ܹιx��
^U~��|�p1����s��
U�Hy��� y�:sT`d9?�]�#�k�x(��K[�b!�-f]Y����D������tۋ+not���i#�Pr�����O�i�+ό��5��	ɪa`�T�n��R@zp�nm��SO4��١7���(�]ƛV:��zX��ڨ��Uz�����/��'�|?���� ��.-l��,�Q3ޓ�
1�n�\����9�6�AK����%�U�L�p�-�c�A�������Ƭ����V�tm����ZWۧ��H����"���P����|�CH��^R�2⎣�.��*�vvqc��ŏݱ��p��5 "�!yү�����H@��> xKau��&="\;��Y�D,y�,��,���a����C��f|� P��B1��r-Q3��Lel��C�H�E�j�w�:?ݢ9��Y��	��#�"B��u�X�v�*|o���I!G1�T�5*a�b_ ;?[B���Ȏ���V��?J�8S=r�_��	�s��W_������R�/�'����g�1o��Z�_^��N\|�B8�s��`Тvy]HL���{l���c�|��Y�&�t螦B�!}S����<��3�w��~�a&@��[<&w��Z����cx�mӘڬZ�HQ�퇨��K\y�bQyba���q�h��>��X�/���H�I��0�NX,�,��%�K�k
�a�sVM��O�����Dބ�C�=��59TGF�;Tg!�5�o	���3��5NjFN�;��4���5���ԩ�����1�2߽�w�)��͛��4DA�ɧ���R=K~�|�� ��e�@PѤ͵(9v:���ێ_7u�?�v����Ȃ�����\i��ﲧ��-Ø�NWj���v"�o�+�)b��]�4�&4����`�u�>���x3_��Ǐ�7���)�	Bm6�N���u�f�����W��i�@�ʢ��(dн]w˺3��	ѐ�[}�L4���^���H��*a�I!X�=���0x�H,�h/�3'��*���փ�F9���:���|��r���#�qU�k�ʉ{,5{C��9���4#1Տ��C|�+~�ف��b�H�$�X7p�I�k���G�`Mx���.�<#[O b1�� �����(���|]��`/�Ա�2��!�^r�EOw雂��醙r��3������y��t���2IBH	5X�Ll��~��7[���B�_G��SAT/p�O�7Mԝi����S��MJ���
Q�[rL�Y�A`4�B���)�m9������k����=ɵCJF�Pk�䟻����IJ&Hӿ�<̍7|�!�Mm[�}��eQ�x��I�i:2��Kqݹ���EK!�'�D�x}���ل�����cn�I|]-.���%��ÃMCχ#�:i�M^�2W��K�S�%���':�e^����]j���B�� �&Srnpf|��h!���E�����&AF'Jo4�b�O���*��Z!�(W?��و�
hF��L� 7�C`�ΔG"���$�O�0dtxh��1±>��Mŭ��'u�mۭ�=iM⸁�6�xR1�p |��#K�ک�M>k;k����;��Zf�
&h���ƅ���F������!ɧu�i�� �w���n�~ w�Կq� 5�Z�sI>v��,~>5���n�D�X�;��6㢾D����݄��=<�N�W\ �b�I��:N�
S	�Ϙ��m�G
����K���m�Kz���gɔ �J���f!�X�V=j����v��B#�ao�,U��;��cB�����`Aլ�[�k��T��eh�W \[�$�y/4�-�KB���[<�{/�M��G�~�_G��zʡ$�+a�I���� 6u,�H������j�Q��F0HčW^�����Y\�F�3�X��y�l[�NTO�:�\_���c �`롑����/��}|Dd~8"L6�<OR�閘�\�<q�������-9Jo�7k�)I���|k4WR���>�o7|��,C%~;�TǏ0������Z!w�S�6Ȏ���Y�^�H
�9�=�\������A�$*�h��b{"Tnt*ocW!ӗ�K�m��C�K5�u)v'�[�j0��P�S5������fA�G�oF�{Z��諾w73��aUD;�cpZ����kV��W,�X<� ;�vM��c'5�as�S4��bvz�0#�u�å�Yi��cɯ�-$
O>Y��Vy3嚉�8K�/���8�yѱ\�̀%�$йq���0�}��#�u3��X���c}e�ṗ��EHvoKc%��X�8�J�v��6�3%�r��	�F�����=~윜L/FO�7�ѭ��@�����;�-#�<�7�W����s���.BA�A})
A���=�T���o��f�H��D2ʙ��G`�֡c��\,3
�NA��_z���Ex��Ix�s �D�œ��:�z[9$�$��s4�Sztzw>��}���]Kɻ�ǸG�9��M]Y���"�z�Uċ�Q�SF@W��{�*b���xa�el&`>!��m�њ���������~/��G�o�Cڅ���eXe%�(Q�-��;�O�&!U_7n�B�#�Z�3���睠�M�,�'����rđI��*�1.�4���I���!E�En���E��9(U��B
�H���������[�ROwج�qP!:

�Ha�Q�g��.
]{|f�}� |_��^�
2�^,t-2O��#),�5�^�xt"kX��Z�$���8BE�t���[)ܨ��Z�!i�38��;��u�_�t�m~���&��&WU�*�#�K�<�t�:�O��Z�6������u�W�A�:�!d1)t���a��į:�o����O�NN}����o��X�|��m���g��˥�^xN*���IZ���x�[��pZ�`���@NRA�)Lv8C�`.D�ꌡI��	ӵ��G@�� 6E��D$�^l4�3_T��.Ò�:�H��kOL�U�l��<c���SzlJE�\�s �z-��k��|D9�����{�f��l�ɺ핗$纨Co����%9应�녕��ϴ���g�~��Z���M^�F��`��ž���PG�fV���;�`����<��,�[Ѷ�nuSM����u�I�rv����n���"�dU���>��h���]�L�����	ZE��A�o�)Y���/�LxID�R���S��Dl	D�{	|/����s߫U�赵��T{�0� |�`"�Jn"m�RLvL����w1�4�T]�m���pd# 1B8�m�e�].�sAWl@c49Q�*�Q��'����}r�&�6A�'�����F��	�BY �Z#���F� �X�G	�	����i���b��N��U�gMZ����NJXT���Y��ƵS|ʽ�(�{~#�Z�H��߮���!�d�*�V7;W���_��\L*g茬v��z����X!�N�ԑh�j�p*�`�r5_�rw��2<vsD��:Z9Pm��(Z]�ˮD�^3�oњ�y�1�������
t
k���[R�y�R���ܸ7�GH`�ě8�L��?�]�-&�4�'�X���}�_*{
c壍Ic)��`U���J��g�%�,-�R ^~���&�n��r����Zn�K0��-����H�f}�,eJ�ن�����J�_s������m+[ �?��B�)e����,�����BE���h�u/��0��I��`�ve[�yՕ�ᐮ�hPq�{y��b����N5�5�1[=�(@iU@�65�t%
�: >�`�gz�"_�@1N�\���@�c}�gC���i���	F6����F*W6]i��V<oyڄ&� X�<˂\�m��>�c�)�K� �����}xh����.^L��A�踻�L!26a���+����z�.Q�D��.P�v�2�K'G 骍�=I%Q����)ۓ���P?dZd�#Zt�ެ�JM�f�gJ�?��A�
��
��4�&� ]��z�L���!f�%��̈����x$.�]�X�"�V�q�����LT�z�둉�~괷�P疆���IP�E�����G�����&"w���؈A)"������XN�0n��I�>�<W�=��1H��#Ì��_7���ᲀ �OȊ1�*@ 혥����X�Q��6g]W3�,)���
߯Ll�}N�6bM�ņ����u�h�ө[�q"'�qZM��˭A�Z����Z׏lM���DG��4���m�$/��c*��F��х���v�1h�%S�����*̆��#�0s�mz\VԶ�l�78V@��B�/CI+�B�i�АX�j�z�2;��T�s>���&�y��i���P��']��g�Z�1�@?�	P��V�Y��/*3n��*� 
�h8Bs)����	���e%3_�?\g�m[�=��Ϗmky��1뻅���`L�$!_w��ܚ!{V2Ũi�P/j����(Ȣ�@A2vB�k>�����E��Kl���m��Q���ƛ=�^�J�鷀�.��7����5#���fԌ.V���Z-���O�,�E��t�K!��*�0ޟ��o���fY�U��|}��-��( �K�b$��ޓ��YR=-����tװ\���L��a.���7��j��^���m�_Bb���&uW�3��#�>s�O��T}?�~�x���B�q��9�إ��x����K_/�T3P��k�"l�d��m�1d�ZA�->����;�E���N��͒��_�@��s�^�:�lk��b��V��!H&�#�p��~�@M���\�=��.n��՚0Q�M�h��(�:���bʂp��G��� �����N3E��v��vקg����?�y%Rܝ�x��.�P�t�L��|�p�����4��ٞY����ss�t�����C��}�TJ�lȺH^��Zw�#���w�%-yt��D�ˍ(}��B} ��7�'`�ƣ��K�>�%����pLkW�qf]#��������X��� ���;��[h?�9�� p�?S]�b�rGڒ0\�U��o�XD4���s���r��}��B�%����Sj�٣�2\$4ĭ[n:�Hhu�̵���T���[͆��
v�c˪��	��X��m4���&����7i�s��� B�K.���6�
!����"�}B��.�`���I��Jn���(�Ed����D�$+l�O9j'r��XpC���G�ay�(����F�ExP���9�i4m�'l�p:.U�ڔYjHq�R���W��C����,�����r^"㛍 �� !S"��K��v����H�×*F�n�õ�4ß�+G)d��|����(��r�e�(Zh3!#G�h!�`�1�]�"�ܼ������1	l�(8k�
���c�X1��?xށD `:���T�h���(��'C�y�+7�n��|��ӝ�x#�3��m��Hǡ�2����f9�#�D��+��V�t3��n��7<��[e��$�RCgQ�U&Yir$��%�=d�x�:H�_���)��sWO7tt7:� ��ʌ�q���2=� �l&��5�'ǘ�z�\����Xn4sA�V������IYן�>�v�. m���ÏV�iLA�V�4�v��E�g�k����)�B�dc�x�C�h��S�(��-*+�*����T�>�:
;��{�^-���8�a�塢��ʥԪᦿ�t���~ꕿ�r�����J��.�kZ!l�/�w��XPW+�f���%EQ��&��y(���,XJ�}�z�f0�V��uЗ_�E}��7�6��/7��u��_fqq
�������������TnU�A�="kh�+��������&�1��}�����	���Z���)�㕸���좊�&��+\A&��;���F�^���3x�s�L����j�˕(8�zcO���vɂ�|�Ǹ;dyc:�WۑUA�r�ހ#���[b{X`���}Z+�,2�+��&?ka�r���fQ]#\��������;�oG4�� ����F"����'#��I2��]}eR��-�"��%�Pv�y���N��MV��C����%X�l�#٫���q��D�4���&[pnJn�p�A�ái�d�zyg�~��6yϲ	8�j��6)��~	����#;�R�SX�S���U�P5݌�Bą�yZOϓA�7�F��D�J��ժ�n(\�T��E���rQ����\��w��	+�*��"^�I}���~v���0=�@��?U��z������wlH��<�霨�����=��`��6{��M�Rfj�J��B>&���#3�4�ͪiE/(1hA�VI�}ۺ�tcA���gF�LO�%�ؗ�L���@��1y�~tT�/9^�����V�9M��z"�F_�?w�V-@�X%��;�)a��>�:$G=�;�PN����]f�vi�>�T��E'X��O�;v��҄A�8`���f�ݢ���;���a'y-1�o�rʞ��jE!v]H��Y-<Ų�#b%�4��%�����{o��Jp߯�_�>$�d��}O�����������(���f��	�;Zc0Ó��^�W2��7��Hb�|=�*p�`���х�`�G�&0�x�F��B���%yo�8��i���:A��bՌ#��Fv+o�������ړ��g�Jfu�� �|�W�Mk��wUK�]Ճ��l.ëL��->9̱غ�|d	A�oF�tUY���6v�����{mF~&��^� ����a���~��� +��u�
mY��0�V�R�E�D|?�����Z���oy��S���U�}�2H�@ﷴҬ ��wM�d�M�@�S�><a�5 �&��MLd��N�!{�����ɔ&��p"+�ה��\.�B��j��Q��Y���$�C�Q����Cb��"���cN�H���+=뗸_���AFz*:�K��fѱ|���������I��E� j����b�:�B���v%�S�������^N�C���!�;Wy�q�x���j&f(�2�g&Jr�\��8���?�e����O �/�2�(��ea��U`��������)d: /G�1\d�c�ٖ����15�Ȳ�÷��0Rh��sE�`�9YD�.�K��B�):���G~��O��尬"iRf̋�
3�N<ag�'b"�--�����M���܉Bv�BC^��e�3CO	�H���_��@P�Wʽ\9T�����ú���B������N���S��Ƿq5>A���d���M��r@]�*��6�PsQӡ@�fE܂~LyV�œy��]�����=��e0T��X�����\6�mDs��F)H�B��o����Q(��M�G!�ִ?�C�qze&��f��{�{�S�֥�>�J���s/Z����ڔ�n��\FI���F7	l��u�.�Y��|��)�����+>���g<����δ��ѪA�z�؁?�հ��悀���{^I��ayq��3ϛG,<a��\�����_ާ�<w�4���"�i/��z6ո�4�̔��4.~�gՂϵ�|=��}g�HztzD��7a�O�˹"%w�_��M-%/��a�� �A�p!3`�3��d'k��n�Q��{�E��"�J.�]��<����9���NY��������M��;�+0EB>�S�I�������+'�8��ylpu�3B�[��b���y�B�9�B�o����u�v�f*�)*:��0��5�w��'A+%���	�U�[.�3g�늀~
���疮��K�v��}b/�悤���[���i�˥�p�O�u͘�Eu��������v���2Rz����d:[�T)qE>�[?����&�똾
�W��Iz�M
D0A'%cT���(g"���6��[0#��� �7{�,�r$���7`A:��';�Q�F�R�$���[P�����و���{�����v�J���K
g��WW�:�EL�ߔɢ��b�wb	�v#R���[�MK_+����D˭��G�=�m*�7dy,ɋi�kmiZZ�Ɣ,�?���8�;@�����"@*W�މ�Z\���9���KO�Xˉ��F�6��܌�$<N��Ke�ؘ��ƪ�(RT��b�{�t����I��AWј���s�5���P�⽜����c_����p�4��"�Dy:�e��y�/�{&	.mq�p��z�����ռ�� ��Ȟ��E�V���U�5�*N�"%}�mZY��6���^$��D�p?o08�>��NbӯBo���D�Q�\턷�H�#�8�߬9����b� [IN�-����>����邮��T���s����K����������9���X@r�(�o�'����K����(�'�ᨅ`����� o'�{��r�S� a!��V�b�̨�ټ�0��A#��v�@0����}yv�1�6�4�a�ޓ�×2��7�<�3c���O��b�:�_G@S������M��(-��Ř%�ۧ�����\����t�y�Vl�<�Yht�ӳ�P @���4Һ^R���]�zn�G�t�	�Z�����b�W�����>NYǑ#]J��n���Sw7@k��^��)Ä���.���i�lҭJ�
:�����`Xw	nI��,���Mja���|Ӕ�fM��G�k�Mr��y�qC���u�a�Ѝ��-�5��.�E �Q��iz�'�%��-ݥ��{�b0��{3SA|�Lc	�6��h�[�C�2Ľ�2`�j'(����hT�$�5�>'xۓ�n���,xDO�g`Bbp\ݮޮ��?��i������y�Q[u�]��!GZ��7q�m�P7��i<p>�䮜IB�GUbĠK���"Q��c�������Lx�E1��/�{��q����4��nW�R��?�f��Wu��r����FPZ���gI=�C��|�n���6�Dl  �o�&��\i�����i����ؠf�V��ǆL�1	�ٓ�U˵�|�]
���6�;W�λ��d�ަ﵀_�g�{��r�δ�A<OC�ꟲ%F���{�8�J�̽_i�Z�66�R���=�\<��Re��W���5�d�;��us� �%PW�l����C�f��H}L��B*]�C>�/A��C�&�M��ÙS��aY(��r��+���ާ�K&����$p?&A׬�"�{��#[od�;0$�68EX f�G�Q�heRk�=l���-_�X�)���p�B�k���� �Cs3�X�p2w�K�iT�,a�p�Ϣ�K���Gm
E�|�NQ ��/�'��W��$ۜ |#�������rL���~}��Z�ĸ �:�r�t�����\p�,]l���(S��a��Q�� u�6CYD�-V��a:/b�p���=�g�t�{�E�9��3w����
z�OJ꜎(����45��喪���q$�����{��AFO4x A˂�{�]A�y�{~[Hk��SS��7��s��o��k�KD�(� V�V�&%+HW�P�h����Gy��rqC��F��ܢ[���T+�>��;�ǵ찰��l�Ռ�F��vʂ���9I��*U뛳���Q�c<�CfD�a ���  �zM��4��u ��d�MOmBX����R:m鋭H�0`aΣ-�4H�?���܂���t����$�
34}b[J.�sO.�ue���2|K޻�;�̄1�����n�O|U�
�j���	�O|!nUX#�7���$�uzy�u�q��L �;�c6�p�<��#CMT��[T��5F�A���*xV�y��ZR���������k1f�1���)�˪����|6������Al����)N��Jb�c�J!V�7�[�sz�����mz���t���"r�z��9�'�b^{Nt�a���l�7(�� ��Q�z��΢B&���^��r��q�bc��<�A^�/�<�,�,|z�+���F�
�+�K����Z�ڞ�`�?��d[�r̿��s�p7�cOx�9XQ�O����i�-��	q�K�@�8w�����7՛2����D��\UǤ�PPe��$Ar���0C`W����/:�;��-j<-�?9ay��9b]m5��]������ƫ�u; 4� �%�<�?u�:.Lº}��d��s6����b�8��56�ػ=���󻕪��M��؀��c�S��]#��1-�;�duȍ���K��7��� 폙�)fL,p-%r��Ċa=�0�}�������7�M�s�����c"E�\Gd1<R��Gr��8�f�g�t�G�X�z����w��T�� ��Go�)v��O�d�[�jA�����ɜ+I�Z�&\��N@}/h�\7�]�J����+����I�q�"��[�$`.���U�qr���K�Ǳ'��Rbi`�im�^xۑ� �,E"�"�:$<i�À�<��v�%����d�\�ⲑ��&���o8e�g�'T�z��NR���i�������=,��$|���bផV�ހ�{eC�&!�@���0� W=`�� �;��H5c��`�31^��*�U:��B�����,�\ ��~$��ӏ����KdB���j�V��2Na�����w`�������ꏔ��.���� �T�Ċ���t�[���:��m
��
Q�,�pb��%���(���aT����l��'9�%d�>2 �	�����`��3��mt?<Q��K̾d�z�� E��9P���Q;O�h��w� ak���H!�p�fG�:�-�ݱp�XR���_t�<�PI���t����/Hd�G?��+�6�N�>�M��xv��5+���MP�������J�G�0���>�Bʻ��`0��^�w���iEF7t ¢�e4�Vl�b9���C�f(�١�f��BP��
Yb$un���7-Zs��k���J����ԟ�'�(]!4�~���ے"Nz��(�Mve�8���2&ȃ���4ʷ�J���a�5C�����>d�Hێ��B��uo��q�؞ElX1�;	+���q_eo����O���U|�>�l����I�+ ��ց���k�ϗ���`�o�\�Yq�$ŀ���=0��RnX
#��
F��Xg]+˔?�,���j@BT���Y�^�	�H�ة"��.V�3�L�g��h?)��z�4��֖�M�I��;��"��@giq%2��F�a)�y@K��[#,��z&�i�G����Q^�a�����²\�r��02Dʃi���
��^��8u���Fj� Y3}T4�*;�9��tv��l�	�|ǆ2>Z����U�E�U����i���
m{��̀��Y �d�l"[����09�$����x3�'�2>�Dqo�O~�6�j�C�����RA8�>���x��/�e\Za��6d��E�*޿���>�N�0$��B\�K���'��Q�Oo�������x��I�`�U�N!lI����R�zx�����a<H�T"$1ѦG�\�8��`�>v;"c��uc��ZI�j�g3�7Xx2�D��Ċp�s$z�(��x�v����=��^��)�{�ꆐXL�<���yTa�I\{I8Nw���I�<[0K|c*i���[�o!������9-⳰�3H$o�w��ΚZ�����5z�\3��`V9�~�\�U�G(���1^ߺ&�M�}K�^�<��g'G��m�v�·�݀6`���t7J{�Hc�Eod�+C�Y��DA��-E?�QpHִ]�(	��'�l3��1$w�ؽ�c�S�h�@���e�ٗfȎ����P�Ԡ	���S�����(z�M� ȁ���y�d7����ɘ,�X�<jG�4�@e<�h��'ӌ����^�*02�mR^#T�����k;��c����`�Q�A���ok��1������.ߍ&�=�M����xt�l����3V�%@����rp5�Ă��p=�a2�����}�0�g�B��0���cQ ����W��?ڵ��'���� g�4/�X�:�<�x4�%W�Y���
s#u����X�Wю�#���*G#���_"u�+]�BLc����kF� � h�	B"��X~��r-1��zU����1N��yO��M�u�⁁r$����%�	з�\3/`@�G�o��}kN�맖���MH��샌7{���'%�
2�?w�Z�~I���0'!��}QoY��t�}-sj����r���Hĩ%Ȅ�{��
Y'� �mm�"V� ���s�Xz6K�j�����~_���V��(.u���4i����q�; EU1�IbT����D�ST��_V���R��`��w"4�`����DH未D�O:1 U��_����R	�^����zLd}^0�*?F/͗2[��Bz
�5�6��ǕNFi�h&_��BG��(�vz�0��t��x�������m��ٲ���E��wZ����&CT����O������1'φ/��.]���kNH��m-�h��R��s��E�����:C,ACm��7M��Z*�0i"��2�{��� ��ŗ�8+��6Rݏ`I��z.�C��݊R(��XV��n_n@��r~��E�	�*�O&����F���(3���Q��;��Sk6m���9ۍ�s�j���^���K�k(D2��I��]�d$')��y�U�����B�Kz�q�����|��u�U	.ԑ]�Z��-��4��G��~�˄h?�\m�0bk)֙l�beA��d�wEw��@���g��p1b^q`�eX�8n���w����YK�"C�E�d��Z^���Y� �:O%�oI^��@����G�B�
ﰀ��(]%HA{��9%��U��������'��GX���Q?�%�Ĩ��1�k<bl�֛!�ּ�ҥ�q��;���͆�D�=�*1��:	�رfx���i�?��D���~����ΆY͙���*���ᘠ���i�ǔɱ��H�^K�;���q�xl��"8�G�}M���d����/ݚ�c��`m�Y�n�^��Г�B���]/�c�y�͐h'C�N'd��d�׶��@�Z�\�D�$�
J��[�d�e¤�5"��i�7L_�( <�Mٷ�NT����h>�5��oz�9���Z��聪
��<�~$]��p<|;v����q�$��%d�����i�5���؎1�$&�̽-@/{#3$/�.a�P�j�3jP�Z63�p��󄍹�@�Rh|6F|���C�B�@�p��
�g��,��^"},q�F�	�Ag#�!#���IO>�jA�T��Q�h�
w�8���������\f��^�7�%�'�����$�6a���f���ʨ,t�˒IM�gb��1�� �垾]������m�Q��(x{'���12Y_�^\��Z�ii�.�	��?�_�S�P\Ǽ�Yy��ѷV�H�g;�m,�#��6���2j2'��}�5d4���.R[��sz7!Pc#�>�|.�%��� 5���+�m��)�x�#�	t$�c���{�l��!�	�sS����`�Jah',�AI}Ū04?W���&˚>&�YQ�(��#�1���8�D�Ke��m��Lb4׏�$�4�!�.�-ey��T�ޒz��X�����ƥ�=���P��jܾ&��U_��x�O3E��j�h�n�T��(�a�d�s��|�{i,%�8�W�6�T|��4wҧ���m�9���7B��])����j�XK�C�t,�Xa�CQ��98��2��ҝ+-u��wz���>L�<����c��w�>ƾOP�DXg� r�p,���`�~5���6����W�j���i��������ծ�T�vN2���|ce�&�|x��&R2`��ީ��5`z�f�ߝ�(���;�p@'�*�n3��I��B���	M�D��m���Xd��ՙt�x8�$�/&��u�д+���$��ţ�J5V�{U���F]�n��l!��"ˎ���+�{y��W��Q��5u|�}]&.���4_�Op"M4-�b��/3�ŝ��ɪ��KXx�WH	��L�N`#
"m���ف\�M֥f�P�v�m�axDǄ��#�:�nVZN;_"�	xB�u���e�%��/��\�A��z/�2C�.�舍��Uc?薡� ���ش/G3lha�,���9	�|jBG����͝�)�>��z��a��O������'�SA�̖�R�p���'%B�u\2�$�ד��N�g��w��/���yx9�>�T�i����kI�iN�q�u��y��$S�C�E#��%W!�#��R��e4�>�.�T���:�2�j��ӘR_?96��-�烑�
eN�`�8�6��\y
�7�F	wo�T
Q߇7؟ت�H��s�@�نH0�H��S�!J��c��Q<�:��Q_]s���9�N�	�+r�ZI��G�f��I�1�"�L�� )3gO,\�\,���g�f�2hB����EB`b�h�CLMVe��5c^�yĆ�;j��~$٣$�1|���sI����2��h1�����X��Az̓��r�-3�#�D�Q'�q(���R?]�mq���Q�B�T�;��rs ��S�
�m]~>���Tb��m3A�y/g����ha�θ5j����:�t�Q�-��DZ�+������e�<(�{v�ț�|]���Ӷ������S�Ṣ�g~�ݡ) ���Q�@=
C�b�<��x��:mǛ�r�6t=@Wx?,k�<�*l|
;��S��|jHUő�w�),ۜe����s�`���m ڃ �47�7�?�P�:���]q�b9�U�Y������O?Ҟ�u�թ�*���^����˸!����=r�k��@|�p���a�FM~�ӗ��K��86���ͳ�m2�����i�Ws��!A�Z��0v�����=*A�4��D�I��b�iy��E��B��m��@���x��&��z��뤶l� �+�
��ڨ毟KP�[$�I��ۯ'�C4]07� �"��D��kn7��:/���='��5S^`���e>�olZ=w#gU�����dl��p�j���V:芅(���u��Hj�٨�q��=���ev��7���!.�D���i-By\�j��l�KR3�q��|}]��ibUc��VL�8��'��!�jz�K��K�D>]��c��uAE��P�}�^������u���Z-���Px���QÄő!9�Np�.ƥ�j^�;���w[`�-�MS k;��S"a�A����х�ey�
�f�[�Q�g�3��_O��������u,}����r��QK�z���������K"�I�X|-��=3|���gň�ܵ����e<�+-�]<����e���Պ�"�<��;D�R!��7��g�E��Sg�4�儂:����e<�����NO4�-θDf���H�N����S��%a�33oj�d�!"�-E�*�_j�a�x���/H�d7?|0y�;/NH�*� �&�ء��0�lB�zQv��@����ޭ_����EҶܮ�gt=�S3y��r�!+(=aT�?�0��C[�w.���wQX`�xxUPmH��e|��/Ho�A&Q'JZ�����ñ�5i�����m#�D3-Ԣ����E�=�L"x�l�C�S�fJ�n��$������H[{Z�pc���L��w�\��=)�_Z�2��=��2_%����1�j9V	�l�v��u��%�y��)��c���S�c�tk�����˚;a%�͌�f�'�y���M#��Ԍ�$�E���3-�%xf8�b��.��p�х��s�AsGE#�������l�-�A�Hk����o��H0Bu0�?�,�����c��U�Jc�Y౸�`+п��?C�D�;b�H������U���?v��L�v[[��M,�9�L��yu��҃�� �L8Df�[�u�s��m�4�@E�`�W�2��ӧ����I��g�<�./�׾i�E��؍`I�F���;H<)��؊U0��ݿ�Ǌ�Z�~���Vߊ���IB�o�)-�k"7��R�#��F�D�;kY��c~B�N��o�0���*ИQ�[*}P���1W�&C�%� ��hÝ�V�i+b���-L��n�.DBb���t(��F��y��F��q����E�P�K4x����o{����>ˋ��E�aR�SO�hX�}Q+ j�ާ�uF8��g������U���^�g_�ѽ�c��H&#�$�6��)+0�!����~B?�*rdN��	�����*�xd�U���	��`��"��D
�~���6,F`�Ҫƅ�Ag�N���h&я�t���� �����m�S�q����`�]�y�!8�f�s�$);�{q"�ӖY�?L�8��x����H��Y��o��@��/C�w���eE����e��O%����p��~?�L�^_�P�g�n`+n��,�#�	�3���6��K_���C��#~��P;i%SN��f��*�:��O�m8:x@��3��-����z�eH���9) B��6���3҃"a����d_���}G����LK���|i�&�Yqj��+�]�������w-��%TӦ���qW���HW~(�z���뾡�J��HE�P3�4u�Y�C��V���I��j�v)���NCV�$��$�(�$����9��Ⱦ��Vc���F�b�?0����ɫ.P h-��h��<��{I�m�~��t3�����g�#��z7�������[1����>��^�d�p�p�;�Y��I�7����o�J��P�5i��n��hpe=ֹU��\�Ť�O�S�p7�֛�:���՚u��dq��BuϪ�8AJS�!�������;�0n!����������0k��#�X�M�Gx�3|�j.q}{h�FJi��
���&g�c��6
�+"n��^ ����>���ል�QG��maټ���ByP�r$�7�wk��[v�R���Ƹt^^�q��fss��lF�`���H%�[���������Ʊ�R�Q3��~e��2�l�|���d5�]{��[�>�L]�;j�z[�7Y���ep^cí�Do8r����ys	�5�Bjq�u��ҽtN�:ٌ�}��o��Z��%B�qa?���V��9k��%��S�(%/)��Q^fT����n6
q*���m��ү7�⪶U���J�:qȒ�����[P���ynr�PB���unn*-j���eZ���C@�'��(��ڹ��i�
���%ݎ�(/��hP1�S�ä��B����s�m�?�v��M�kT��>�f�o!�,Et��>���}Ҟ@�-�(O��i�ΒE�za�6vU.��X�GJ����%ͥ1�,-&$��	��,/���G;F�%��Z������<5j=��._�B� I�1�����hnw�L>�1u!s��n��t��)�<ÄX���x=`Ԏ����K��j.G@iߊv�O��o\񗕤,�m]�CYl;�Pr������[���e!����������%�H�g�}-���B"GPA&P���K���}��r||�$�b�����y��/;�ӭ�G�c���kP;��x{�1�X�����~���J<�����������f8ZD�9�G��&������҃i'��chj�d�/R�^ׇ���_���u+��O���2󣼙q�"U�K	�aU{�����O�g���R��{��K��Bġ�tU����,&�����pc������
��ď��8�טb��y���lg��` �v>�g� �$�a�K�lS��3�I�j�MN"�����w��.�/`�u��e��-�젗m��C~���!9�[r:���F#^�������i4	3Ɯ�)��?��3m�W>�s����8"�9����<����
��\�c,Ohؼ�F��.���wz�/_7�FV�W���:�9l�V�å�R)K*���^�-4�����0@as�2F_e��f_��˴N�r���?�oY!ݫ��L ,Б�^��ov)�S9:�<*����ѢS�өvh�w�8,�4I�A?�2{:9St*��[mp� �!Q����<��I��]c�LӢ,��#����~��f����{n�`��>������&�d���7W�p�h����YooH�o�7��4�]�Xy�P��q�쳲���NJK:���I��� �x�ڞ9D[M��R�(~.�֘O��Oo�%����]����Gk�c�3�U�zb�tu����	)|��ҕd�;�����#�p���p�;��ޱ2/+ƒ�Nmd��}�TDjx�֍ _�MW*�sl95_��efՐ�������R5�w-���)��~O*�-2�V��ת���Q'	z�5 "e��Y�.Z� R41�,�D��� �iѪ�))�(���k��	�PЩ��L;�o��}�y<��9/����	�̢��{��
ϭ��I���?(�=Y�B=jR��*;������<�b����h�j���U˨Iֹ����i�������%"���E�����vX6�D��������Iy`-����W�٫��V����xׁ�c��X�@@����g5yۻ�kb%�����%G.����I����M��=�œ������D�;���(��M��Y~��:(�����\M���Bw��  8���'��ɥ��_<��}���o��c��S�+���Bߣa~׾)��&�rO�=$}� Y.�#ኍ����1K��qg����sn]�.#�N�ө�"9�iwC����%0���P��`��C|�m<W]��Z�r���D�  Y����h��I���L���$��]7Z�N��029�E$���3J���M�,ڪ~#�7�����y�L���r��G-�;��/��B�7�?��b1��>"�6>/���-rzqQ��H�,�Y��r�e�q;���` r($�άM`�.�vޑ@+�p��&�;��$~�l�L˧�+��2 9� ���A��@�ĝGq�U"fo6�'
�!�ޣ�4�7�����Lp��Z}�(�}e����u��_�7�F;Iqዓ�9$~�9���w��XrG}�v	�5i�´�q�Qk D�˾
U�?]e�<��L�Uo�"����z�	��@윮��C-"��J}� V�ť�<�6�d0m�A�O3�e$���fΔ�լ�Ae|(�pw��E�|ר��9~�ު������dq7�V�S���/�w�{`��:��kt��	`P�Q=�ޑMU�f�U?m6)@d[�Տ �&��^µ�jA�W~��JV�MY�+|J��%eg��=s�%��W�_w�����f`��h�;4�������g3l����+�ܝ�Ŋ$�\J4�%�P���7�L��<Q[l�Y���l����-�gނE�ǀ��Mی�ݼ��Bp�zqA�"��e�����i��?��QXC0o2�|&E*"�M�SX�FIǿBe�1�ݹf����#�Ϡ+�h@Ħ��﬙��Eڵ)�&ֶ�IM`oxC4�t�U��1�hwy�� �ְhqmc2�&�;�\ek.�ŌN"B!�xՏ�1�h��/�`b�U�U�I0�D�G� <̔�zQ���·���4�F����`����;�*���<�!��2`��{�6�ш�vK����\6�X�� �*5q�&B���
�lG���\�Z�L�FOH$�$kV�6lȆ�d'�ϐ��"4 ��XnY��)~�|�����M#�|u��-��	��O�7��B���Y���d������A-�v!��F��6L-�/��K�}�w�^{#���; ӥ਍�uT�Mn��38���^�>������j��ؕ�'�y�Z}(��q��y��~��/,K �1[[J\|kf��´q�Q��F<P7��G݈�d!E�FA��-V��p��a�. /��F
I���P-�95·:x�_ƪ��+�-���EK�'�.���P����˒�iSթ�2�@3�����{u�F����2�1���o���Gc��r�tw7� ���^�N��i����{��<�|��wk����9����b��Y7�N5�^�X�z���������h�~0�)˶�[ _�3��4n�a�0�5��o�F�F8�{�q�M�t*�e�E>��O�`ANu�V�,��N�s2�]Yؗ���&���������g&:��.d���󳓟��%���O���'�gX�Z x��w`���9f2w��nh?�U|���Eg�@/�Q�@�<� WZ�K8�x�y"���9�(B8�?n��Aiwp��O��2H�{� �r���w¢���$���h|����(�6
���"�Mx}�e��f:�3�s�*N9��jg�ؗ(Z��7��s���g@��S<�3����.�c���(>�-�-���$�j~����LK�Hh/a�2+��������s���hU1㸌m%G��W	�&�J�m�W��Y�e��ŋ`|���v������B��0���;���_�j�$D��ߞ�qp�h���߼��a�Q���'�v��w�����9���D_����ܢgY�9�A;���'쾕 *�'��ҋ�A����s��`^��sO�+��ý�N I�d�UI@�|�ŵP��W�PP9�k�m����X��W���ʾ���I3�v5@=aW�#��	a��M����O�OM�����jҖ�"�����(9��Q!��s&�*uō��v�0�f��%�j�����ӓ����(@3;�m��
:- C�f9CD����=����若�Z � 3W�/��@�C�����7�E��Ջ�$��V�ʝ( ���00���ƌ�K5��ro�K�ࢡ���?v�94��	���aSM҄��3!��	��5�J�E���щ���+^���o��KV��T��� F,�r�v&�'�ݮ����z���ER<)N���2���>c)�mӼ�E���j���{M�1 ѥG�p�����#����n�ձF�o�v|6r�,G�le~<��&ԕ,Lӥ��թ�dO�A���_j�'W*�[��h����f,�O�w�(%�p_*���eE�~1��c�2����A�7�!�bIJ3"
�I�g[j��k�qۧZ��2��Z���<���u��G$��k2
V ��B~ʭ;�t=�2{%�/���*y�a"d�eUU>ϳPr����q�Z��E�Ր��r�g�AG|�<7U��ө�'G���vi�m���E^\�����
�~�m��j,�3-���f�c�)	�Q�-��/�cp#��L��*�a���s����[�������8jS88I�ܡxa=�0�����ƺ��m[|�'�>dQ���� {ﻢ,ǀG���{D��"6��.����]*���^�&[s4Z�m _�>_�Ftr�T���&Z��i�wAw�B��|�Xs�.����clzpr�j0g˄+�!�}*��߶�������\��h>�b�^�(`7�)(�[~d�Λ�8����zEHW���<p��p)<�W���IF������C���	�a#3�|�x�9z�m��;^�Uć�9gW�U�@�XXc�ʹi8��U̐Mh�H{&14+�6��(q�2CĎ��T��HǬ7A?��Lh��o�S�S$�O�I.�j��Ĩ����Xf�{)��C@z��k�C�� �Пq0SY�[wL����#c�,:5��&��5���+ ��@n H:��n���Jm��xw$�`c|D��o=�G�I(��$;*��s}��6�-��JMj�n�d��\"��H�4��^�MpzL�c�&�xF��rzT�c~���u�iÝ8�Ԟ��4�����.�?%�K��i7�S��F�z{ ܔ�J�C��ŬS-�S[��K�96�VT�����)Y�%rzW�̅XMZH5KE�i�r�s؜5{/!��5m9{�l�L�vcY��wY�t8�bS5����#���x���KO�.���GUSk��/k�;&}��.�y�̺�n�ۭ6��@:,������1!�:^C���=q]�e04NX�<>�R(�_O���AD�E����o�	ZE��\�V���j�TW���Z���O��8�X�mf�h{M�PS�8d��~!8z6EE�n+�bc0Өj|��V<�����V]��K�	��q�8+����b����6 C� a9���\�q�5��G��q��S]�7����B���dO�6a7�h��. �ƭw�t��P��3z��%�m)��J�cfh}WZ;�J���E�3L���7�?��F������~l	�#?="ǆ�{�-{�ŧ\<���F�":Q�a������gg�������P��+{eW��Qu�'8��A�V
��sX͞@��U�*�p;MMl�p\�r6� @����R�
9ى~�ج}�#����_�e↸BF;�0�9�]k�R��-.cy����=����X[f�6�)U�@s:���%f�w�{�*'ј�Ќ��^�W��n%�jM	G�4T�%�?���!�߸�O���-"��I���<�V������$�,3�Q�C���`���3��<�Z�Y �+,��Z��ࠡIx�YC<8Q��XgӲ�n�mz��6�0�2�n��`�:�.X�5���l�*{����#�ӄHL�AGRR��t���S	�eȑ
�^,-�~�l�x�%쁮C�X��F=�pP���%��n�Qm<��8'��1��<�R
�Wv�J��:�т�������/����w
"�>�{v���*v�a�~�,6=�B`k��b|�{�v&��	�nnU�D�PC�H�r(y3��rn<�L�U���-�F�9����<�K��J�~^�i�<���c�K꜌d,�J�7%�u��� �QW�[�t����Ǐ?�><l�p$ԓܻ�qk,�8[BF�iO�d}`�}J�a�y"���t�K�R8�]m$^G�V��"9�_��Ł�$M�7���6CS&`�"�=Uv8$J:��ϔ9(�b4�`լ?�N�r�Q�SYf{/��P�D&)j9�������F���V񢱘�����o����tQQ)��B����7KX"�k>}f�k�b�b�iv��0�`�YB~ǰ��iȆ�m��Q�1	ZX���C���\O�gs�`d-��b�-a,����E����_#������'�׃���g䞉��):���_"��٦���^�t��|��o�t�j0*R��-���E/�ҔF�V�\�#��K��8�>�O�Bj5},>M�h�"R������ �q�G~8ۀiy���21@?%g%G/������:'x��k���1�X�;����N�c/%��2�C�a<)�w�=7 }�|mʨ$�0���'�EK��Y[S��h��q�E�y�Q�*�wX$�LTP��pa���L�m�$�����n�D���.g�_>�&�lRl�^��Ϊ�t#���-�O]_1L\��xZ�	�G4 H�@�]�j(sb�s��8��MA���"J�h��m�!�TP��
�N�u�gp׫z^�I�2�j��,��5�Y�N�y�>�����F�R�T��6�@X*�o���N�S�����S6�f~)�:�z"��qE'y�OG�Q\&����sJ�:���������ɒ?�W	���P��㣭�L�h�S�H������zE�3AY��T��� M����D���҆c����R��ڡ�
��2�AW>)��
4f�i�Bm;d�EJ'�y�h��"��Ϲ�g�
��<�����v��I���Vqe��v�^�	�$4�i�O[�\�wJ����f	�&�PeYe<}Z'��_f;l3�@���3����;�Zĕ�^��-i�GyO6���.�<�{�@7-I6Ь����U�����:xI|����}�
IzJs�cBhDτ��>�3�EB��J�l(�J�2;5W���}l'8S�/����FH4e��0�؇���f���8�����_�wP�沀�`=���>�E��J���0 �Nꕙ�����u���$;�P�H�xa[}���9"Vߴ�o��-��4���{_v:�n��F��Tcy~8��Y�(C�ď<!��eX�#t�/!�҉-�����h�j��a�B|�`��A$i x�O�{vA��~�7�z
�eT��p@A�&��2;�V��3<�f|?b��3i?Y�o����N�/����� ���s<-�#���y��6u��׵.X0�s6�\��M�9p^���4@B��>���Ț�ɑf;�b֦�)ؽG��9�l�IW%��I�R��6\��_ٛ�Fk��;����-�����3"�Ɔ`)͐���jͷ=��;�0�)�E7��O�tv!׼%��7�'"�F�7��m�g|�N'z��6Ce�:t�RF�At�e��O�2J��TF��p�G���me�0#��E~��>$�1@�,^�#�I���w��`��!6�A��
����ܩ�8�V�����n$�r���Q�Ud��Qep7<p�PP�����01%�%x�17���t����ʪu��Z2:��Ƭ�T��'�>#IR��Bа����s�l��|e�FQ���Wwc�>T=����:[<U�G��Ob�^K�DG������V�[�Pލ��F%��ƛ0�^�b�{�qv���Ͼd�xz�G�J��^�]Fc�wGɂ{�³.ѭ�;uV:6�_����!!�<,Q��H2�y���O������@䲳��8t�f&��FY��+V�=ǆ�W�8D��6fp*�xE�1�DQ������O�,pO���~��b*Ѹ�g�������1	����uK�j)[x@wq�~���~��"^z��=L�D�b8ޙ���=O�U唸?��B�pJ�����m�@�K�������@�ϣ�o֖�Ο��Φ�s]�t��$�d6�;�SGk��JU���t|�[[�iג���_��:�|����`�
#h}��a�ӿ{5C��=�5α��M��0�q�9�\=��:��c"m�`6��i�H»-�β�����z<�72�4\ 5n��Z�����=QM~�S)���]���[�q��e���!l%��Y��0��<�I�	��Hw�U�y[�[ e���� ���ۀ߉�Ci��.d���Ϫ9L7y3�{a�7������m�p�\9��阰��c!���pY��l���O�_�>_�ެ�k�������`���5�����y]Q�?���A��IVP���ٯzx�o���!#�&�,2?��q�h�V*�#��d��ӫq�!GwP� �D��.<C�dQ>��kT7�1�4`!�a"��v"���u��Ԓ���r	%�b�ཪ�b_���a�!�74$t�!�٩�k�G5�=̖��-��i��#Y��VB�L�3�9�����*�nS"�ޥB/ �s�!,$]�Z�ӈ�3�n�������(_�9[5���q��x�E�AV�_(B��=���ľ�w�\+������r��y���e�L9���M?�J�G���j�ڄOW�����e�hT�p��Q���z��ٸg�d+l��bx�[p�]�9��(�
���=,!�>s�foy���[p[��$P�4��[����2��=�j�%��6I���U���%��ٲ;���yM}D���J����Q���p�
�ʽƿKB7�����B�I���ʆ���%�)���@Ր@K��᧬YU���@�g@pp\`��k�ā֋�+����ɉ�t�<.�a
���RV[�(fS�����ct��������N3������ަdu�����*�Q�r�S@�<q��hL?!�:G��f7k-.?Gհŭ�f�Q�h���?�8a% �~OH��r6�����,k�}���iMg|�� >�ZJ��9Z�#�X?A����ۓ2,ΰ̚��D/n-=�d(-�X��Yo"&C�bze�':�r͵=s|�������5�q�q����R����f��r� �[x	�R�9N�/���Gt����.G���h9��D1�L&�8D@�b{���+��H �Q���Q���j�_�ѓ�e�}���oSӄM�2����k܆h�8�y�:3�K.#�����!�K��/����J�7���s��Z�r��u�7](��3�ZӨ�NB��(�X������[�u�"�\S��2E+čqI.o$���;-�e�m�vHuFi��������1
1�!��ğ���<r*TFd����K�"��<�n/����O��[wg �g92g
���$Q����D����	�#���o�uz�}����Y���2�I������T�v��%��8-W� JzW^AbQq-�*Ʌ�;r�w�D��Q؇��nZ������F~t�=J�k#ɪ��v��޳����yM�{�˸&��je��5=�kZ�h���ڎh��֒�S$9Uı�݈�����Al��H���ˋ��2k����;�%����֔�J�=®=��������,sUO��پn�_հ1W�c5j��Й�
��]��ͪ�/3�>آ ��dl�s�Y>��jy*�,���9?�w��o"H�_��_],:�uH��/(��5������Y�7��z� Z�-������u��$!���;�6%v�	?����1�bgs�rW<�ñ��G��X��g�ｕ�>2��T�Ji�X��8�-G�o���(#��� �Ӥ�[�����S}��T��]G�.��{��_��sT_|o��-t~��W+ _B������ �<O��D곬�� &���	9��� ��L��HO�b�@��DE������S��<3�����&�Q����#ᚵ�:#T� �uV�|����\}����6�~�P�P��3��h�V�9\~RBct���j|(Z�Ӈ�^=�������+a���ӟ��=�rlg���n_���.�5g⿛�fk��Y�bY�	�`�L��=©�\A����]d� ����%�J<Z]��DV��8�%f�hJ���Ҩ��VVDS�޼�tS;s^P5 ��9a��isa� ���iV&2e~tL��ľ��N;��L�E:�(HBXX5^-�x�:7�-����T��n:_pʬ�xbE�z�n�Y�+o�u:pS2Ys/�j�2o�n%��| ����C��.Kk|D� �#��S�	�ͱ{�.*�*��FB2�*�������O����N��ҹ��F����}i����C��>aH!�-o� ���3PP��F��U�O��'�G/�M����<V<5�J��������a�������~�1]�D<��F|Ժi���P9-�.����d`|���醂���Ͼ+Ls�$z;����+JL����aT�$��R���W.���6n%qk�)x~�Ӽ<�T����b�զk�J�fO1%���=��, ����P�:(tK�ss��1�
�6c��q׷ޕ��
p�0 ��f��KwӶ��&�n��9�>�]@�D�1�a�$4ySӚ>	2��y2=:���k�j����`�ȯ~��#h^���G~C,#;�hc\|ԣc�E+����nI'Oi`?����ON��O��"�.Z�LTWV]��9�ː��z���I�,�"���ȼ�LB�|����Y�׷����U?rצ����`�Sʜ��t���j�����dxo�S��K�pz�f��jS?����?f��)��/2��7o3�z�TR���<d��]����Z�Y�8�B��g�tc`,`�S]�/Ä]S�5�	�����]h ��x��<�Ȇ��)�w�����Y�O�4�6�&�|Jx�7=3Q%�f����1?m��?��*	Sœ���R��~�'�:�K�x��<����ᘧ*a�Em�;�����t�(f�'��K��h]��C�v/BÆ�ޗ�o�I:�&PQ�ۍ(���JT��w$Uҝ1r9��C�b:�^���S6hO����į��w#sd��sguoK�W��o8��U��t���FJ�-. &8t��g�07�]zfz탋� �S���"�0K�{�.�
X[��g����$���kc)X�(N����n�
△�[��s��*�V��C����9r#X���U�K�\��:��~I�n�:g0�6�q�Ptu2�D8�G��C��qdz��//���t;�M�z<J7���/Y��F��n������͞A����Ľ�;�=÷�s�
b��+���8p���.yKx�i��Kl�ߝF`����$]�i�J8���(�u,�����:��᦭K�tkM�����]	w;<�ZbHG��{H�.�'X&WK�Ub�w,�:I&�4w��rxE��/ckO'�ﮀ�y��(���Is��bA�A�����ۜ/]S������r��we�yhL8����g.U���2_fIHE���\]޴^ޏ�hU�gڎ�,;��,g�=���	ƍ���̾�/
����Gb��LL���qHP��B���Eś]��'����ƛ0�╙@��!�J�}g'2�^J���3�x)�t|<�L@N�{�ͰJ�妦MI��9 ,
��y0�e�����ո�`���!�bc�X�����2��(����ϚvJ���HpM�g�?�Dx�9%R�+�����#�S:�^ Vg�Kc!t%����F��G� TG`�P�D��_dFT)X($��b�&`���V��T�VX�q�������M�B5AƴKB_�N�ppteY�8ol�6�Ϊ�0��W!`?��uր����I����q���89~1�����LQ�X@
\��{���!G4�_� �'�(��"��I��2d�'��ڔ;#`�C��ͮ�3�3w������#8CEҌh�9�u�1��pJd[,*����4�,��]ղ5�e������/Nzݡ+�^�>�W��84��^`$ĵk �m���*US8���IE��TQP��/3}�$�'ʄ^�pd+�KZZ�gKN7�)��*��{�S&�`7}�Ac�
3��*����Θ+܂�f�=b�9]�6�"\��g����}��xSx?&�'ސ�9�XՏ���e��X�L�EY0�f�e�w�d�NU�:��$H����=��۶����n0Xi�-1�5�谟P�rT,E"ַp�ô7�X�V��Y���cf�1ԃ�P�sI�q|x(�������^-LZ�TB�D�mk���914xűp�
mqA�Jw����b
z��}F
qV�%��8�	(IQi6��~$9 �My�ɜ�
J0�c���X�-��=V�}��z]�� �X�:�g!�f�4��9��q�r T�{%J�?,�Ye�� �=姹��A
�����J�W����m�o[`[�C�g�k����5�F ���ӏ�z5��_��V��	�nI�U�tŰ@�wj�*=��H�ɟ����Wj$Zv��}T���6�h}�����>J��X;-v��9�N�x�1|��ھ٠��)^��>��w���l����������@��H��٨�o���`Z[��t8�ݽ��	k��2{���������t���k��]�?�����M��h�H��8ls���HZ0���Ǌ���`s�]�d��\�j�k�@9U�ݢR^o !�=�f�q��m�M�뫃?XQc���r����hd�S��B~��)�Y�re��6T�c�����E=�����R
ϸr�W�]1�v 5{,d�}�8`�����+��G�puP�_��l�K�{
�:]�\m�4�+���r#������&�:ɟ?���"��2ר���y�w�O�t37��.��I�u�L�Y�WokDH�n���Vɖ�f����D
�}�F�UVܜ��LAh�w���4����NT;~�3}���.��B�Xθ�Lh�>�H'�k������� !,�U���U��(w��_��ј�v��Ph��y�Q$��t̯�b�=��9˭ԽW9�ux����]U�������~<���\�d�n~<�� }�G�>��U�s��ۃ��	�WagT�u"S�'���T9�6o�k^+1�B�y��I�P@H��or�, �����x�(kEf�����L$�V�2sU��D�l__y���Z�/��dT6��))����-���#16��m��z���z�Q9����]������qgBJ����iR��$~�9x\ �����(�x�� �'�##p��h�l�X�t&ڀ���wH���6ӥtي+Zc��k�H)��}�<��*r��p�O�$7-��xLl.@�·iPs���ŧ���l}����Sς�b�7���]-��4�O?XK��6����B�R8�u���M���:z7���W<P/�y�����J4�����"W��`�6��_� �v�A_z�>�=ό���� \ß^� /�H^GU�鶗=֝1��肹�ٌ�^�+��q���"nx�d�����cw4�&>�X���hb�4�:���ɩ<�^b=����Uu�ܲe�ʡI�;��nh�"�E ��^&I��e���`:8��+2Y��|��E� Ʈ��w;�VWu��U�=�pE�8�����@���j���xf�	c[�yV�S��:���y�2Dz똗��_xؒR]�l0�Edb�"�}��3=dk.�H�?ڤ`�X{ۼ���6�j��)�8����u�Ar#Ӹ{�D:;-G��Hu3T���F)�dbj
��rE� n}�s��*��^Uڵ�K��3�>p�F�8b�
Vx�"�Sկԣ��N�����i���t��!�����[�����jk��m`�:����K<N��y���2
	�<?��n{��!��ôz�V?����mwۙ���^g2V����yxN�^��i�Hib�����pW��|j���Q<,�a|��6�3���`�:n�[�X�S��C�Ӈa>���K���ݼ@�Aˮ�b@|ԸP�Z��b+դ�Bx`f�f�5�g92%�f7�������,k;#،��/�ב;U�KV�X�eK��ד�JE�n�n�^ׯ�l�o�$�$�'��P���w�t��ӒY7Ya�j�����1�zإ�G��h����b��QO�H�䤂=�C�c)\�����~5�߁Lǚo���_�n�0�a��T_���d���L� ��>�� `La��V����7�0�y��VvI�?򒴎lJQ �k���n��nņ�hߢ_7㮛��ݗ�����"y=���7�#�+&I[1�K�^Z@��;�x�1)�?�O��c7욧�w��Ug$T}��):C�?8����R��]������|��
�`V�O�e_p�'�vϐ��������N����dIܖ�Q⋇ f�4$��s5���D��;�N zm�npJ�m$�A>6S=,�ؐ
P��SD
�
�A�J�d��X?F	��>m	I�S��ѐ��RG������ ��D���a�0Hɚ� �N��TWK��<MP��dj���e�Xg=S
�v�1���%@���@^c�:o�����ъ�8�mV5ya�4}��?98,s�D��7[B�)%��V�]�<�s���r����D�����zr��z/�H��IuW��&��J��8��8#��M��<��-��n& �Hϵ��k�]���X� ��x��j�"̮���\?�L����b[�J�Iڶ4�nзf�����'�+�����,��lhIM0��8�)"�~��9�q�Q��]CC$^����2k�F�=��'�2�Ř�7ł"l���(��;B:V���[	6Ո�{�c9��h*&��?�5��5�>��c�����s��h[l2P,�zd[���J�#^3�f62J�'�O�6���Q�F�ؽ�=ྞ�䫂&�t�.1�w&3&���˭���@4M7�3ë�����fB�H�k��:�������!��2yw�zv� q�w�X�ۛ�F�/Int�5�^��g7���,��/���2\�*P&KB~�B,wU6�|�V#�����F�4t>,gEOf�`��(*��čj��n;^�w4�*
.x�/�9gP (���(8	�����������>/���G�S�Jl�Ơ�������;�e$�R��I�M>��R�_~<��.zz�=<��l�8k�hq������KZ�Q�=�zTLsaDlZ1���ig�Ɍ�]��T.Od�}�Q�y�N1�t��ƵKā6S88�eD��U��["4(@�����|�PC����͓��N�DMC�%�iu֞��@)	�����"���7�7�\r�Tan��fTg5	�%��f�R.p4���*���(/.5����!2�y�M�~c��"��T���%�'0RM���4��H��������t�Ī���ӑ��	N����s"d,�uPO�T#��4��iǤL/������ຬ��u�б���
n,89���*�W06�NP>��$�/���kt�@�`�h�#�.ݾ��F�j��
��Y��S�Në��fh|:[6w�s>̍���U姉� u��Ó:eD[ϋf �y2B�'�o\3�Td�Qꊚ�T��V�-��8�"���~��B<Ϯ��
=�D��7ٕZ���"w��O_8���y����Z��~����Ğq���(���l<�c&�X��:��9����P�c�i([��*Y?,Xԕ=�ʾ�>���/�y*�v.�fQq�Ն�X�,�s�%��ɦ4q͒������})wh��$� ,�u���òxBѺz��ǂ���2B�c�AE�r#�9���" ;�a��y�6z�ki7��_�@��d+r��Q��֛؉�O"��l��t�PW�������S�P�MU~ɀ�g��о��`u�*�Ȅ��S��Ĩ<���F�?ʃ٦��~?a:~��5�@�8����N#�`��4p�ӘJa��l����ވ���e�����)d �~� vM)a�F�X	��ƒ��̥�_����ѕ������w>����JJ�+��+�j�X}�M��Ǔ�/�9�F���=r�z�s�ET�]�@oR�:�� ���x&i���Ҏq>�_�B�n����B�Q�m�u�*O�2�Z�̩�x����f8�r�{XrA*�(T����2��h�J�͚��x~芦|�,�Z��J��BR)SI�	%����%KD���O��OU��^��JA;A	��;�����j��b�j\`��ʭ�\�[,(>-����B��?���W$Ax�N�Dk����'1�p���m�:^8G�FÖ�j�����&�3K�ظ~�|@ot=:��M��WQ�~�����L��nyf�}Т��&���.oKਨY��5Z%Q�a�9�����CW� �S�8�� ��U'����$yz������^#l�:���֑�#���q�����q��&���=��#�~���CC��x_�iY�Z���~a�������Uxr�a$!cK�<T:�h��F�y�ɻ���w�������J+e�bu����LS=�f ������_����]�fo���J�a�S�n��o<��CQ�{�br~a�����Q�T�o6rӷ�#�M��0�":���Q@D�`��_G�#�am�Nq��KRz�\ϐ^Q�S�0��V[2�cc>P�H�#P}N4u��z��Urǆ�_�1PD������[o��t��s)i����ؔW�nQ���2��
V�f�_��<�4�Y|1I�P�%�����>�vh�����tO�8��s��)�7@2�\�6���� {��������^oW&��۱.6��Ԝ�j�:0�hx괰����]ocLO��(����lO#�y��ɣ��C��PI~��*�۴�Ώ���,��[��mT�#!��)ǐ�h���4.Z��@@0�]��X��~�62_�	��v���$iv�[����1��,K�B)O�i\E�i��ZX�RdK���X�⡑ȉ�^�B���L��ͫ�Y�WVgǰ��{׭٪�A����UK�_�r����c?�q��ws��iU�� ���ǌ�BJ�;P�4τ��v��E��;|B�A�3��&��{�8�@�}����W��)'J����Y�t}x���2��Ȍ��!����RD�t���o�y������I�N�k�0��n��DL�}�6+�%�S滤�[��7P���)a��	�5��s��3�}��O!O]ta��!vk�h��ќ�Z�o����Y���]~pΪ��ڽ�����;DB�	��#W��x�Ʃ{��2�3�x���x���H�z�����r�pϡr�^�2*�ŉ�d��y"���I�"�:�8�?��:[a��Ž �9/|D�*�\BA3��HP�w���?0�Yړ^��Z�Hǁ��9���\�?��(J:�sA�D�(dޯ��z�ֻ�ˌ�b��=�g����r��b$��}4�3����p�R$�궿�',ӥ�Xn���/tB8%�;�M�H4��B�n��y�������O9j�7��%�a%�LI�9�=�����Sۖ�ڨ~K�|���F컰[�~_
q�{��4�aْ��e�펇+n�]�tF��%�8O`.
�J�T��ׂpM����r���Lo,����3�>���v��x�b�S����ۄ�Ԕ�TH�ª���A���Y��}9�+#$�ׅJƑ�Zf .ٽ>1bdߦ��\j˂�@�*I���y�|��H��{�x�\�>���tͼ3�� 46I�U��f/��P�_�#��B����Wa��BG��4˸�y���$�Ёk�����ˮ�^�Ճm�Ǚ���6p�W����6)@'1����&�l��X�%�]ET�K���`�rUD�ԙ.!愂�".'&m�m��mv(r���/�}u4��1�]\ȂWθùL���U��d䨡7�yPr������&�).g+7�s�ʦK��ӏ��R��f�T?�>x0�|�)C�`y�].V>MX��L�г/���§4��F ��^^(9�a�|ɫ4�NP�#���I-{��Ŵ�h�U�)��Qof��[S���Cw��	:?�!�R� �zԪ����������oV��~��iL�3��	���,nfm�_�� ����&J�S�t�JW�}��=��h>�^@�٩����$��;�$2��0ȋ�UŗP�WW=��^����1��-�v̸ȴR.P:(n�Wp���ֽl�A9��.\�x�l��^a��}�����u.��5Ϥ�p�/{!Ԯ��'�i��n�w��͏�Ov�t`1H�?��sұ��|u�E;	݀����Bv隙ٷ��w�I�������я�?�gY �����Xq$��*�$>̔-��:а��մ�[��L¥%fY�:�c�D�~�O��3��(�E�#R��n�KzXt��hK���B����쇍;�5���G�~�;��0����E���1��w(A�LJ�:�+��^�N]*r,��ev:q/ҩ�����h�o����$PT���l�Rʗ�m���UEM���MB�6��O��2��`l<��Ȕݺ������b���p^ts$���b�|��r���7ڎ�h����0�lHq�����k������[j(s.F�6݇��g���'ݎ�Em�C<~ڱ٢�i`�z����fr�(ף���tc�Ds��O#Mى�4����B��B��A@���ͯߔ�=�	n�����  ���#�����w:���\,O.Yw#`��7F'�?�Ǽ�6�[s�O��p�pDk�h{w��MuV�	��E�pj��/���F�����U:�Vʾ�r�ը�ecY&lTbQ�ݵIR�ѿ���U�)����O�F:��wXs��U�a���ʙjR�ۗ���p]��v��6|�7�C��	��Rt����#\_/�1�>�������,� ύU2�)��_�����aFz��iƭp2�F�O�������T��i�f��BX��c�ݔ�^|�܄�>ig͊D�\�M�q����y!L[�ܚ��=o�&Y4��0% �[mR)f�c:�B�ZT<�V�3 c��	��k9����R��G�eY{�UA\~�Fdq�Fƥ�*q?h!���J��F�����}'N֡����t�q��]���2DTS $��"-�uG=��4���E�+_��g.u�B6b�ED�����}'y����>�c1�8�,�UʴM��c̼�[��<SS��mx��B-�����T��c�P�[ɸ*���KS�\J;b�_;�FV��x��t�KX���-xi�u�桅����E��)�H��/�]���os����m�Z[B|@��/k����B
��"���*y�������y3�	��	���������G����1y@���p���Ļ;���i���e�#�{�}j̦��
���Y2�m�8�) l\7#�CVX�v IG��6���%���4�i���p6I6S!"-5�x��9~б� �[[tѿ�-���X0^5��a����%�¡& �^vc�<`e���Tf�l�t?"!�A��h��-�K��I����LBZt��0(;@5�¥ÕLm��`Q��m�~�S�=�Q�
��z�$�/��1ۼ3�~}���`"�G�7s�d��_
�����#�"�KP}~.ߟ^�"bL�1%��}�/��eޘ��K�.D�g=�*����wy������8橱��ֽ�knw������2ƌ���=��Y�l��^T�R߰��n,�rQ{�T5���a�ȇ��ơ%� |iq�^��gfD=�D����oׁȈ]�'��$���?GZى(�������8([�=��8���V6r��!>}�)�>n�r�<a��V.椞u����5'B�o���>hO���+]g'���������K��)8�,�c�L⹎�.�o���*�j�֪G�f%!�΄4�ӿ0��iAk��cѐ7���}@s*��c��Jo=�����G?"�2E0:�eYK1�X��U����E.���"^p���+xr�O�R�M����tȪ�1�"bw�<U��i~�R��U�d����i�,OF8�2�m1ڢ
|�RS�3A�~9��z(�+�zz��\�x�r6�:�G�g��҅��)��2T��+��kc|c��i*,��������OК׺��	m^z��a���-�箽�ޔ�E�C�����N���Ҹ#h����iB����ؼ+����vQ�^=/�7�k�:�/0�����s�s�h��o����iX5E�'��y6B�R�x��߹N�>f��!.A���֕73��Z����Y�C���D&�l9���5��(�oԚ�^�)�i��Bn{혬"ԥ�K�vaO-���&�I���`���^��SQ�>����)'���+�4�����݀��މ_L�oo29��Ͳe/u[��ɨ�7�\�z���Wu��K����sУ��\��qd����ck˼w��yH�:����B̣'�x��q�`I�^�+M@&o�yt�\�!M�%�t�d�7�8e;�]�(
k֢{QrP��F��H�GɜϹh�zgs�Sy'DZ�s�ڛx���V����Rt!R���߼���op�K��t�-� ���E�zD[nN�b8)�' ���!�-)S����	Ģ��%]�T����
���`��
n�-�u�	�J��-������7n1��;�?������8*#셜���qWؑ/\ <Xq����	�9t�IVo�UQiaH਼���^���Xa����=�ok5mp|={��cG��W��*�A�����F �`�!i��������y��n�� Y ��9$�aN@HH���f.o[�2�+�±c��F�\U*Y 8}��Ha��m;3w�^[^��\��py�:˚���A�s�C(.^=m��L��A��:+�J���~b0�9N�C+�l�����`ř��B7&��h�6`q~7،��.�ϧ~(�S�#5y)8k�N0�	��=aՊ6�����xO}]�.o�N�+N��T���c�+�&l�7�~�:�����=��U���nƆ �9C���C�yP����#>0��[@�ՙ��#�=�9
������F>	Z��J���^��-ڴ��H 5��L�V�k�6c�ܼ�n�![K��?P��KW��V��y�)yE(�:9�S�^VG'k�E�n��Å�zٱ�2G���aC8��`�-,�4J�m���	ٞ�]_���V,w�W������CF#� \_X85k�+��a3��/���C`�(ndS�c	��P��KA�D}��=?no�9�jQ��n�.���NwB�w�3:m�P����w���ݬ�!��%\��NvP`P����x�ĺq}���c�\/��fjo�,�c�=�d*i�q��1��C�ūc�v�ӧ��?\:���Ga<-Ng���I��k�~��O���#h��
�am�(FH�� ��8S(�P�D���Y���
�/�B����2g7��xH���o�O�^i��~^����S���0z��K<�7
eMi��U&�@d�L**�����da��hI�����Z���	�S;�N�bUѦ�,�Aa�I�������"�@,�:2$g��g��`0���*�j��&n��F+�����m�)�>���WU:��WpU�m�~�Aj"�X���?��S�i�>�ɾ����������3y���+;� ������QlY_�
:�la��P���$qf5;y6�x�rqݾ �v�d[
V�?8��;�s�ǘ�c\u&�(
��G�_����ȧ�H���]3��nd�}�y�kՅ4|<��lu���4�\���ʲq� ';RC�E�p�ȣ�x��3u���w�z��s�<.1��o���r�,��"��� �Z�V�q�ӏ h��Ņo����;V6��<�n]$CtL��p�g�aWnڻ�e;�l1�ז�I�?!h�	���Ws!�������cm���DG���5� �^�VO����[B;��^�r8�i��)ƃ�1R�O�z�)�~�ϭ��$. �70�SyҤ{�D�n��ο�^���eN��v���q�i��J���f�������*.-̱h��k�~�[�M������uο�Q��#
v�׼��h:�b�F8�/ڮɦ���G�t�
`���� �K�=ˇnh>cO$1ו�a�4-v3���C@ߋΠk
X�-IT�.J����z��:���%�ps��⼬��� �o+��b��Ë����;�ظ�uE%-"XS�����F�X� 0�w�#C���C��XFϣY���#�� X߫���@@`�A�/���[iB��K�ê�����㇚�`O�Z5����ǳ�h���1��뺬vNR�	]��K鮟��ǅ�U)�W�3@�
#A����� 'Y�'�� �W'��=W�\����ٹG3(��$#���w�=Y�L0�a�c{B8馔`3j������ts���L�C�w]��P���Ͻ���(�vx=�8����-i��k�i�q��v!}��=�Z(�<�O.I�6�U�V��`.9���
+�S�X.�����>*�.S�y�����f`h�;$4Į�h��(�5�;wM^�Jd⬗���t� �Be}Z����]ռ���eﾭnh�T��� [&��C��,����Z֛O9��Iw�]�I���o�y�2\��
>�Qm�D�Q/M��P�8�	��3���@��\P4�X�
'�h���3�S��n�2����hD�w�V9G���yp��\b�h�%遛�R��	���ݍ�*w���B܃:�\ښ��~"r��x�G�0Ώ�!xAG�Cپk{���Ÿ���Q��7��äF�6F�S�_�~��m$=���$L�<�ʌ :wr��x��:V;!ݎ��
(����3%Lo¯�"Kz26����آ+r���� E�JstO���#�����J(�:~�7��� �͇����w&��vqc�O	�O��hV�im�XSv��g�6�����R������P�����U��7�$N�j=(l���q¦��$�^6�ľ�i�1Z���+x��`��䂶�<�F*�D3�$�o8��AZ�Ue���o���Kal[�!�=n*��>c�h`�Ö� A�7��|�5זx^�ng�c)����Ԥ?�~B��Z ��hA�|��Ҍ0�H���0���;���Y��;�k&ˉ|��C��zK�>Iw�d��8f��WuÃm`���|�s�Б����>�e	h�/C����a����~��W�AH�"-�����am�N	��p6]��_�{���[R���sB�]/
�OÒ`|`��	���e\����PĈ��ė���wSa�Z�st��k�L#�|IA�(���<5em&�ؼE�0�"�P���&��u�0�i�k�G�Y�9���*z��KJ�����z�D�b�md��e�Rڎ�cc��f�\����� P�9�r�����ͷH�y������W+bC�Uu���u�������Y3����gh�ꤪm������p��Ȧ6n�D���0d]h����d�X�T8t�-�}L�!Ŧ�j�e�RC���:-f��Mᎎ�\�,��D��(Qi��Y�D�T����%��_S�-h�lF��8��/��PEWv�<�Vq�Tr�>A�?��7�nA�B=m��u���?�K��p�,��Ms��a���oP	�@��0�?Z�j]��ZJ{��E��\x�h f/���7�'?'���t�V��8u(�0������M_|��o��u�l�n��W@��K����M�w2��磙�O#��P�F��2*"]��j�OQn�j��([	�(!����j�0Hא�짮�C�}�]8vCB �'���	�\S��#r�5�h�S+*)]�/��y���h&���#Y��LA��>ą�z�������+~w���*?�^������$͜��;��nl0  ei����9��=Ww3��(Wׂ��\x��Ƈ�1�����-�9J��'�(����R��`�Jn�a��
&�)�=+nRKF�QX������<�fZ�h��f��+�A���_������W�H���<��1�_�,d�^J�ܠs�=���U��3B�F�9e٥(�j���kM����Ô�f�<�_u�\�!���؛5�����G)�yzk"N&��{�"7�+'����9w�v� _��(��$=I�za%���u�[��[z6/�4 XM=���H�+U\�~�j�Z�k�׿�V-�h/�D&ΐ�����W��e�$w��k�=�&+�j��Q,b�ʥvR��Ow���.���%xD<��D�5L�� �2O��D��"�k��-��Ě:_U�7�*�q�Z󜪿��nkS�+K2�pK��ί���4�?��ƅg��¬0M,j!_1'�m��rU;���ޢ��@���S��6t��g���pМ=�������lT@����	�=��
�H��+xH��!c�
�v�
�1�770)�0���D�V�Ȯ�_8w�x���:��5��R=����[(��������02ai��~�}����}p��g[
5���з�D7�� �\�ZH�,�jط�CQ�+�����!��D�
��I�B�����6bH�/�iZ��Yx�!D�'��]s/>�8�]n�&ȗNT?u�ޯ�:E>>�	g�	˭�7��j�nb�!�Qϐ��Wh+�b^E�
t :֔�S�t2�˝&R����T��7���Jc� �Kﭹ|��qih����IE����!��%Y�/2}s�*����>��-,NZ�e@�r��@-AĪ�.汭��&�P�A8s�Rv?K�&�*'�}c�]���@�˕h�E_: �?d�(kW_��fw��d2D~O�j;�/�J%"H�-�'7���d���.\�]6N�����M4	�zKާфH��f~�M3x�H���̛<;��AG�>Ce�{Wޭ�$���Ζ���U tY6	��ܪq�P�Z���ew�<ۦ��a�$�mA���p�ț�!)�xqQ�j��9-̕$��ʟ�]�G�Z8���U3>Z'G~�m'��`�C�[������Ү&̚��
�2sO�V�f'�D��V���g
<��rQ��q���ț���w�SQݑ�c����=�g�0Jc\˛���L��
�~ � XU�j��;�C���������ʆ+���%v��5]pΐ�}����y�E´+hp�{��m7
z��n��+p�MoH�ř�I�>Z��Z�dtx~��(�������uɈ�O���ttDaT�G;��� #X|�l`x��oG7��c-�{{���R���K��Z�A "�@�f
����#-��w�AzR/�M�ݰ�RP���2"knsUçB�l>8��[��ױn.Y��NNd����I�,���Y� ���e"[�=�54o}�_�_���1%s����{���r�W���1��Z�Ɲ��}����Opb�46�1Q��-�H�p2X ��<�0 �"S-�{�56 ~�s�#�����6�0�7�������Je"�D�s5�L�OP�/Cb�3�����0 �!0�y�zjf�	55&NHPA'�����5'ݜ��@M��K'gVN����i���B�UU��L�P,��r���R��U��_��kV}���ӕͿ}�- Ꟍr[��|b�5�I��Ȋ���-���5��u��^�%u��LVd�/}G�>�B}�n8S���hנ�&�����koE�����)�V��C����A59��g���N��j�u���g�q���wF��d<ѓ�c��d%�}�����K�k�ÍL�l�\U��)�V6.� N��?�$���A0�>�Tf_[D��rl#��h����bW-��Fί��˼}��شK9V��b����mZ����
�L�����V�.'���!2��_��@�62�������4��1���yAd&� �;`@�.BKNU�z���q�Ζ���?���nQE��]����D��U:V��m� �հծ��G�_��+l�5��ֻ�2�
�Wp���(؅Yp�&���\��.�z��΢���~.	.�$c�ŪHW���G1B�e���[����E~��w�3�+(���RW�0<Igq�p�<'|Loɤ�s��Æ�_�G$6C�h�4fUE��#
�7f��X����$��3�8�|��{f��/���j�U��g���2��溱NCٽC�翯����hK��[��җ�����@�����^ȶR5f1�.K|�����Cz4l=3
>-�����7'm�$:4���P�_��;��<������d������k�$8�=��YsH��U�4@�l>L�j��W*���n�dа�q�H��x�J�y����
҇�'b��Z�`�or,�d���S�q:��ҵ'�w֝��6�����?]�܄'�D��HzzՓ,��"8LaS~��jU��T�D���.7{^�&��CQ�ˮ�V��K�5��D����t�ܮ,�����$rگ�	�e,@��mM�,oM�	����3BVo����
�w���鬴�z���	��E4�0$2e�Y9|�?�V�_xN��C=`�g��y�h���{t(P�sm13K��i��-b�	�H=�l�^*��,�l������7I(�1�V��e=��}D�������nav3�GЏv;u�;�XV�Y[J�`㱅;������O�H'��h*I�	+G=g��
H��<=l�V\���P?���.������������ҏp�rG�<["���i�	�ݠ�[�vd��6�3���R֫�~j�p�N�#C�)��)���~�h���.�����w�6��Td��i���� B��ϩF��l��Ȁ҃=j0���Lmfh���Zxݥ_w����[���rB�v�?m?��o�߸M�T��ʖr?Ѣ:�l�܀�Vv	���*��ЕK�)�8���Z��G"M�6\���1�E��TƦ�	#�0%4]��An�j2�؊q��R���b|��uR���'�t��{���*��Vz�������y,,%�î���7�5��^Y�Qﶧ�i_S�����l5��Iq?(����pRs���g6�<E���`Q���+\� zB���rNqor�@�P�6��ɯGb���0��R� ���gR4�)�Ż�\-e␺+��-tԊ�4p[�7���'��D-SCB;��yp�(+RdS��H|^F���	�����¥�@�e��ԛ&���-�f[��o0�-l��p`��D?]��D�>c.��h���Ke�zY��чG�hp%�ڄ�|QhD���O�iX0�F5�W@�T�#f�*�큋�:�FN1z����,J9�-u/�6�+P�� |�\�")2���a� *�4�&���D+EZ��� MxbD&.��A��=
'��h�\i�_zք�f�"M��3��d<�,8Q�N�Y��p	�q�>�����O"Z �c>�L0-ޤ���ՙ`��R�/5�<o���~��|I��T���a�� Ӂ���?��K]5\��M{6y�	�`;���vOyB��y���w��X���N���2�Pg^ڤ��M��]ڞ.2Q�ؐDK4/�;& OA�-�9_{�A���ja���ĥ���P��E'v��g�(��e&D�iMV�!�x��$  �Q�Υ��*ʭ�����!�JMI�[�3h-���$������p�2am�FSB�AV��0/��Wo�0�R�}^��H�3�'Eyr�{&W-g�+��>1�s�E�+�I�U�>^,�^E���Nɂ2W%ex�r�Д$�!d≻Z_��ZWpEn_��6��S�gY[8�����K(��ͣ�h썈'#_l T5���4�!���B��w���6��� ׂE�NJ �ǩ�sN�y�h��@�t���Ih�o�}��꩹�-�ܬ̠]Up��Y�.Aʴi�5���P +�4��<4�*�r�g	<�TZ4u�jm[�	F�0Wݠ ��ܫ��\(J�x�����_��;�ʹ= ��~���Tw<h�D,,~�C�8�8�o96>}�A\�}�ܱ����o�4s-�j+ZAY�h�B�{Wr���^�|�y�� ج������,�7j��c��-gB��݇�C���niTc�|f�Kiu�pN{�1�O$i・Y��K��?f<LߎHե�4��BQ��Zt����+�k���B�ef��9�KO]Wmy͡!��QZK����ڵ�	����?vn�_@۶���{��ؾo)�Iv���ܩ?�~|���![�P,��1_�D+~NOt/F�x����y	|��$z�v.���i���%X�d|N��`P���#$�U���q^��R���?�.�=�󽙆E"�
�h0\��l4kٟ���T��<%�h%�ej��U�)8�e�)S��O9 ����7i5j�$_���̴�p��G��c���<��I%���I��Ə/MB�=C�����Ψ �	�סr@�D�"���U������u�N�.wTQ���[7����K���ɔ��XB	���dv,��� �3��V��/���IG��I ��l9��|�6w��Oш�Em>Va�>V�A�+i� =.Axa��i�}�;߃P��§M���N���H���2��'��"�v��Thc���EE	�i�wL%��o��n]ܤ����� ?�)�X�M|6���챯y��.f �1��5_����SCy���q&q����}�zw���5e"����F2k��'�;���4>hE�ʈ��������&�\���F1CĠ��<����I\��<t"��32���!�E�!��Gn�)��ȧ��ʓ������R~��["�_���_@�����58��5���H+l�D(U-0X�gEz#X�_�{C��l�V��v��X��L /�/w�o6�����}�h��� ��B��0\
ͣ^�J�Ƭ�����E��:�	ծ�$ӫBĞO�
�)��HVMU���}�0U�=�t�J���y�����5��!�����V��eU��!�*��B[��J�5�F�*���i5幔��jv��.�L;4=��m^m噷g��XWFn+[�/�X��]�G���M��N�����K|�S��~*5�CF`�A�Yz<�8fH��2��1+^����c���+�T�Ǌ}�%z�����~�O�C
�����q���7Ɍ~��ZQG���~-Ж$�Aѣm�g�v��}�"H4���l��g6_u��w"�Zt`����j	'�*���FuyZ�p�-v�҆H���w���
 xs�Bv�#(�a���p�R�r9_�udA�3�c�<��$L�$p$.p�%�d|�y�3���nI��Uݫ����8+�BN�~�1h �����e 䢞g,�6C�A���ܥyy�U,o 2�YjW/�f��E9ǟ����/t����u��ȨL'��fs#�*���>�]������`��pj#�&t�+�P'�84G�ʔ�L@�$6��L	�� ��r���#���c��4��H��"��fBg�?�^(H$��_��M����� ^�""H��C��V&�A�L��Y���a�9������V��=��,y^:������܀2�OM����^��Ȃ�zob�K,�o��̱M'��Ć�@Ҡ�_�`����?]b�����E[���i�:�{7\���82
~E�F�/&-D,\�7��ɘ${�"�s����O����{#t������(���4ʻRJk�t5g��Ӓ'Vq�σE��7���:ٛ;A:�`�k�����R&��Y@T%��nk�@G�.mM���꼬
�H�����N�W�F��?�Ж��}�6TAW2�Jx���rm;` ��&���{)q:*j,���.40�y��O�4��}i�]м)�s(�������ɑQ��Ǳ�e��*.���X�I�/i#l�#����]�B79�-L������R��/������H"-hs�?B��5�fw�/��{J�V�����c3(>��~e�@���G���Ɲ���0�*_;�~@�5-���>	���������Z�\=���=8�e^��џ��w��n	�ۍ�0>"c�d�[B
��F�5��޼gї)T �,�zI�Ϙ�-��6;LB�PV���"���В0FT�T�E��d��J�X;�:����J���K�ED�5Ea��<��v@I�(#2�Հ��V���Rz�t��P�E�g�{�en�!�J�3o�QѰ�<Lb�,)Ӗ�(�~}��g��Dn�����F��	�ɿeI�_�8��]��w�JB3��>Q94�T�_��K���t��D%�%��ČA��Y�V��r3;x��dm����V�[������mZ��p\��hO���>�su>��L�eWW>���M�)�Ter�6����! ��U�Wݸ"�MJm�5R��/�+}�����X��.���q�^�)�57�~�a�IH����.��	'Y2 �2@�B�mδΕc~x���=�h�����Q���g�ލ��Dݏ�u�u������G�IMe���͊��7�WY�1���\�*�ՉP\Vy����Pd}P^��P�8+��?Y6�#ρETu����1���3�E�z�d��~>����*ۼ���
�|�w�'`l���:g�E{�O�8M���r�U#����M���Y��:�(9LL��.������v�y��>��ﱐ6���4ړ�n.�� �H�R~eJ�2z�;/ˈ�\t�+�5��W��x�]x,�n���v��d�GԳ&���0���.0@]�4M'���3L��+�<z�W��*h��_�yh���)j�?�<��7����&�nm�߮DP@+���?&����B_�+���M���V
��>}CY�;T̹d�ˎeaD�F������S>�D����s��9��=2��H'�)sФ����<�T4M�G�8ٰNp����mSEkxlS���h�
1����{f;-��!�t��O����y:�> �����*�q�OrL�˻���1Q�oG�����P<)Y�H���� s�f�(�Zъ���
*�X�p���hK���+W퐤}@��'�h��}�8-�ohgq��z�LI���<"����	
y��U"��*�^��?˹��ڧ�q�^�Y.>�e1#��ŠH����o#�G"�vc�rf�g+S�s1Q4������Y��=1K�m�6w9���p屩�7���.w�����5�ɯ]g_z�F����۵(u�[8�Om'�Mf���2��%\(�P��̟���)d/��_h��`�g߯�y#�s�P� n@v��b�8�n!���]:���Z7��(����X�I�����&ڎ��i��q�&�H>��GHl`���z&���J��Rd����y)WMn������0��$��?�$�w�W�UY=��N��X�gx�G���;'�~�H�:<��qx3��:.�tǉ��#7��5P�!ax3E�v\�ba3��S��o��k�z����#�O}>�:Pߎ[E��@1�k{$#��A����fǐ��T�)�G������|�SGq����������n�m�1�+�g�:'�ed�f s(n�_�y
C��|�u	d�*����r� z$!F��Y����M�}��v�g*pʸ{�l��[�����=c�:�c���ȩ�Jy���+��H�\Yp�O�+��$8�p��}�S����!ES?M5b��)��|���}�.�:�<J�$g�­��ͦ�?y=���ZD�;\���A]�6wBh�|{���^�x֧�g��W��Z�LM�C�Σ�V�u�D�Y�~�k#p��|A��e�& ���<��R���vM���dܻz߱�UG��p�z�r�h����Y'�6�4�aK���!*�<{�
O*�_�^?A>>�_�b��HNX���ڡ��C7L(���͝*꽡:""mz��7^�Ȭ�p?���6w��~�{��5�*nd���M�b��ٝ?秅\r�ņ�#f��X�x��ƈ��m���H�f�{5H%S"���F�ܾ �����[}�B<�?g������ڏ�ח��� ��:�_�ƕKLv�� �y���`j���nG���R��]��M��X��������N��+Jk0��i��ɿ|���F��q1 �.7���(l�l�v�b��n���T�*%fpx�(��BG��� n�%�i
���^�-�Ѩ��>�3*��+��(0�a�FS�H�$~�ʥ<��tW6��I��P*4S`��>���+Us��ę��A�x�¤��ԉ�.!H�?5~G�I��+b��d������!5�t<��[��ԉ�yeV�sϩ�b꺛i
7�\��8N;s�}+�P���$��H���>�(���ی�jN��fBhI��|4E��Y-!r�b`5���hx#`7e��r���5lv���%��5�$������T��J��߷��PF��J�e�
���C����r��%lW��mge�D+�TD��$�jv�JAF���lsaG��f����^��(�f�*_�+�`E����cL� �YA���w��S_�x�^��h�8H�ƒӶ5\:Q���q> �yEO��/�t����N��Ƥ��U���H,�'�X;�� Ch���>X��&��,p��\�!��c���yW��Җ�U�% �N�qfW�x�%�PI�k9�7�-O!mҼ$PX��]����鄤��0gU�� �!�|��𫞽����p^B��B
#=�)����IH���p�u�)V�f�ݛ�* �(�@Xwщ��w���'5t�VT2S��'6�`!%�,�͖HN��<�B��4c:*w��}��
љ�������g��F|
K���%���I`�G=H/����|��h��TAHtOϖٴq��~��󀫼��%��c��կPW�`�ʲ�Q���n��K�eu�񲴁��`� ��rm���d ���t�=C-#LBEp�0�}P����0?���1����|�0kk��TfO1�Rs	�y�I'"�qkFL�����p]�W ��B��ܼR�n�k���e���k=�Q����%a=��� ���Ł+���a�R:|�zX:�`�z5uQ��ӥ�V�z���N]���B�C?�;����MirT���H�r�Q�й�!֣v-��Hv������.��L��bȸSA�ʎ�8��:?|�+,��@&9�o��`���%I�3r0'��d�?h	Xo��u�H ^�Ý�h�ݢmBP���~��ѤY��,�61O��B�i�:UkķE<���p
��8N��_�jU����T�V�N��y'�:$�lTg�~x}9��#�N!��k&��I+�Fp�
	�<+F��V����z�]^#H�#|o\�����<��@��<
!^&��?��s��2?����V5�D��z�ѕ���.JeC�d��dz�/�7�v�q���Z�B" �թ�*��2�G��C��n��.�*M��(����	$�� �D�uj�����*���6��yH[8rfr*���%�qP�3Ra� ����hZ;H�v�E���$�aݕWb �F(�8��1��o�r��P�����.X�&hף��̞����n��]g| r?�Χ/Qx�9~�VM�쀵5���;5�u�M�2����(?Q��w�\	�xR/G���E�5io��,yd�绨 me���o�~�G �I;�Z��������@��ɝpk��$P�R�7K�X��=Y�����Z���Y�d���PB,,���Qu	z�D��M�>�+��~���Ǔq(����F`g�p��2*����6��z�
L��8����/i�v��k�[[Zi�L��+!,��n?(�|�I�W6��spҚ������aF3�=1'����q�o�&��$I�մ���G|`s��3I���e���\ ��UB��������}�+c�)5h�c>I	�a���nE�j�bwc^��߉u{D+'�?Ŏq2�ҭ��ڌE��t�-��0�o�9��.�9�2�(�-�s8H"�F����8��\#�E�-=��Po"�?<�[q��B9F�������'�7é���BdR}�;%�/<�LS`*�w�pH��n7E~VW(�Ny�}%��h�E�(ϫ杤��pK�^�|)L�i}�*7�d��r��0� �ռ�3��D��ֲ-��
���N)²g��{}��8��h�t�ϬO��/����E�l���,�-i���3?c�����Z����.�Nz/S���cM	Ձw��o��{����A�p����^_�U�܅H!=zvČw��)o3��c)����I�O������|�������=�]O��Oq G�#��c���\O�D��!�o{�E
u�"�Di�, ��&�T��*�p����7|��{u��P��_%[Q4)�C�;�岶��н�� ��-K(
���#���'a2e/�+�'W�G�X#��7�K2t=�wf�G�?٢ M�����
d�M��H?زR��g�/����L��n��P�G���ե��+��������r��a+O�?�L�� 3�":3�����x'�RV.`IV�:I��,5��Y�<ۓ��f=�_�i�*��whg��S���*��A5CEVh����h��6]U�<z�ΗK�Ey$T:圞�,+P����+�(��(��̰�-o�m�"e�)�Z���H�1�R5��"���?,Qŀ�=��^釭��VvÔj1�I�/��׹2?E��6��7"^�	�ʴ6q/{��q/��� �D�*ޮ>`.�G���4�@cWuS3�a��'����e�hrBt� ��}xϮ{�l�tk*��	;{����r�yM�اcR���Z�J�3A?����3I��^�)"��q�����I®�=��51D?�G��M�IhN�zCvԨ�>�="Ƶh�:3F���I�D-��սڋ�0ބ�c0����<Yĕ\�l@IZ����>)�����%!:��cSJ��Ӧd����Id#I��FU)�d%�LK�����;�(e?��jB/v�SL},�%J��v��Ԧ�
Q��Fс����������~��X����M���WAσ��A�9$w�����sR��lz2,�9�o� �\܌���f��������k�i^�ԡ&Ul9�-�^�*K�Q�C�9�b��V��O�!,xV��N-!6ĳ4�M�]�\��/MK�=���vXz VZ �E��'�L5���	�)؁����D��7F�'���Lgs��-L��v�#a����Ѯ	b�`05{��UT�����MJN	I�^�՚x^��x�O�t�OvӬI�ĩ2��ڠvkp�=�a�����<�r1�(v<�⬄˒�Ϫ���#a��4��mq��I�m�3��Q�G�W0.Y���H)����3I�K�4$r}�`^��P6�+�\2lB�Q=����2�Gm䯏�&��Up��1`���W�f+ �"s"���t�b_���c�	t�d�]��,7	�VI�v�܏����M	���;�2��I�0#[�ӛLP��W�#>�����9�JJK�h��g��gk��݀��싯W��A��%LR��G��l��k��� �k���p`6� �&ms��r7�_�0w>����w���+.��q��5���ش�jP�f�+L�f��0��J)[T��0R�I��+����U����ihq�M\�?�����;w�^Y1'N[䬌Z�J�j5&sǀ����H�j>4��Q7�.ӭ���Ð�Y������|" ���g%^&���hֶb�N]�i%�MKڹr�aQ�[����.�qty���#�V2 "�X-��]�b+}��^7ZZ���BlC �h�ņ<��Uvm�o �e�x�!t8ۦU0U������'S1qo���D���`D�A�0׎�v.�dA�7pWxTC�<|�!4��]��{%;&�[rƂg��Y�*_?)Ëvk
���Y��Kp?1s�+��z�����^1g�U�h�4.�zD���*��kc_8�zЊ\,�@>��a�S�a�b#�2�$fP�}�ː*�%�ƌ+ �y�
C��@ɥ>!�N����q���s{�9J�� �2�6�ڸ����P`���@	����Y�f0�� 9NP�e/0 /M߮�p)��B�O܈�z�T$��>%9)�'X���}�8H�5j�i��H�����W�+k�O]uo��1��ʲ8�N\1���+S?u^�
��(P���hR�5ʥ�83�Ty���g�,�\�8ͩX	���ëg�$���fo��}���}��T�6 ����ƾ��f	�e���8�����v~Pm��5���D:�4�V�-uP�/i`�/��trv�@�H���w�,�R������f��8j���{?��ZzN_�09J���8t�����F��v �@��V��5puy��Y4���&Ԓ17�.��p�o�cn�φUrm�"� �$��Xz�G�3� =Mg���w8ψ��y �.��SY2m;H�ȇ���<��La��T���kMo�@D[��zMt8��3�H��8`O�� $G�#A�D|Jݑ�3�������T��oЍ�ԣd@��S�#�Crk�չz�מŽ�JEo��V&�6�@/�|H*��X��e���rA��z�w�v{A�H.����]��!~�"Gi� �Z����L��)�rU�J#8��夼�ܫ������4�|�Ʊ���|�+e8;>%B# weO���Lm�#���`�6zV2j�)J+V7���rf��Nߠ����}a��4vG�E�k��	�M|)���h��(�V^��:�j��b�B�A`L�O)�HT׉��ղ���/�W��f��\va�������Wt@�{+R-+��Tƛ�hO"��D��$|]�=1|�<�-�_Y����M'J�=�@cf�"�%4L�U2�G�2s̈́\�c��B��4�?�A�E��԰$!��	��<��M���$�"��ॊ> `I`�]ŀ�A�}�.������%PO�FM(P0���2o���'��~E���o,��rj&�t��<Vh��ܫ|k�,��o�����c�l������5���(�͔^�h��ju�O���Yoˣ��dy2o+���d5}�JEBk?�P�/I�����B��Z_S�[C�%i�RN����K�|#reZs(+4c���
Z����7�Z/!�Z�%���&�����a��МA)L�F�P~[�L�"�ucL��r�'ĕL�n�5�U�G�-\����ڇX$'dN�ȓ����t���~@�Leg�����o���n�[�YX�����Á6C���HB,���~�AJ����,�5����y[x��NV�����>�멹<66�M�����p�w�E���em#@I��Oy�Ⱦ�}W�f8Oa�pȑ�Bj�r�UV�$Z8�쮖	���1��W�5�ox/q2���n��ѵJ<T]�?�6��(8De�ۜ�Q'=�1G����r��$2��m�I�=`�v��I��萭Ŗʚ'�7�v>�nd�&�E	��E��9�����A�2��L@��5� ��a�����:w��`ѧ�X��ٮ:[�<��.6'\L�'b��yD��u���f0"Y����'I]G+�mo�w>Y�upޕ��3��$66ON�[Wۀ���+��r�B3Ȋ��u)O��)�p�ҥ\�dYJ�aͯ�_�Avе��j����`S.�$�H|i�I��o{�y}t�.�tp��:	VZ f���
���^�@�N�_i{4���Y�`��F���%驂�Ǒ�N%E���s�_�^B�����܏5�\wЀ�dQ֚{�H=0��\�}SO��1��:��gy�pp�iW9_�^�����]8W������hW0�z�J�W:�7&]���'��X�3cֱ�����=S�z@ct@M����R|ت\)e(��K-e)�%���*����້�(�mǕ𭣇w��u\�|���\u�y���`K���(�ߞ ������g
Ez��V!s�`/%��c�3ّ+�@��V�`�q�!�@�Q�<�߬0��%�����e"xm\(m�z���xi�˫��{���ۖx-�q�"V�&���g��{̵>���̽g�聮ȀFK�Vj�d!�EB��+[�	Zh��
�����n,���͂h��a�mYI��ZB��?n�\l�嘂��].-�#�&BQކn��B�H��<�i
�g28��ݮ�"�3��k���(5�Q��������T��9m�(�y<f�l���(���_]M��������~� t�0�U�5�f���>��'�'� ��{����:�NQ|x	���k,gN6֚ ��Q2�S���Rr��Q8v=]&O!'�8�� �<B�Zmɹ� ,=�!�g��K�Th��9�=m�!�XՇx��:7.�:��\��7u�j�&����Ѫ��̹�K�0��I�UԶ�4�����?c���V	���G;n�6�E���\(�b�qvsO���8WJ���^|Ճ��f+JG���!��ι�:ߵGu=Bu�D&��:-Θũyų�5yc�N�?�����$�c�i�Z�Ǽ��ۉ,����py��7\���I=�%>.Xj�	
�/�&P����;���O''q�A���jmpZ�9VK�x���j��n�ߖ��]�[K�1,��o0E�CeO!��� {~���.�W�����B&�xC�M���쪞)S��\��q/V��W�*۰*@3D7!0���KAR[kZdR���˥#�ރ.��@_�{��9WJ�9�� �X��c1F���e�]u���1�K�"�/0�l�(�Q.o?��$��{D�+�r�5ib�ᖾ��w%��7_ªC{�_o5����'r�pzE&�I�t�ݐ��dc�ަ�g�<�*l�!�-u��vKD��=�C��k>]�ڱ�/�N���+Y3b����a�E�0�o����E������5x����}��6��`&{��:u�=3{
"�K��>`;�����R��P��?����$�Zε���,25�d(	�$Y��&���v�CCV�hW���ܰ@썕�x�LqZ��,�����n���T,F��4T�=T��$��@炑�0�ׇq�)4�Kl��{�w��O�?�ffm�:�D>" 0����޷����V�?�{9���q�l��)-ݝ6d�Zsw�7���O~�y��j_H���r#+��Ͽ�����ß��/IЉn��.�9�����w3�D�˸�0��׿����
�5��ڍ'G�/HO���Ta�����ܐ]��PZ�yp�g~l�H�j��N�0���14�5�hC���h����r��wԇrb�Y���y���H��AS�C
�F���q����Q��+�& a/��󷘼�3�/��v��M�A�
�a�HK������l����f_����k���Ïj�����n��>c�,�؎�-B���o]���!m��h�õo��]��gz�V�>"�ʾ�{� i��A�5�?�K�n��엎e�`,7�oh��}���^�?��k+N��H���S_2����J��m�!W�XI��m����5ǼdK�����o6����щ���/��3��]�7�9;��2[����#(��,Jzkb��n\,�TW&gp_Y���9�%�n��{ɜi��熁��.��\��>۹�+��Zm���h��-�{����$w�󣎿P�j/�</)S��1�N5�im{QQ��gj7�kU�ʵ�n�D�t=qE��;>����غFi^�'I)���+C&�ks�t��.V��g�'A"�ԛ���{[p��5&�`4D2L�RW�O����f�x�6@�_���gA�8������ˈb�e[y ���E�<0ce�'� �_��_袟�Ȁ%�Y+%�76tl&�0����|kN�^\֘���Ʃ�!`�V��j�����~�����M��r�M��o��۹��I�Ձ9����\�g�����<�h�;v I�c82ց��6!�?[q�!N(�=F��|~`m"�_�ɵ[�������T仪�p2��@?o�����Z�i�b ���!(�50g= .�A�Z]���٦Jl3(���#9�禗���к�)4�րv�옯)}���/�������֭��1�Ljأ�F� �W��eb��V0�n���>�ԅ��e:�w��� ԁ��k��Iwy�	�A�^�K�n�H4���1��h�f<����T����-Ao���,GLh��w��w����f���w��GkU��ɿv�z�JA?;*m����w�6���k��u� ;[ ��鱴rS��|��	�!��=��6[�M�
0�D�m��e$����!�v�A�1�+�6�Dv����U�]�,�n�<��@&�3	�f�+.fW�k利��r���;.虆�3u��,D�}Ȍ:H�\w�tg3h�����+RA��ў�`N^��"]�@5��ˬ"��E�� F\�P�����evS��_5�ˆ�y��?n\c�c������%��f!jp�	�琔����� 3?�*�<�'��tD�*��`����4u������o)6��l�R�ґNn8��: �kaҡqj������L�!jǬ�w��rH#X�[q�v���?u��W��?���\M���1# V�Z��Կ
 y�O�i�/���j���3ֳ���tp:���-`16�_��X�Y�6:�˱�1�f��_� �^D��P����eU����8r�ߤ�+���"i:���-<����m���_B+��?Sdh�ňw��>������v�.�H��s��Q9w�PҦ���G�!����ǰ~�V��+t
C�	���%2]��o��C�c��e.���)������t��z��c�۩^��[�Ѧ���N���/N2|�a�� 2L(8���L��U�	*��)˝�M�08Rn������7�W�������s,��=MD*���4�r���@���~��6=^%�#����x;�mC9�z������̭"���2U�x���:5iE����2p��A;{�Z]Z�����s��wb;���C�I�t�����!�V���{�t=�E�]�}���ф�;|�!��"G�ޭ	}�Qq�ٳ�������b6
_O�������-��8�&����(o=���CKZ�����}�W�x'>~����U�=�6O���HG/pr��	~�8B�j�m�M5�Ҫ~^�V_8�)xN^M�e�Uj����y��u#���Z���(;ީ$��. �����&BhK�e��ݤ�v��3[�?�ڔ��t�Mo�
6�%ޗ�3�L��ќ��ii#��@S�)��Y(�E���������W� {�R��̋�<�^l���N�k�bԖ��n "�����6pH�����B�u���>a��R{�� V�a$M"[�]B1y��l�W( ��T�$�PI< �`�R��&�@�#3�
�\(+�*�.�f�>���l�+0ʼ��g0�˫[��H�#q���~Ce�3bbq	ޭf�NI��ϬRo���N5SM��	s��$������g;�Qa�����#�6#.�"�o�dёĦ���Y���M���ޕ�1�s�64	�U4�.��H��Č�MF`� ���P��(�]R�Z�!��y
�]5�M�I��z�J�d����f����#�`���3{�Jc��?�F� �>.�7��;���OfhZ~�8���d�-��!m��? �1Y}�|��q��B�)���k)ܴ����G���
��HRt��Z��"J>�G�yC�9z�igG��C��]-���{@B��q���콞9Mo�\dՌ9�#��ڳ�HN�����U�Y��VA�{�!��7
��F�:�X���i1���,�
�\�[Q�`�mE�u�=Y�}�b�P����uތX�������\�iƑ�>AX�n�����1��Y_��V;� W���;Y��?�>��Bʱ�CY��7n���`^�0G��gU�Y�h~/V�&��Y-���+̮��cF�e�Vp�{"I��T���`�����h�#N'�_t�NlrIN���sQzCG�9��$�x��JW�?׼t4}�IdȔ�&�����ݵ|:./�+@�^��o�s*RX'{�O��`"�3tX�A�ƀ`���x�i�p�N�$wTu�40�S,��(���O����'���@�n]p.�;����π��O�H�.�,��ơ�L�k��K��b���5OT?���)�����Z�e��<�¹}KK�1���U���L�
���*��2Hgh����L׍���l�z������F_�
��E�����6?����p.������Eu3t?_�y���L�q��M6l.ňvs+`*Ʉ���vw�~���ꈱ�e��m�㑒���-?L�S�rVL������:j(d�|����ե TSK�`��F��|�i�q���n�+X�[�TOŔ{���Ϧ�Q��:��*?�Sp�g�p
f�����x	 �`wSMo�1)G)u&7�0�t��L����q6��9(a��p����s�~0.@
ѐ�=��c�R1:�)5��.�>W�P���,�'��͂?a'2}d$
�Ϧ�ll��p�<�V�����YJ��y6T��Ű�-��g�y��/�S'��{����bL
c�ސ�ybL�F�#%�Ȓq�x��'_�n��t܈mufT#H��8}���@��q����׷g~��a�I>z��4��8c�&�+�^�8�I70�v����;*ƻ�e���e���8W%�8u�^X��Ū���.@��5b�
�*dߑ������ƻ�4$���J>�zeH
��?Jù	�O���N��ox��_�.m�^q��P
��%؄��̹#�B*�ù��Cb��e�Ջ�4.�U+�qW��Jqh���g<���[ ��~�-���bB��O^���a����dS�3�b׹I��8v�vk�#������}��c�5�vI%�Q4b\�ܴ~X�����U=��0�-�.27��@�+��byE8<������\c+���}iZQCЄ7�)d�輐,��6.�9��A��d3��^35ւ�"H+ڽ����]�(ԟ|���V���w�����lN�
NYj� }8�	'�Q�\� C�k�ѫc,��6��� ͦQ��/訆f_��"q�QYK�)���M+�)P��k�����R}�O��<Kq]��Ea�s}9����)�_5̥ ��f �2��Q��8�pNR3p	���=����HZ"lc|��3�`\�i'Ic�0��hy���\�'ι�& A$_�ܵ)[=zڃy��wx�WRrw�$���{�¸����Ѳ���İA�[��z�kي���}�� §�.ni����@N�4tF�4���C�D���\�Z#����_7��w�2��	������*U�'Hp�U�4b�_�-ߎ��W	��g�O)黚�7_�+W/!/e\��!�����=5@L�=���X��ز&>�o��$P�שWY�gf97��pҿ��n�N����� �'��ynHoI�w�EIm�u��H;J�s�1K޻u�f"�?��ǆ�:��퀡j ��΢���>�Lw�����PgK�U�$�0�Q���w~86C�5Q^K���tcd�T��@E���.��IE1�_9z^�EdY]�mT��'����������I|Ȕ؟_V5d�vI�[���r7�ڷ����g/m��8�6	��A��bb���"є?4L\����11>���z�&�uf���&���4�q}rQ1��ѐ����:�z��)q���bb��������~`j;�\�z���,��ꐨ5�m4���z^������i�n+0�o(E����)��Q�3��W����t�!xX�7�,.�r(� ���I��Z��@��t]D�������i�^�W�-�8�r��"̝���?�Sg��Tc1�AeT� Q�"iL�ж6}�Ĉ�����֠�=��	�3�c�8���Ba�(��js�=���R�V-��|U�3nz` {'���Է2��8IS �ý�zV���#�fJIOEE�8�SpЬ�U�"c������ڀ;�ȸ�\'�Ƌ�0�\�%@������R!�`ԟ�L1(,.o��)oS	���s��_{�se9o":!f����k��=�>�_#���p�]Ow�h�9�?o1G�l|�� �]��i%����'=]K�nk�6ˤ�����L�z��r����E��k�)o��v���>�(�o�=-{ݻ�9��W3�@�*m@v��;��6S�8����I�D��0?�d�B-�Hf�k���1�ۘ�:/2����1 ����R
CIۅl����ڮ�@��$����z�1��
�����
���!K���`�4uQ��1d��麼�
��'��������q�er`�J���hM�A�nn���Ϝʢkg3�=Qj�ˊ(?���0(��D���	eV�N��;�7l��U�a��J[^�[��V Yr��e�.�u�.�ϊӑ�RQ�.�����o��BI	��#w�[�hP��F�2��Y��V�5�:�$>4�!Z�	"�]�nŀ����.��Q��cU`ʦذ�A��!l%,��]E����jA�Îw1x��7����;�)ӽ��}�[�����l���ȃg����-?�Fb�M��-0DJ��-jg`rG�=������4g��3������ڼe� ��컱��f[�|�����?̰�kla�Q�F�	��A@�0y,��E5WX��}�3p��:=`�(E���m�#P������uJcK5f��X1|M�G� ��1^q�=5a^��2�zƮpcf�7g>�
~(��r��+Az%�A�zs}*����k��P`��v�t�(o��r����o"#[�G9��q?�bJD�p*���J�!�-���Շ^�I�mz�/�WK:q�!)o
|;7ѱ�/Tv�D�Mt	 �G��)B,�>\�ra�q}�q�(
��������bV>!�6�_�/G��c�d&����Q�cj:���j�������L��g�K�ꈱ?4�FS	�,�L��#?�Ǣڙ�l�ڛo<i�F�Y5��仐��2��g��J��'�zؘ���S�g�y��]G�˱�<@mz����Cdљo��G�b�Ʌ9u2��9k}l>N����O�����D��nWHe�ۿ�=| �ʜ��O4sG��}��Xl�fo(���.)m�&gS��ڳº�札��ݎ���g����p7�C.�`�]o���sS����A5��_�V�`U�%A�tIf�Z�� ��.�Q�oZ��ȵ92O����O�y��	���S��bŬ�^�T��a�L�(�kwu����Fչ�s��3I�Ჵ��ٟ:B����'-h�s���M`��l�q�zǕ;�NTd� ���_#[nE�;�qIS���e��A��%�_�4�	6B��G�ܵ�l�2f�mD��FUB;���V��V*�2�=h��`�O�ݑ���X�܎!� ���mR�Ț�T,f4AZ���T�gi�b缃wt�T�|�=�v�ڝ;A��n��x׹�X�j�	y�����Ft�y;h[qۛ��/�������~.�	��@�@�u�ݯ}0hO��o2��lD��BZ�	���2��H1'6vj�bCz���(����4;��P拴�
�H�qbT�h�����	tG��_kF���}o��JW*?-��J�i��
�ڣ�0ɟk���5>+]�8��zp�"��_C���J�	�W	@|=�)L�&M��	1�?9�����iNk-
��O	�}Dk�G;N���=�*Od��h�aO�lp��V�y\���Z���{y��d=v�³�Õ1���?ׄKOV��h���)"J��y(�����0f�G�W����|�=����rG��/��/��˖����_��/�Sgi���DD�����R6i��S�ʂ���o�����	��T����`�n� I�6���{^�GgU�	�dZ�സs�TC���ʈ	&�E�Q�c�z�����v�������T��l/|�ІL�8§AC�������@����\�^�x��Hv��2��s0���߼O��&X�E�}�=n���`	0�+g��3j�R�\��>i��~�v�����[�%��޳��?t�jKq:ۍty ��8Q�Y�'�x���R�����f�M� v!4Nu���p����
uΕۈ%�ʛ��Kji�0����z"l$�r���j-S�
lT���Q��^�QqD���#f�՛@�3�=EI�pwq�D=U����ߡT"�~��A�[�jLH��#�&������6����%~��=�B�����G�OJ��Bl��b?"���QX�ڟ5�c3=�+�8�a��P��s��vY �{R��$�8 iN����j�LO��ef��rl}�ֺQ��N��`�ѐZ����Y�Vȿ=���E7��uPP	���Ul�x��Da�)��++Z��[��oT�y��G`?����+��A���WtN��B3�ٕK��� iܭ �S����0 �F���>O}�8�L2�2��4��'�|�8�������~�������n�X��n���/�,r�R�g:~�w��֮@�i>��|a�&_V�1�Q1���#�a�X��rbe�=\�$u�L����$�/*Tgݦ�H��}χ�Y�hr���r=F�:z�ʪڦ����Qg��{g����#+�0S�"�*�h��m�"m��e��7�*u�d;w�0z���������w��쀰���&��L�^��*�1�u>v��g��Ġ��ͬ!��p	<ႅ�Wk*zJ$I\P�.HC���;M�B����e
jIf�M5^�<�.ӏ��@�T�>�7��KAv�h�i��zC���P�a�t�;V+���������z�G�ߎ����B��֔������]?��Z/"�,BuY��M+O����O�ֶ��t������z�ݏȀ���
%�=���؄���Z���Ø��o�D�a_���;lF%�ʢr1� ����K�t�v�&�xb*O/�6<��vkoX�$���2�wl�m�G2]�mi�ѥ&�A2�W3lDw��f[�ѱ�����H�s��j���JH������/*~i���cW���"�<�e�X���>QB�]�Y3�.vD�U��AW��έ����|����3f�T��˙g�4Ba/�ֶ<���߳9ךZC��w���~Q�\�	��B�
dl�"[iKZ���Ǭ��c��,08����bR�(rHJ��=�˧� ч�*�e@+6b��-dz̀c�#]�Y�9d���[A�]-����=.����jw�z9O�М���B�'ѷ69����eR�EC�.nH���^4��ߡ�<[5)��q����ۧ�j�.���<���tܲ������&��<�Ky������i}�^���ݿ�r�u�ӸFE�`.R����`.>/�*���cq$�Wa��%���z�쎱��Ex-��W��~�)�er��a�ciK{1}�ŀS㗥����Xhj��/q_���v�>�43?�ղ�0�U7*�v�(-�ë�C[/t��R
'��0Kr�]P�R���n#�z���VatֵS�|�����j�՞a�nn��N��`�M~�<,"%�UF�l�sO'�WL�%�BvY��j��]�/�q������W���\s7J�U�H�I[)Őa�"x�0��_"��=�?ɡroe��i�7 ����P}}3��Q�SI�]�B��3��,vmk�>���.�U�f�z�a1�X#X �Gu4�&�v�G�m�0'Ekt�|$�uJ]!��+����CN�.\hO%a��K)�&$.�4��nT�a�o0��S��`�oT�>�.FK�&e��a+u0ž�`�<P���wA3T���5�f�!�>恙:�
:���̎{�n��i���eO���cbz�t<�{{�l0�P_��k��SG�� �?��< p���.�('��m:e�5�_`$�Eǫ����N
���c���A,�,�\�Ee�!F~L0�X���J«8Q+�mΈ#ݮ"Rjŕ�8Js�9���5@��~՚S:t٨�V�N�*�� iq輨���v��2�dl_�����	�%�����z"p,p�)t�8�t�y��<� ˡ�)��&/��Q��6�Q�c[�]��K�y�SD鳣�1Q���sGtO"a�nJ���ix�X����u����=PƂd��i��@4�c ��_5�\-��ҙ�U���W@r��$gv�^o Q��۴��k�m��3���i���(���b��q&{��{�"��������K!�8��]<[K�_�_t���z�T �|Jx#+'S�\,6��Xl[if��r�*��ԀD�p�Qe�flJ��gW�0�a��Y�XO1N����B��!�%RUYJ��Xv5�����������n�h�~�4{�bp" ta..VB?%F�m�����\�~%�քo}/�'�u	6���+29&)8L͎5��vvΕʗ�R�J��<�>k����9т��b6Y��a:�i����-3E�҅Ie(Y�8Z�Q�܈ja��h��\1�pZx��.�{"0s�Sz6V�1 �;�4	��Zw��݊HDۛz�n��rxj!�~W��lW���K8:.�e)~wy����UZ��*N�^*Y�c �"���D+�����$/wy�$��f���@{T����c�W��W�fK$ĝ|/Ͽ@���%���a8ub_� ����%�Us��U��@S=������b��\{S*�_�AQ1���ٳ��2�7�-�1�S���@*`b�pK��)nW`�%����}n�����M��-��׻]��|�m���WPx�eI�wWg��.�r��Tٵ���%؀GV���n,E��ȗvYN�s��՟]��#�z7��x�'�U��s�6���q����7�VJ��\Bj(]DwUgVl��Vf?$��چ,�I5���Y�#�F�&/���o��2B,���a^ ����ʑ��X��]��u��&�Dd�qWC��(r�a��k��]�]3 �:p����Q���\� :{��ŜH���}	���)�P�c�������6����n�nZ7�\⚨��ȭ����6|ˌ���;�j��ce���h��K'�j���%�7����Sr�y��ʬB��e�p�gM~���3'�<�~�Z�#����zq��˅�ġm�~k��ˁ�=}�v��W?��G{���������Fp3�vZ���.�%\w{ײ$K?(�/�xi�/��;\����ߙ�E�Vm�tj�^��~V�xRl�8z&8Q$�-'n}�κE�&���h>���h ��V��ԉ�~�P��h@���R}�os?o�����%�H���)�9������`���Ujݬ�U���ED�"|:��\�~����;P����l7MЫ�S�97H�f c���z���١�9g�眑S�f�O�K?9e!b��;���.����jVY��1G7���'B��I��' �`�0;�9v:J�')^�V��*�J�`�W�l����F��U�����=,~.t5���_��S���Cg�տ_����a����f���7�+�R=4�K�A�[�5�Vwt��0�`٬��������{t��S�-���=��|���d~��>�N�յ叏z�b�WQy�n�(;��� ?�J���ol]�Z2��Vܖ:	��Q��4��%%�)ݙXҙg�oCl�o ����^w� T����e!���dՋ{����3���U]���U\n�;�%���%��-�qiʆ/���ҁD��i1+L#�gn6s!&\�!�|#��I����O}'�jzjD��D���7Z�L�q)#�Zk���Oy	�u՜�K� Aȅ�s�*�m�yf�|����FW|���*��x0zt��΂*-����y�`��=��F�Uϣm���¾�\Sf�4[r��9�� ��G
*��-�O��(���* �����Zأa�\u!�5�	�-�k*� �	/�r� �{֤z{m��j�gF�(�41���E0
lrk�w���c5k�Y"�#j�( &����	�����R�9P1�9���-�3���sqbC^4�~1B7;�@�ztQ�3�QCR�[��
�π#��N���L�yJpo��1��-��7�ѐKZY��n��)	�ݵ����\g�P�&���fUiQe������Hj�3���P������v�-�N�L�;������戹|�M6'H��ȁW�	;{�Q�E���.�)�>3�RB)������g�F�\�hu�3 �R���HȠ:d�Ⱥ�p:`�m��oȤ#�3G���-؏��y9�F����XC\�I��e~I0����5��c��w�tb҇����z���T�?ѥ�⹰�* ES
I���8�s�/%y���gƯ���Ro�F�[���vI�v�J\r2��u��}^[}����+��"Α���I���#�"��񆂍�ۑ�o�������:+1B��6U�
�=�i�7?��T�)�9��Hؘ����e=������� ZL#��x�c�}4��W6�R�����)��7J�U(,wv��n�y���=m04���w�r�E��ֲ�R�-��J���2<U�=�|��][�ll�$��M$�K3�������q�[F���o��'���m��E��}ݛFc(h����qZ ��j�y-,j���._S��AE�À;]��J�碓.�IZ?�;��|��#�zЉ����G�$FMQ�^~TI��S�3m���FR�Øa�FWS�fW���Dn�ҫ76̆#9�HQ]L�2�i8C��F�*_��hɱ�=a����Ԑ�"���)���*g�sb��ﯭS��rv�qf�Jh3��j��C�M�v7����9˴
H^��E*��g�x��3��H%y�Y	���n�Q�W�V�_��j^�*��Qw�~ȹ-�����yt� $�0TX���@��x�����Y��m�X�J�>�Q\�����pX�1�n[`��|v�D������̓\[i;j'���gt�UG�$v�o�2��qO��sԎ���㱠�Y��@�/��g��%�?�2�eE�����!����pV���d��	8����R5�̷Q`X{4j͇�?���I��id�[L&J;3�5�q	0^����%�Ta'#{�M��� ?�͋�W?�'߼�K8<y
�mf)ت;���l�����}s�(`7h�;�*t��\UU��^~�>tX�$&�����h��o�fl��0d2�k��_e ����9�rm��P�xB^�pI������\z�o%G���@�>}��&�1��tD�,���� I���DL����}E�R6MD��8��/,d�+rw�6�*��U�Ym�LÅ�AY~�a}�\ ��X��`��=rR�A(��+]�
���ۉ�U����l�'X%F����v��A�FO�>���_jZZ��p�r&ߒè�d?�_3�����!�bC-A��ȑc�QV	#�N+xD��-�/싘h��h\���כ;��^cYꙢM!q#����Y}l.�oA`_�J>M:��͞�a����K��MI�S!�������mH�#����.-�PꢮؚuDZv�mu�fDY�㮘ۉ�Y8�D�3����8�R}�p��}�ZM�(N��"�ڥB&��=91�lZ�ȴQ?�=�֕-չ�������W���e��?d�$�Gn�wC,K���]�sW_9Cl`������в �N��pĒ��HĎ�U�9�xU�!��u}_Dgݳm���ˑ�f壋�6Z|ݛoK��#�Y~�H���� �?�ٝ�
�����&�aC \��fZ��y(H�\q��a4��/螝�c�y1Z���5�C����d[�3Pd
���Su�%�G7LH��¹�.���%����I  ���'��y:N��|q��OL�3�"կ��Dՠ����S� �l��]�>J��%���	��*H_+8�x��;y���?j5o@�K��$�34*^ĵ����!��B�7�򡪙j�������ISo�N�S��wg��IWp���tD�
����~�>�G�ul���z��<��_qw�ɭ�i�A����,�q�E��a+22		��E6�˟��8��{�DD��z_��^�(m�3����p!˽|��y���G^�	�vp0E���<���"��bl�$.��P�a�s� �`/;�w�W)RWU���Z��@?�.�r��]���~�n�nqj���f#�׊(.�({���|HG�K�:�U��b�hC�]{�I1�f�2]:�R�@��a쨏�����3%������N��E��ZU���=i z.O�U��	� n[yw�aE<��&J��h!�e�@=���]���9��GgxU�o�y��D�fm�)�����ȫ�!u��ﲀ����p����qN��~G�����Lng�5W�����\��pz6�ު��q�5ZPf+2!�3����oTx�Y��K��FR�*�!j���͎��0�^i�n��@��<�?�K� ��̅�j��qN�����O�(r{�L��ɀ����'�H����~��!��"���[����2ʧ�p&*������sG	�t�sH$M�a��$px�]��W���pt�ssH��W0m��1�C+�$a���]���i����".I��8��}�m���'�%u ��D@]��'�r�JC��Ɍ���@��a�,)��?� K౶��J�UCsߧ�yO���y�bY1����1��<<�,S']�1���k���Q�'��8@���~όJ�\��ҟ v-
����$��ɟb�N���J�Z�<MͱY2r*��y0�]�b����	��rK����Hzg��s�L���*#�\���tD�P^@�D�P���3��7��>�-�@��4��- 4秽�먳�ːPh�fXg��͝�����gT�;�%��-iXCz
Ĥ�à���q���eQk��!��!L�U��R݉��Pep��+IM�V��Cy?Z�;B¢����ZY����j�����$U"�NK�����ը�}\���6���Ǩ�X/�3=��]a��g�S���;	��� ��1�� �\Y�_|B�����P�P�l�J[D�������LM�
Ϲ�=�����8��$Hn��&a�L�D��������*c�S=�r`e 31�8�:n���i6.C.ڲ5�Zs4�7�m�m��>�� ��?�F�Ƭ��ş�:��_�VK���+���˵D�!}�d.�p����D�d�ѫ�w9���/m��w�V����kC}�j��p������?SF3 ��&�@lZ�e�l��!�{�J�I�.S�I���˚ק#�/+N�4���a�i�&v����r��e�b�a�P2ٙ��N;�F0�l[

�&��/1�j����Nb�'h���(�`%l<��i4[����m9XZ��::�Iuh�,�~��^�V�^R�@���j��/w��ލ��g�mt��?�oo�B����y��}V�P������Zs�{��|��	��.��ׅT�a�����B���^l���E���#,���@&j1����k�m�!�n�Xn���m��]���CW�G,oDy���HG?�ͯ���ld��^����X�x�L��F>�A� ��Fr�4�b6�<��1�[���gq����!U���P_���b81�������<}�S��5�C��7S�B�kb��6��`�H��t�%�p�w�q���
%�p���0d�>�v#����P'g:��.�]�ﭵ��k@43���W�GF�#��7����! ��}F���z�<q��[�V���C#�c�1�mg�ۚ���̃�(�_Ȥ�@�7	�/C�@��!�������tU��Q[<C3�hS�D~�\��}�8��5��~�w�o
AM�P�a("����}���v�ՋJ��n�8�o���y�D��}��L���&
y�N�3w>�
)kW��� 3
���'��(�e'�*�$XC��ٗ*3ыja�D-Xc�՜�wc(g�����ʌ
V���=�EwC҄���ke���$�s���KLdM�����]op�_"]�a��L8U�������[H.]L�t����z>���h�[�G ym�И���6D��Q`��5�˂I�w�y��E�U�T�XH1YT�j[t"?���9S�����^���>�W�c�HJ �(���ڳ��,8��C��vq���C��uFܮ�8��#��5QHg��[Ug�lӿL�^��ЂNyy<�	4U�:,y��U�JX'�|m���3]��b��/b�(v�K^���|D���U
���4�T:�?��}wւl��:�H�Fb�ۮ�T#�hWBK	����U*�\��H��Ћ��>�9ͧ�1�H���P���.j�2|7�tjM���7��q/.�e�"?�{�4]���*�4l��~h��yx٣�
��RHU��]���+t}?�"N���N�L�u�8�ͱ9��M#��/g����nΉ�Û
��$Nv�c7�U����>`�G��	��Q^\�橗3��~���J��1Śl��8��j��m���Î��@WKU���%OT�hf-��~�%����(Eb(Pm���=�}y"D�c~@��uʈ�o��`33Ж���Ɵ�iB�T*l�j���O �x2 �{�M������W!�-|\�ǚ�,����% q�d�[���MA,=aB�-�pw#�c85A�I?M*1{�<��r�ђ���e3���xϐr��,��ŋ�yb��;�ʅȟs�2a�	=�h=��^j���(_�4��sg�Ms�R�y�\���uM�F��}q����*�I_��g��Pay��w�1ϼ�剓'`�(ms[�!�w�c>�J�<�D��G�9��@�5	��*�+%������Õ\i��7
֎���{���k���eV�^E�6�#�Xa��`2�$�Y Ew�4:n�aA���u�=��կ���Oo�R����궖.��Ki��`@�W(��ɹ��n��+�����q�6E,��[��B��-J��Wo�%����D �f*(��p�h0�%*��a� �A�7�^�{41~�_�<ԡQs㞶#��k�v��{狲�)w}(y�%ä�+����j�x�w:�t0ڸyܒ�e2у-����A@��q�l��O�:��^��/Ͱ dU�+�>"�T��ŢJZν�+R$��\!WT��r�R&O�(�\R���Ց)VE�^��i��5;VX��/�� GZ�a��$�8�p�=�����]�U#�����P�Фre��1!(��G��
i#~�� �����jWF��α�/�`�����3�ą�	��T,=it���m���j;avk4:R6^�Q�� |�B�[��&����o�X~"K��QGm��u^�b����2�������I�m�2��&����W���%��M��Ʈ�0��#��i��PŌ�$6#�
4�������}�5��AUP�
���4��W��S�3M��VJ^2i�`e։!�L�B@/^@�r�FT�,c}��6T��3����W��dey�g7�!��5�VGw?��2�(�)@dg=^,�A,�V.������X9ݟ����ˀ��-���
�t�2s�P�i8G)e�8���Jh�p�G�Ot����p<�8G��˺�TF��}M�4)�t�yɾ�L5(ނ��e�~μi�U5Ya�C��hD�JW��P< �����附���G�ZLF�_�ɣ�(%��o06k�Ov3����G���|8i'�~�e��]Q�@��ȁo��슦�����1d&�L*�����i�c�S�`���b��� ,+�霚bʊ�"&j��5�I�J�F�{���w����>B�o��q�����;����!j�Қ�"U.J�%�9��]~1�8��Ƞ�1Ѡ�v	��]5�r( ��qr3-o?�3����_<Y/W���侀X�zS�&�����En���J��4�-��8�}89�ødb� �:DyM�d��-��O�zx��_��kC���&붾{,�^��ܠm�Nh\"ł����������0)�)��:q��ɼ���,�����E��.��Ni�7/y�������Ooiii~@��b�9�ë"1!�=��v�~ӳ�C�Q�ְԽ�;���qU��N��0�x_㺗������gHh5/�ر��E��Tgy4���~H�v1<�[#����0����u���EF^��mG����)3b��dq�k>��N���\9/�Q9���E���z틛����������P�7V�dJp�%�&�?Jy	����{�!��5����S?�k��ΊCI�͂i�T9#��e�&7��n}ʯD����8zYv���w��I�`m��cV��lt��l5N�3��ݱ��M!����{�#����`2а	L)vl���Y�:�W%�o�.s�=*E��Ə^�g��=j�G"�ڙ�2B��o}A�G�an��3Zv��O�uM���%k���c��%<S_����}�*�$�N0�ۻEUYp�&>ZM��|�h�쳎L�8��I��v,gpl$'/� �\�}��̏s�_��u�m�s� 4 �lk��'2û��$;�"���1�w�r��wQ�����Ӵ?-!�3T��H��(�Lt�[�*�s%Lj~qA*�e�\�I�7�f�Y[�m�E���sC;���˰-G'}
�mc�o0|N��(��u$H0��ұ0�gy΃\�ź�����O������q��-E]m��͂W��@{CM@C�㣸��]�m(�#li2
���'A��@U��z����A ��+��9��/� `� ���brL(�p&ۃ�ug���'���C}�p`���0'e����F�`��5����U),�9�e��(`��5�	�0K)�7��<S��|1��Ea�w+7���ě&�N���!�1u�K��_�H�\x��-*����ri���ZXл�Ff&��s�Y����^�&;ŧ����
2�,׵	����S��9��(6s�l������Ӭ��c�N�z\����W8���8qT�;��/�+~� ^i-�H��'�W��o�A��`dI��PW�0�و�#�.���9HN$�B�Jta8��A��+�oE��<N��(�w �m�ki�0vrc*Gˈm�.I�3��U?��`B��hT>�a@��9-\����F	�J>�dR�#�������hB����G61o�c�
�cI4�5�]j����z�r��>����� l7E7k�k*��ܗ�4h��ۭzy����&�,�WU����ڔdr0�(�:�����H"06y���}B!��Ŭ�M�-�S��L�24g-���Wf\� ��K|�qy�X�[��k��!p&����/�`EG����ۉ�
�.�{�%[c�W�R�̶e��@��T�4c�9'Z�!,aѨ�ty`�9��\��v���e �������}P�V��E��#�t����P�$��5F<���A�K'@����
����&���E84vf��k0"��uM[\��H���3�2�QDF�������:�ߺ�R��6�,��=���^�]��V��:H>������_��v������D�p��\��BG�t�G_>�rVC��AU�졅{W;�U��C_8��;��[@[$ݏ�����J����� P�����!9V��8�,��J��q}�{�f9�.~j>�/�&�б͊v!�8g'RfX�.}W�d!lG���](�!8�D���=\�/o�V�k8�|�V\� �t�K�Ť!�(ߛU0�Aa���a=Cv������q�c3�"��ק��	���Ҿ�N�v��ENE�b��'��?�){f[�.�;'�O��=���/����������ܜU_d�/~u+�߾����;��NDv'+G!��~V}������9�M=�
�:��1��*_�z�t W�K(Y t�q/�b�� �T�L�C]�B���X�L��E�Π�q�w�Z+!�}�X#Nx�'vs(�����+4\LYB�X��n s��0�2s�X֎QXX��*��J�S��R�}��ͧr���<���y]�*�C/��[�w`�t��¾���53[�ռ�i�n#�
�Z{7����Z����r�Om3^��Ԍ˘{�����^���dN�!b
5�F����J�޷�ݴ�Ŕ֩w>�gجKWn� �2��KI]������Yܣ��s|����$GTp�f[>����5U�I{mڥPn&���,����7l3�9�9���m�؏��#T�a�Q��lU�B��R�'T�}���I|�u���1�ơ˾5:�h�$^�&N�	@��^�-«�vV ����>�S�Ҁ5!�6�8���\�ͨq�����p9�����Tx�N�<}�m>�Us"RaA�4�S����{�)o�O5�@lB����K�\޹O�i+9��W�����
��ɰ/F8��q�F�G$�ܗFn��J( �??/��Ľ��ǐƵޓ�q
��aW%�:&o�|�c���\�T��#�ȣ�﹚>Y���"Y�oC�l�Ǵa���+�n��`
�Im�u�|�3��������"%W~"�IY�a%�?�E�)�e(���VB��P�wC��#��g��P�D�������zm�P�j�����I-�ܴ��x3�|�3��Hn�{�d#@��p
D!�p��FOm�,ra�����5�6���+��jSh�.wהA�H	�A��O�)��7�Z�t�C���'>����C
	1�ƨ�s��uB'��B{kD9��f��١��Z���7���8S|�L�n�`k��j����)�4��ZĎH'���zz��V���B��� ���v~"%v��p0�#^Rկ:�,ў��uu�BFq(l�_�Á	�3�U�:?i��s}ۦ>Ď>6�o�mI��OM5���=�sv+��mi��RKe�^����1�<�ϸEPL<���pe��c��5W��Sb*��Z���r��Ag�]�cj�ޔ�D��C'���Vg�m,�jr�)��bW�\�I�m����b�fK��n�������,�p�&Q��Ki��u�n�/ya�lɎ4\�~��k>t2�b7��$�?+}�-ݝb���PL��%vە��HP���_9ق`s=�K[I.V��|�"��ڔO�q��_^@V����sX�*��76�G�ۛ��G4sm�K�-�B�A�c�βc���Z*r ��X��1�E+x.ܶ���{����������b=0B�PG�<��6��C�L4-���+t�Q������5�^v�M��Be���(?>��B�*�\��m���~�E�kH��c�:������h��� ��H����R��Sы�%9������E�a����.�|a�r�Aw�8L��$�uᖹk�}.���鱎��B��V [��K
U���%����]��*���TK[��g3����n��ў"�|��QAhEh@I�J�w����љ��c�� ��#���Z�:����\4YqU�Nv}�d�0���]���S�K}�k�������E�s�F�[�~iY���gg�(����v���&��P� ��N�.\v�]�1��P�0xG?G�V۫JԞ�6L��Ǆ����ִ�I'�ZAoM^q��n�jg([@�yȃ�ϢgF�!�v��=2Q�P4�`��l��&����8�� ?�X>lX�l�"�a�������	Kܿlq���}E� ��p�frc�h���+����0��߷:s�F�$n���L�O�I���֊sw�+1��_�G���D1\�Z��+B��&-$ᴑ���Y��hц����9����G��aB�JGᤋ�}�FH(��L�
-=L��0��8���Ky_�d'#}�d@��y�Z�i�ٲII�݉��<+��������yT[6�f#��u���r�B�V(p��fp�(�Z�NӦ8��'��8�� �fb K��ǻ�(rIkN����VбCQ��Za�,�1L�o�5��ج��g>�s~)�be��d<�":��Q�_gB�1���7嗤6+��%���Q��F��N��/�I�\$ECZ��G�۹EW���9V}nuѮc�냬���+�wҽ�}��|�&�T)����/��r�M�K� q)���� ]T�o�,�"��g1�=!�Ǆ�}~����w0�^���}b#���̐&>u�o��a11�-�<j��n��ȫ�+��/��KڳB�pݚIWn���惵"c>���'e��F��IIW,rWB�q]�ă��b-��,�����4a�������,�����%l�4�'�.g��D�X�t����~}}�!I�O[#�f%������ԕ^t�n�93OlP����/�<�U�,��頻\`�x�܅�e�c���bm�l%%���Ϻ]��݂j��ck��D�����R�ht%�M�Z6Ij3�(����i��~�ƿV��6>>���8{u��/r���$$������m?��?�o��ll�lBӚ�das ���/��VE;��B1HQ��xD4����'�rhDCE� %�
 �C�d�����<�l	~�Ӗ�=�%�2�c_��lIH��*��n@�\Z���.����Vb>U��ێ�PK�)�%p�ֆ4 H��F���yW� >E�Iʐ.�kxH�kJ�����<xNI;t��6 1��Z�[={~6�r����pB\v��uoW�R,a���|�.f�) \N��Xm���$�Y-���r8�aw-�Dw,��.g��i-�p����&�؎��9�$��t���L��;,�U�G�%�*�x�e3���!/�]��Ud�'�<�gD�D��:ʲ��]���@�1#�Z��r�/�"��	rݜ�h��6��א��R��
*-.�F�0�Tx�W�J[74���!Jd�G]�}
g����?f]���IU���3iE��<*k	W��X{t�t�:GԮ>h�2�J!m5HCj���!�_���� �j��RG�|b�heh����BW#	t����~
+d�N����<d��TDFb��>�ǖ��y����J�n���K�>`^�Q�.n�g,��Sz��N��=�v�@.���M��8W�������OCT�^��ɑLM��F��[�L���>V�qyh��&��<��yy��f@E�J��cS2��慥jrL��W��ٵ�s�@Yti�/�������t�5u(������g��k�C�R:σל���9�&"P��B��[��6���g(D*p��k��i�lB��0⿸�^����v%�1X�jˁ�#���e��O{2Ю�j��Pb��g@.��I�����=�0�Z|�f�Ar��q��.#0�so5�\Y&_�$]���S�ٮ� 䁍>s���j�����~8����TI]V��i#9����{����gA��a���W��0g3�#��t����@�~˴��p��S>��G��PxE�8N�B/�
1�r"y�?H&mmw��5𫝩jZ570��}mk�B`,,v�7T��KA¶��nº!��}�%�RU��u"�J{m�N|`A�*yMPE_�DL��!tu��%/��ӓ�D�8UbCenZ���w	Du��\�FTb����UYr��<���_�_H�R��7��p&�a���/ك�>V2��zr�e�g݆��p؄>�V�<�`��_ٲ����K�>�mN<������7㚤Lb�*:2)������t�S=?�J6�$��E�4 P�e�F�z[3��O{R&m�(�*8��q@�L�Wf�%���p��\���p���������<���œ�V�z9Hd�l�J5\݉���X���Y<3iՆ��,��X~i⯛�R�eK�Ǥ�(K��
�Ws�'�����;�����a5!Ê�4��a��� �����},��k�_,w�O��Y��8:�6Z�[��%� ��5���Q�+�%Uv��D��~�BX��5��^���@t��9�g�S[�֎_+T<��a��ԮX�k�*,�G���6:� �fD�/�褐+{g�Xl��庯���f�S[cg��=��lU���Rh:��I�9c�P4��%^�J=��[���C�oC�����)��ZA8�t7G=:�$6Ҷ��̋���6&T˶����)�J�������i�m�EL3�i[�&Hl/�U�%����B�v_�ֵl-��t){v-��Koz����4�V5�z��dB�����7n>|�OQ�p��ߌ�[Lk�^0�[Q*E�pT+�Z��%Mq\�m_�{D����K��o���3�"��.XOe�)���qK����u�bׂ�\K/z"q�'q���������f|}���ld:��Θ������
 ��v2�yg����ED��.��u�|��1���R��V�VxB����*!R?��B��T�&�	��?�Л���'LY�R�E�~F�ܱ$M�,ve���1.���q�J=FˉE
��O����W���$e��'�k4��kY��i 0b�Ʋ!]�?xO��:�K� e ��K��3�hs��L���wd�K��
��%��8@�p칦,8L-��T8m�` �|��l7Kє �D���x߾��F����,�']dU�Ue�	EPBl�b���+'�EqmbpC����^4��w�8V�� ��K�
���UD��?p$ۭr��[oA��j>���Tٯ�5��4��7a��5�^����5OT�չ �s��J�H��$�U[�E�=e�7���*ڷ��k�P#��i�O�lg���l.m����k�K�M����#��i��qv�A����M��R�9lL�g/�f��{s��� ʥ���f�l�]h���1�dN��n,�[۝+9z�)?R�8B�2ڃ`��$5�������]��F����_��.X!,����pLዺg��z��N���Sܗ�DN5���-�O��^w}��WT����i$��>�I�������n���w¤N~�>��v�^!{]�1��mYW՟��V�\�qxF^�헦K�/��^��BK�D�L*��8/��j��^W�?+@[�������J݉Z���N��A��'ES�i���4 W ���E`������q|���Fm8l̵�}�Ð���C_��o�մʿ��Qv����TS��	!QeV�hz���h��aAE;s�=Uw�wѝk5FLs'*�{���]����6U��/o��:t�rh[(f���1�Sv9b T���]	�0���[�;|�O	ܲz{A'<5p���Ք�ْ6������������"Ec���5�Al�'��r��:\�Vҩ�5tG-����6rP��c���`V:�]���N��:� K�ބ�B���i�����񩬼���G���߇tR��J�G�vA��F^B�DIA��2W�M�jy�\E�xCE�X���=_T%���Ի}Ɲ혐��c���F~]U��dS���y�����z�,_�T��?�k��h��et�+3R �߅b� �E���Ch����0�(���K,��ƚ�����W�խJ�A�H�W�- �!,l#��>�s�ŉ�O���R���u�aJly|�\xlr5xU/�;�S��H�$���	Mp�X��\�5d��P;D:j#෵M��R"}����	&��-��B��m�+�*
���@VB��W�� ��"6hH�w�	�I9��3�1��Fچ4����e�Lc��jQJ'j�L��C73U�$��Y^Ѻ��	�h,�^�*�h��?1�/ie����I.KJ�ċ�$��I޳��R6?�5u;OETW���?�8���Q�\��ڙn�z�8�j�~*0G{�v=&V�O��=��w�P�5�6ˡ�{�.9)�eR1(�������C���(ho����Wz���l���b�m~�o� �WOt�O����
1c�������k����L҄Ч�c2�:SS�	��Z"����]��]1����!��d�d��`���
��J������i{�H�v�m��IffJ�h(z��L����IS�gw�-G7Z�k��LT]� �&���dS��-ܽ�)"�
3��+��@��D+T�;.QO��yj
è)h�%���2�n�Q!T&�k��KzŝzɗN�q�>�ѳ����xЃ.6H�X?2Ȕ���?�-p׹�Ą�B�807�sly�T�%[�q8犐G���[��m#�׍`���Ÿ�2�dyҥ9	��ś:j�?��d!��y�b�T:_qH��]Gq#�����=�>%B����2�'O'Ķz��xݐ���$���b��֒�����&�i��Z�,�Oݒ�����z���{��d��3r[KaQ,�|r��0"Tn2�t�EV�Q�}^��v�K�Y�c����w`D!v�U��&Ӛ�x���"&l��Z��c�ߐ���0�k{�^	Ԗ���b�jz%&VV�X鬦}�+��3.A��e?�s��6�L5a��Y�%v�0M/Q�oa���e�dL��tz��(g�O�0[��a!�4�|)H��-˪G��Ą�������%�"�^�V��0�Aۭ:� ]��N���B=�u6 ��`0�vR����F�
rԞ�K�!R��[y7�-Ll_��# ��3�+=���F,Si-��ǲ<�cfreC����U�A�d|�O�y���/~�F=�y��̂�k� �ul\�iu�*��(�Pw�<o�0[R�����!�]�w?H����VI�W�ѹ��Ş+] �P�Sk���f���/�� 9ӻ�_�1������o�5~g�Q4sRc?X^��.R ��3|�神�.ʹp�g;�g����pS\-�vr���E��wB�<�M��dwT��=};$�ȱM�XJ�L�}��E���s�d~�_�D��A��ެW��^���m�ȃ̡0��Rm���n�n��0�"����o�}Ɩ2kt��6;�1���<��d�d>��sK�N1J��y ��.$`4�,����2f�1-�YEW5�.�)����/X��,@1<��XwU�lc�N	�"'�=��OI��4G��)�a��xxq�������� � � �́7�����7�`�N���l�A�È��,��Ũ2�c�:��*�|H�2 �4�W�"u"",�������>4� �"�8����-o� P�~F�h����r����;���p��D0B'��W~`����qQ]V�7���}�BC�L5_�!o�D%�X�I����h��}�Fy��-+�}��z��	�-[����P��x�M��A}hmc���a6 ��Ƹ��6��⥤������V���uO��Z�y'mK!l8a��ę�
,0��$�G=��P_�a;�q��d����vˊ�3�&��\���M8��>�1E����H�N|�4Q=��
��؋F�N��"3T���2eue��~('�	����	D���	F�%fʹ��{`�3�]����4�=u�)=���D�+1�#��e*��t��|��'��K�;RJ	��*�\������"=^�T�� �{=|����Κ�d3�X�b�*$��Ŋ��T�6��崥k+G$�ħe�أ�AOvI���k{�oq�E�垦����A���|[��ѹO0,`�����ߏ����4�&a�/���5%���_E��Na:"i6;�%��lF������_�[7��x�0(�-z�HW���;�v�Bf�ec�6d�d[����ƞ��ʣR���$4:vAf�_)��[��{JM��
rT��{,��nt���=^��Z�<}n2cR���M>A΂
�=���d�����$h�`k@$��{gy��V3 ^���"�gpK/�VVͥ��!ʽ|�9��$�f��{"{qZ4L�O~���ˬ�5�Z�����>���ܠ[���E�q͔��K`�u���ĎY�;�	�j�T�]���H�^ZV����������<��J����{Z��y�0��:��L$�n�PƯy��E�d���f�#���jޯ\j����A�H��AA<@vdC<��uY�2?��ǴTX�t?��<y�Z*�,/��6�~��<���H&��b����C�Lh�Y,C���u�u�|��Q�h%�*�;���~q-��MǱ�as.���>��n��3D@=_P�Y
�h�{��2��SPuR�����?D���=����b}�z�f�]�M��o]Y��]�lp]��Hs�os�:��L '��?�v���J�+�'ܟ8#u�T�ߪiv���&�e���8s7�'��~�݇���Y'�oI�;�z=�N@)`k�x�����Q�,3�^��M\�)�	�iO���Q��2ÈTEUA�~����f��f^ٰZU
�b�ګ��&1���v<��?�!�d�b���Y�=���:B���9'�J��?`�@����pߦ1@���n�2`��������H���~tW�7�CL�x�M�I�*�{��]XbT�ܻf�����GN�*o�y��D�>���n������$˸e���퓢��8�k�'��`N�+�u��]#��A~�]�e^/.���j����L? ����,��3�W5�tVn�;IR����9&�*3�q�}�)ϵ��6^�KM�:��IJ(��j�X`�����=\���@�k�2}~�O�:��9l�@lK��������V�&(��#�rA^%Xmu�^9YXG�%;?�� �W��1
�_��W��Kj��T���vtč����hL��=�7�/�G���#?@�č�<��]�����@��L49*k>�a��Ղ��1�tJ�'�6l�ǳ�=��0�6 _��v�!v��=h��}�.����D���	G^�k�����F[E��|ޣ�]"�LރOV>Ϲ
L=��� r�&謌z��)�U�ۡ��w��[�!���'�+��gn3�)���� 0��ځ���B#�̭��M�l�ҍ�Pqg��̃ωN��G
npF�v�oݻR��
9����|�M�3zFӵ�B>�h�o5�l��U@?vo�^��`$�+�Z���l�N���zUX�.�����zV
�{�n�_9��n� ���m	�dn̺�����5����M{��{�ߟkR.[���N����\�./Y~�PȾ}�~����1"Q&�SI'sޔD��Rן@�:���͂R�5��z3Y�J�s��6��?ɴ�mX��P��/�σ��&"�6^���������R���l��Gv.b@�׊�1��x"(1�fHu��S�d���I�q%'�\B[D�-��#��S������Np��1y'�z�ٖ�A ��@P/R�����j���Qڨ�v,4[˲*P0�+J~w߾L��YC�5��u�|3�D  ��c���A&����2y���p�1EG�1*cD�z��\����	�T<�������5���~NX������++݂3�����B��ؽ9ͼ�3�v�1���ی+���*J�h{�cF��gs����Rf�(���d�i�<J��D�� +%;Z0��x��7��N�[�i�_\Ȗ<i�T�z�AQI1�n��7�*P 9���*��Ġ�.�v�H��m��1�w��.���M�*�hЮW�д�� ,�g�ቦ%	�?�l��:X����jk�n:U+���&�3aMp��U[\�N��~��f�xΡ_ԍ������Y.��C'Mp�������H���E���j<$�*-�,��k�5d&�ɕ�R��%*f'TjNC)i� �E�X^�Hʒ�]V�|J��/U�'n���ఱ=6�n\w.�H;���YD���Ď�qd���7�(��9D�n�Qr��P0�4��QYu��F�1�땡�ͥ��
��s)g\8׬����'+D�c������z^���=��B��0}����3A�#��3�6�eג����3�|�g��E�fu$��B�z�(8a+�d�J�
�*���ҹ�F��#�0]���`�e'�L��T��H���f�K��Xɪk;�(�E:2L��5ˇ����v,
�i�H��y9��~ �{8'{8Wn�T:��j�!l�̀薅�">l8�J��Z�<V)�S�������n5��5�#����s��gؑ%��'��i���6�G��]ce+��:rN������[���T�^���;X 4}���\�J��8.��&�ͼR�^O�R���Eg���p��]�&4߬%��F��w�d���(�.��!A����B~��#�G�����'^��h})y� ���HPq4<�J)�ZEU�j����Y���FL��9�N1��K/�j��POҰx�^�׷�96�@�B�pGI6�̡���Oϱ����ܙ���k�	�7/�ץ��]� ��;�X��]x�����zDԯ�s�-V�)�['z۟�|]��FQ���2�X�y�������*�%��fa~���ݴ�3j9*�ґ���vW���.<g-V���iu$��;�H�_g�s�ɚz��"ش��N�aF�T����U���*���6�y�R�f���i|��G�7��X�`<��M>c�����7c�ձ�W�;R���~q+���q��/���X�
[w[��������l��<ڑׇua��������64F;z����#��;�i��P��G`f�d�k��t��@m���vo]���٘<�in�`�\�l�3�=:ƹ�Ys(�`���]@0�|�G���nњҹ���ϐ���O� ߲��tf=R)�^�˪7�vB��x*�]B�/p8M-?l4;@��+���D�Z:��J�����U?F�Re����~�cP20OW�8�|��׶���Q���Z�h�Mv3syl�KS��j�A�-��(­�yj�V���>D��;K�;L�K�T�x�W���B�B�X����03����&>/o��`-��_(�3]ɸ������A���k����CV��a}�$TP�K�_X	-�-5�t����[6BR}«�f�[rs� ����!j�{�d��Gc�1��:���E㔊��K2�L���5�4#\��@�O|UIi��n���-ᒀ�Da;"`R|�
QD��������ZZLf>�P��}��2)'��M/z8�����갎@��;@m��l*!G��[+���?�6��2�Q���h�9O�ܺ����'����;��Ŗ�J��̧p����� c��7��L����h*Ɣ�:�cp����oN.��m��ge���'���Î�nH(y�����*��7"�0<�gǻ�E��P�5��I% ��7E�3XLd�J���Y%�'S&Q��\�
�Q��!?���t�!]��o���8�U�L�(�͊1�Q  �&=���@d���|���GV���c�n�B�-u�[U{j�މ��z�Z�`5qD�;'2�����B��v��fXN�X��Y�L���:�z�*��:J2pSu�1hC���E����.l����Stl>��^�f}���ܺ�D&Hy�f�m���y�lv7���Y�
P-����/�2���wh3��H4;�a�k��J�ۋOH��Ǿ��V�#]=�Փ�U�,R&f�h7N�w�t��K�6�!P��5X����e_S����n0¢X��q���T�zy��{��-�Q���7�����c�w&p���/���w�?�Ɋ@�7P|��ϚmI I&78D�F�ͱ	��� �,�2�]D�]�PN�c�	 Y�l��% z��<����s��e����݋_�SSc�\e��C]�0��]lf6�C��17�D�MM8iK�@�D���,�9�y<�;�)�SB�PET4�~���9��i�.P�>��Q�����T]�U�@��l��r�ciP��&�g��w��]����Jز
W5a#"��Ԑ��=��8s���*ӯ��d_q抭S�b�	@��[�:QQMH��hC6��g-�� ��	���K��ՅK�^<S�x���5����`^(σQ��X��w�����A ,H�8f�h��#O��˯� K����Q"����qa��Sx�#��܊\OPX�7�+��p_�,+>3���Ǖ���⣤w�P�2�8�uj�����i~�KAi+�uZLM����f�C���Θj���ɏf��x)���B�G����_�|i(g[n���-��hJ(���=
.�o��׷/.`��?Ӳ���z���>�ʝ�i�ţ/�Q)��G�@�`,�����x�ip���D�s46�;����F��Ip�Ǩ=u��O���\?�����$�/�:�����LL���Q͟ÿ���L @���:��ugi�����4b��3�>�$���v�^6 �/6!�;���,��r��ς#��[��J!b�r	x���׮_5�{�G��)�zA��l�t��D�),խC�z\�&�1�6O*D�����{�u��>����`�wA�t�זmK�6G���3�m(C`�	��h���HX�*J(_ո���^�{5oZ���҈E��g���˰�2�
f��1�7�\�%t�M�
�,�O�츻b}��Kg��ᇋEMh�@�Ӝ\&�;�5b���Dѧߵ톚N�f���ܛ����0	fH��bbƤZ�������b��!���}�����/�W���4{5a6*/%��*tNv1��)1��!d��ċB�]���kϨ�<�h`�k"UD;���a���mT�c�c9����oD5k��i�1c'jJ��0CeN��M�@�s���R�3m��?O�i��[�?� �c����ʶ<��e<SX��Lc��'�U;� �٣{F}��	EE�#̽F�/^d�o����	��^�N�hCq[r?]]'����c��Ʈ�Y��r�O�f�0Ra|�%`�`�6��wN�8(���D �zz�֘�v0qe��wҘ�wΫ�����L��G����`*�C����IF	K!|�A#.	9�P8�2λP5�wn��"P;$m	��(��Xs����o�9^߆���=��>����y����Ӄ ���f�"{4Yȧ��C�>�����k�#D'�ŊҼ#N���w1h/��$3g+��&'qV���A"�¼$"¿�W~�.k���t�B�L���Y��f_9�?�O���},��"��sXvݔ�b�(�����{��
�9�RU�h��oZ���W8ť2���:�˯V�
t���;hF�LK���=7�H�<�xO�_�>Oހc"Ŗ�?���M��B@�|�/�2$ڳ}/����C.��q$�����kĹ��_�z�-eS��YI9kʪ����?�Y�
6�N���0�إcc�WF6߀YE(Z���<�㰾zt�����8��m�WP��/Wx#�IL�x��j�y�u��nT�;N�|`��q�6��'�c�3�R�o��fp̦�b���p��]��������F0@cu���_
᥹^Y��`��~��>�?���*-0+�i�.q������$5ځ�b�uuF�����PImv�Y�3��v����Z��̋3����b��B��J}vW��d�o$�*!�o�����Ѹ�׼�aQD�0�=̏�H�� ^_�WRI�yk ˺ø��<*RΫ3:�uǿA� ��J�A\I
㝧bKo�q����d�+�/W?t�wR��L�/�R���Y�ʰ!i�5k~�r�q����7�.�]\�a���Ru5�$ş�1�)��fM��?|��I)=�Ef�VӳѤ�/��(��=on �3�HmtF�V��	��ѓ;9�||\��Ջ��i���e��0��]�-r9n���ҫY�q�B�%bZ��v�T��������Z�^
e1}�X�?�����`ʷ�E����=)��l~E�g)��z!��,�\���6�,��A,_�3�֒~�o�*�{�Kw�c�?���3B��Jܓ�Z�N? �L��Ȓ�{ʋn4[�M|�$�.�09'F��Ub����FpO���U@��}����1 �u��d��{]�4���HU ���YbJ�ŝ6�/zfw�\�R^�PBJ�Z�9�8R�M����7?��SW#|���e�g�3�Km�9<�C��w3�����o�9�o�����McK�D̳���s��=6���y����c٠.��L�O�b��cw�A�ȺF�ʫ���qqx����@v4���C������j��:���,��g��fz�*X��O�A��!��!�"N��o�ЅW{5'7�ˁdJ��K쏊�Eo7's(�6�Hk/���~�6����%�:oN���a-�;����^c��79�9�O��((_�7h�����z�%�Z��,*�F��o̲_�h���<EF�
{e�h�Z�ь��a�h��7�g�r����z��J��`�rL�«��R>�d��JQ�uu���7���6����Ϸ��ώ��fk�p��Vʉ��RU��Ci�3�~��f��;#��E&�|�����T!�c��9����l|}Fw�K���=��I,P����}^dԟ��D)%��UR�ʭ�QA���=�2j[�sY\��	cʭ#�MSoT�����C�̞�\Qӏ�I<Ă6ƻD��t�o�g^�C�?k�3�ݾ��m��v$�v#Mf��|�{x��2���CP�I &nGd*!nQ�eӡ�J�Q����GN�ծ�V�o^H���k��������3�:BN�~(�,� ���(��P�/"wa�H��$��f��	b�;ޕ�p�(��Y ���lbK6M^�8J���Vt����F�b�JM�+'˗�"M��;����9����"\(�ɜ'���vVZ�>Z\����H����(�N5{bǢ��f��.�uY���� J����a����-'�Ku¿wb�sF��d�9�ܤ��-j�܆��y���-C��㼐���Y����=����1�?��,]l���Y��6�:͉�cP���i&�fz�`�P(��/Zį|!��w��V�Q�c�&���uw-t���51+2��M
sٗ{U�,gS��D@�j��^X�m9�>"fw�\l1Bp�*���  {�h:����R{r����F;�� ,7TrG�^�������m)�\ug״7��ǣ��-�ĥT���E�CW�^�pWec+~v��������,��j+�xw���9���ب-7�����(�}cKh�ٙ����b�|��	Dݒ���[�͠��v�,��>o!&}t��a�N�k t&��+�U�35pA'`��}������y��	��-��.�%Qk(-9ע6���&�c�A,��كn���c��9'SΠ ����iI�ޞ�<���J�&֗��ElR���*z�8XXb;�R�����Ba�s+��ާ���֙!�x��aH�`�£����:K���b�m �N\6�%I�5v�@N|����0�LE}��#�w�2ӆ��4��i�@�hw�=���S3wi���|�)|�v�ҟ���9�/�9[���"��*�"��������h�Y�ϠCФ��'�C@����ّ-�*�	�[f�6ҩyR��@t��\ѽAK_��Y��و�DUS3�AG��Ue�[q�/��4붪Cl��ʌQ|�c�qB����	K.�o���s��{�|)� 9X�j�K�*���X��0
�y�ԃ��-^������Ө��+�2�'x<-�OM�u�7� �8�g��a�Yc��׆���g�6��Qƀ;�+�ۍ�BM���X�|s��/���1ppȥ�+w������T���E㮶��u��e�$��?�'�m������)l�#��F�{��}�$% �R/���k��}@�$� �ʀ���#*i'f���7��?G{w���b��ő{�)�-��d�Uv�G9, U��]g9�m�h�\�V`�K]��r�h��x�HIC� ��}�圙i���ho	�SdB����o�69�5_2
�&�ǤB}�s~�@�ѩ�̾�� ���zi�@�lb&�mpe�hB����FO�u�_�\���x��k�B�-V͇\�\x= �i�s�/m�>��u��dC�L�o�kf���GE�����z��j+d�0���~���7�y`��WV�v�>ݚ7	�@6;��;� ux(���M�����*_��g6��"��"�	
�k����c���ƻOz���򹄇�z�^׈�{�60�B8�Β��K^_�`��VR[��P�@=bP=��!o9f�m#��_���ؔBwT�
���rv�q l��$�y�\�౲ˊ�Pd�4&�<���Ѣu��Չ.zuQ�`�E&+:?(�Sd��W�9�CH.�A	43��_4t�s�NU�k��1nyY:9�L&k�9�c�� t�I0�3�>!K�L��6?>��w����hZ����hY�a@�{0�әڪ��s$�`��z�M6�~��ҸM
��&�;a��]��3�����F�٨����3E"D�.�g�r�v�ʂR_��H '�y�Y�� ��9=84g6����Y2N�O�
O�F���	�3R-�G��><���T+D��U��ֳ9?���2m*�_���yA��@E���Fm+�k�>����ek�fm={��>)	*�� �)uՆI1"��u�t��@�B��KD�jy�V�f����)6ӗw��UB�0��Kc�6�M�:otѨ�Խ0Q��t:�;��ci�Bhb�E�9N%"-�J��;�:��J��ge��gG������7�b�Zp鰚��mz�$&&�1}�"�y��˃�?y.��W�M~0kU[�U�t�{��6P��}�g4mؾ�|�J*��!;���֢�C
/���vo�F�2��ć�e�����v���<<(p^�����2`�#={�\b��'�Q�v�@;�%�c���6�j�Y�L�O.��8�^�@�
Z�
��!f�[X��-��F����t�����L�&k=hc� O-;�������Y����G]	�Dwi@��[eJdtY'	2R��C����.vL�`���pO�_=��4��\�w��\&R�(��}z��}[ 乃��)~H�2û&�6���D��}
�T��A����0�[J�kOvN!*�H�E�ɾ|�C�_�8�8��j�a�a��HR�>�+]�f,r���xn�}�cy����u����/�w��&�^�W�R{t���F-��
=�w�û����\_�*�>g2�a��/�O����4��/ن'�P�|�����gm|2�U��F�h.G$�ʻT�Fw�NAi�l�� �j�c �I�M��!7�*I ē��c��ǒ![D����(xY�7��Y���$�l5ɟ����
n$U2?
]]�&q�]}��eǹ��v�h=`U�z@7dz,��-��t"DeN�T�U�+�f���I^� �pR��H�ޕ�{эRɮ9���;К8�""�7~��97o�Vˡ[#��c��:ך��s�����f=C��
4Zr�$3f�=1LY���1��h>�B,�"�γ���sf��ӊ-x���)���0�?w)W�`e/�X�q�n�J�͒Pj�	ޚZ��ڊ�;t��s6����1n�aSL�>�I�d6|����3j[��yewMD�XQ���̢����kÖ�?#`�0!홬�EFɠ}b P%��O�M�d����؄��6�I��5�4v6th�˒DM����G�����4�(��# �٧��s�qY�:!�BM7Xl�.b��p|t�L�`���#��6�����e��o����e��H�jP�5Q�9�����}�>�4zA9���R%A"\6<ڧ�&evn%��O��s�8 k�,K:�ˢM�ϴ�¹�uz��*N^p��OURT2�л�價z�4T�7t�+2<ȣ���wn��ԑU$��(:�<[-֜q���#_۟W�Q���>7�b؎!'�	�P���b��48(?8�*��-ߔ4���ʯS5!>ځ�z�Z�d�	�
.�<�	�*Y����~�_�ϒŎ49ǚ����|���!�򛍎��%Nm��ν=#�mھ��uȑ��.]y���7��y��������:����F!��$^��]�Qj|<�E��jK��f^m����ă���e��S�kW`,"�u5���E�򗥖�R'o�J�Ǒb,�u�6���̀
�{�ŝu<����煁;��
0��_�1kE���U�?ִ��& �֧��. D���w�����}���,�ui��=���aBM�K�zĞ!��d���t��̇UP��<Zv5nD�-��{��oчT���1��m^���������?�1W���T}s�)��T��[���/U�v};g�RԿ&�G�j��0 �[<�Cژ
�ȉQ�Ex�������O�����Sҕ��~��6Q��ّ�[=��*���	QD�W��ys���!����*�2��."H@ �4�X.}4��^S��E�~9���.\�TA}�6FXm3�3/f�uD���b�B�Ho���o/n��w��6g� �*z�]��)^<�my��,�&l�?>��Z�j�u�'u��|�4A�x�W]��6����Wa��W�"8
nFl�(�DrF��8��\:<���q�<=diy����s�Dtʁg������8�	|Rl����R���}� � �Ot�M��Ԯ��υ��d~4�	6e�;tq�yGۯJ�-eg�"G}YO�ފ��q�L>|����Lr�dC����W�O�4����jO�7�ȑ2������ۥS���(�-4���,.gh�TQ43w}G�+K��<3
��m�#QF�A�QGż��
��3����n��+i��	�����B#EƊ�r�#�E(���P�F�Ʀ��=�Ԩ���� �c���(�����@c�r1�im�#@R&Φ�1�3/ׄpF<�A(�e,Y<o����#�q�d(�D��9�W���J�[�6R�<��S8��A%Þ�T���i\�<z��?���F'~8 ��3Xe/��7�#l.v��b��	~�c�Z�|!�9�YL�?jN�%���U�ɶ�T\��\aS(��?���>��2����kQ3ݥvX�ÝE��K:҃���6�1r��Lo|XU����0��:	�y�ᾩ��2L��QC���K^K�(F��	V�J��Go���D�@e���i���r�i eK�~+d����c�B�F1zc��:��,�Q��)��݇6Š���a����%[k]��Ҟ-�PKYM�r�<I9֟������L���h�Bo������a��uΎl@���]Oa����B{��j��ֳ"0,��
K����x�����=�"AG��� q(�A�$��Α������hu&�@k��u�y��D.���?��4����eu�A�aϢ>��j[���ϸZ^-�d�� N�|{<�bJ�����<�=�WVɹv�)�-f+A奒i�qҧV�Y f��|��G��Y�V�8� ѝ�D�+���!/���:��_���}#���9`�!Q�2ÿA���ڲ���S>s}o(Th���M�����p����UGr�!�\aW�����8�ǬrÎ˧`��`�. ����; �\�^J����e�gU{@Tn^�5� �Z�t:�+lέ�81�T@���ȭFi�3���*_li���m�ʠR�j
�Q��ZB:EiM�R����Cek^�.p#���XP�<9 ��D;������e<����2�ŧ�����d��p�(
N��@ �'��g=������g7��R�hz�)�c�� ���n����=�u#H��	�\;���~j�z���S��D��]Gȵ�P0)� �~�;|-�(��t�^���>��=��/#����7LK�yD��ih�-�~W� k[�*�\A����J�W����
�	F�� �!�$[V��m�?y`x��־��"���D�GS|��
�����,���U�Ȓ�z� ���e�*��m�F��MY����b�Eu+��q�Q|%z�t����T�A�����ؾ��O���F$�4��K��aI�,�k�!\V����)���ø��X���S\�^��;0�E�������N{�M}V��:]��|&=�=��?�u����}�,v�����d�Z���x�mb�
��	(�J�&N?F�xa����f�h��!���RB^��ɠ}9��1���jl����E�R����d�AM<\����n7�H�<��T��Gj5I�(�濯����L]?��Z4胗 ���CI�D�iO�7�-FE��O�c�@�mC��h����1�	:h◾b���΅S>��݇�*ڿK�oʐ/9lI�,đ�	�h+ i�)��rZ��q2�{�[H:�	�K�JxY��zϦ�d�R�x��~��8�������1A��i#"��s8bD�ZEY\<�W"i�?�Ou�A1��Z�+�Ud
��$��UKl���,�*�������\?��XJxԾ�(Y�I���}ìN�?=�dg���������~S��Զ�Hb8���ɥ��6\1�~p���)ݏ1��iOڥ,��i��6鬶��'"aɻ&��i�!c�tj����-�|s+���3�Ԧ%���a֥n}`
E�]�;��s��/5;"'%��RaUDLh�C���3m��#��@u@e(�RO�OM"��?�pL��B�+���Y�i{~Oˈ@w�-�+��'�]�>��!�Qbil)�%��]��KQ�w��~�ON���_{��DG2���_�'(��6V���b*��A�W7	ag��z��׮���"�����qcB�e��d蠑u�V�_,}2�[�y �-�)*�I�eGN�ĆF4~2�S���%WF[�l��F|g:�p��~�;
#i�8J@�h̘g�D�֍�5� ww��T�⢕�\~�q�i��j���V-��CO��e�"�u9��\��x� �0M�����L�c��?8O1.(NT��9q�%��\ M��	��uK.2ebŦG�tؤ3lW�f��������ܻ��VZ��]�����oU�Rj{���H����g߰�f =))fW�˰��"����Ӕ𜄐[OG���� ����"�/���My����;���f�Vk~ː�g��Ք��	=Q��'ˣу�vR�g��|!!6[�ݰn���b'�۸B�d6�e������NSFi���Ҟ�O`�'l���=��~�)ղ^3m]���i�<5eBG��(�i5�X�$���,���
.2a0le
��[
��t��K>�k3���]�7�V�E�E�$���2L�$ǛC�'��?b5�cYz� �R0A�B����_�T�`�</��6V��<�AԬu�4���}����.�-��kQ�"�j�}:��[�5ax�o�;�&g~��^r�pJ˾N�fj	����Qr�� �+3oQ��v�)t$' ��<$C�H1�u
��5C��Ĉ�?�	<�j5Q�ay
 �"�9W����+��3Xٲ��ׂm%�	2n=��O9״���G�Р~+m�z;�u��κ��5�sq4�O{���I�� 0:�xH��R����W�e��`K,��'�K�t ����Ζ�!�������~��
�9�LS���,<�C�;�B6� b�CŖ��t )��&2|]Q�pUT)��S(��B?�XWv�@���b�:0��qz���ax)0-j��0��� 
9S<N�qJi`���@��-;���S���$r�^wK��H�[����`�����Z�����H����-~�U�N��:�	T��&]#��;y�	�>t�BZ���I��,��d`&��[E�+i�O�ݴ�XuX/C����;n���nۭ�l��`��)*��m�B�g�5����~�v�7t��@�U��;^��p�� �dċ�j?�W���o��D�k�0cz6��$F�����N�y�/�4���)���v�CC3�AZmK.e����3�Q1���]@X�H���Er�`8�i'7��l\Gl\��q���%��,�)��V�~�|?���\0�uq�V�=RT+�h_X��˲�k��x�_ѝ9q���4��y�N�z�As*����(F��
Ø)���7ξ9V���!��O�r�	Tg�ev0�w�Pێ�ѿ O򍄳ѐ�B;̳�f�,���y�PNn���CtE�YLU�bNд'8E�z��z2޸�稑.�r��a&J�;Q�~�q�� S�2
�۫U��]$L.�h�pٗ�2��ց�}�Ն�ό�R�|���v
����8;��P,��MI󱢃��c����.��/i��jR���45�D�8���q�C�����m൚b�mE�~�;2}�����%� ��W�Dh��G�"�~�d��jCc\ʐ�٣�Ьo���D�c�����ttRd���Bz\�_iI$],[F�V�$��q�Q 
!?4LY5G�d�������	򙭔L-��u���~���1�t�!�������%�jbJKc�Xn�9�x	nwwq���U���?���4�|�� �o	�\�|ljj�|�s�����[g�}���h�u=��3������k��!y�2���)���K�^���`�܍J���q~�I���N�R��7��4��zS���䠞H�w��JZ�g���m�07AE�<~�p1_���� ,E"J����%�O\�>ނ�S7��|}�j���Ȓ�<���$kR���*	�Lm(�Z6[kt��<��1Z�����b)bNw��ش"��A:\�Ѐ��[0��� ��w3Q��y8�9���H.�f\�#D���.(������%���z:d�Ǟ�_��XDU�2Fқ������Vȋ�;���~fn�h�����t�꤅���2��t"W��6�=׸\��S�O:�Ύ��O��e��j��i�����$�w���̡�@�*�0{0����-%���ǲ�^�qi+�Q���[nU���+���m�f���� �,�(�n����
�N!��td��Ԧrͼ��jU��b�$`�0�3Lښ�Yظmq7v��90��F��l�myBko�f�����WlJ�����wb�XQ`{!���	����_��o6F@ʷ]^n�U6�13)�x	D����֑ �H'�2�BÙ�R�oQ�~ǝ���栢g+�}'���ō>c#Y9���Oh g�������S�f+�zC>����f��6�q��BL_I���8�#םV��)#|Zm2ZtB,��\��Ƅ�;20X5�I��Z�#6�@��[��^Wpj�v�n������J噹�,f�m'�N���ݹ�
�o	���j�c~�_&(j <�y�ڦjU �ˢ�8y�F���Lf�.s���ͻ��R�e�gts^B
�X��11��cB�{��+��g�r*u�t(Ή���b6k{��߀zvT�b[
>���1h�9%F��'�E����V�����P�r���ND8zk�ɦ��T����c�^���f�O����^��v/�	EW�5�/ܲ�*�~�)�8�`�R+w���e���EN���7�uI[���W�b;�Z�Y��#VbP���!Ĩѡ³q8η#��GI|�����|� @7re�,��#�=\UxW1l��{�++#Z3u �YD������ ��L�]3d]�������fhʀ�����q�T�=���FJZS�<aP�y!�Q�kp.�ǚ�WS��|�{n��ctv�K 9j80}n�n�`��9,��c*��6�����Ox��h
!��S+r�R�4�j��5�xv���/U����id� �!lp��z��]A��͵�>�6�vY���	���!_e|����<$�؇�2%;�{��5-��C�ò�oсN��L�^�U��ث�BQ�6w�T����q��9�V�R�������1t��,¬���[_+�\u���  3(��:��RpHQ�A�k�>���N�W�1n�l��X��y9~3;}~/w�~l�+:��G�|Ɛ�yf��U�Ql��ݔ �`�ONި���ރ�/�S,=Й�H?Nr��R5��;S����$����� �lZ��榠�����}Z��!�p96��ގ'�9���h�(̡����9щ���B�g�h���ScO��ƐfZ��L�]�O���O������3�Ou�ۍ�\�d:rUnux��S��~k;1�y�E1 L�T���7���@ٻ�t�7	��xD�����[���­�u���̪�[�YX����5_ȅ���Ƒ�U���$���o�>):�8�r]TG.9~	�=2�? �3�ޤ���P��:�ݠ|c�Et.HE��橦6�`��ԍ�����=@'��3�21��Q�Vu�}|raSY�����X_tdB@lx�E�a��I��fsb����'	���� �Ŏ{D_9by��f�m^�{g� x:��=U0D���w�*3�S�J+���eェ$-�[���[����sN��jNBGg���0��qk���]S Mޜ��KQ��X���C@{MS�Tʅ��XADקs�^h�'摡��2�V���Ԣɟ���r���,�̶�B�u��f���tL��#�3Il����n�a�cC���J���:�M�CB�5�F��N}Ic�u�-�P�-���� U��@���ΖY�&p���b���BNis�6�T����W�g�.G�9d�2��':�:(�1u^O<'�i�)�o�5J�w����M`9g�DV�L&�̫�e��J
ᑫ���l�,�-�9�V @:���x�Aߣ���r|�tyĽ�6$�(a���䲀*7������T��2	h�;�<e4���S�J�=�乇�G�
Y��Β)h5�k�@l>Z-���GS>T�;(E�aD���������O�Ǳdfhj�*��?ߥU5�Inl�]�;~������=Y|5+&gI2�;V�_���PQ�@��E��6���g3��1�;|�h�=fK�U��Ή��C����o/0��\7zH��a/6=��p3i�'9����*�>}��S�,���Vr�e�Z�<;K?�〠)D&AY) ���2즶b�t�:-���
�U�,~�\��f׌fö�{l�t�7X`�A�q�.(�{�($mi;
%��ü�)E()�c1�W�Cn>ƒ�V�{�59�ï%k�ѣR�� +I�ґ�bM`�g-w�=��S#vũ~P���{ftj�**�Y�A$T+����� 2�
$�;���0�<? �ZS�o�&4dz���y�q (���*�m¨ ���ر�3m�!2�j�&�P��SH�aJ�fof��T#
�)� 9��쀘�N�\�<��E�1���}��ٶ?%�znt0�5R����E���`�l�\3#NU0�O�]��1̀��В�I7���@Mc�b�4k�w�����/ŕ�c�k�� �afP04�8�7߁�������;`��@�y������A��Y�Zrvu����j� �4��wr�	��!�7��60�9�.}J��D���rW��o%P����	�����!�l�d��h{3g�q�/����3�*�݁;φKY[��=������(8�˞��xI�z9��i��b����\�v�A�&y5c�k��xY�G����@�b���h�� ��bF�v��WpgJ&�����x�	�m���?v�k��@,/	�A��I��0�g?TŢ�Ԍ�(�q)��غ���o�9_CO$�V��ӡ�<��ߚ4���xeqT@,Dj���f)i���Co˱�PA2E��e�D�ӓNc'���P�=���Sm�#�D �{^��i�_�#�P2�����>&��EN�:������E���B���㻦9���H�j���eD�q$D,��( �HQWI­ �KJ���V�S-�����*�$b�t@�S|b��>R���G�/���g��a����q$��$���ҳL�l�"^̉G~3�+q���&�����kV�w/�i3���`�3��G��aR�,��ҋ���v���aI�'�8����Sg�v��0r��pX��w�7Kuݫ��E�� �
f��ڟ��STU����	�K�F�6�-�ڽL�h�+�Lp&�)	���W��i�Pϵ�v����yxPJ��_���	��k��F��HJ�aD�	��+��^�)(.�c�� �G���#t���A�b��;[7�y�]��3�W�ϛC�TZ���,ɨC5R W�������[�)�h���Dta�F�����&v����C���Ãh�S��;pF�Ѿ��J#s4�)���l����+@�߰�=0���^G��'5n��>��WbO���"��U�EP�� �����NG�1�0*��QN2��L�Crw����ٲ�Yz}j�o*p�3�ؘfY�<S%��y7��H���d��(�h�!�˞������ݣ�/み0��{��T6��F�9���M'�%��εn�c(�6�^��J���y!aK�S2j��aR��T|�6�s�_z���g��
��Ò����.�;�;e=�K�4X�;�0Y��&tƝ��ǵ~s���n��ᄾ�>z�ލ��"�z�}u�J0���]q��b�˳7�OB=��	�j.���-!��<Z�o�� �>K���P����o�f�Un߸��"^�0�~8���j�^�d+����{��8_�xa�c�A-��>�8ŋ���>Tt]P0(`������f�KQȅ��+�Z�a���B����ٳ��KCk��&¸�3��~�v�2�!�E�z�B��u�O�����f7@��h�֫[OǕ
%4Q �:�Mq=iu8��>	>q�S����n3AV���ˇ7\"���i��]��I$H�J��Ö���.;�������(/�r)�**I�o�	J�#��y!�%�����vM\�An�$�c���Da��)<���~��Y4g�gl�L7��42����M�
�+��m�Y� ׹lZ�����P�1?��U�푑G
;��|�xZ����PԌ[��95}��P�)��>��زb/{<̘�ٵ�P��10T}��Z�O�8d%����,�$�o��	�@؊�K�D[�\��6��a� {��U&�jǁ;2H0q��J�D�@�םVY����)�;`��A/@�Jn ޒE��-�'m�qC0�m�H���(nF�]�Q�%_�'��.�2��wc���5�a�՜���(���z֮�� 5�3�o֣>X��A�����=g8�2ʭ��#��֭���4����M\]�����uu
b�mi�t��ׇEG(	�q��b��5Хj��~�)M�����}�m�ؐ��C���i+��L��c�m@�2i�6����a#H��Iۺ����������.��=��BG�H��{�nj��Z���d߁֠�5�^s�BH��(������d�{����E~T��ޢ�Rʿ�+�A����?V-�����v�S��|�a�j�<���q@X5'�.�=	��� <y�t�࿽�?$�w�a�@�/�����ݭxIKN=�QC��A}t���\eNBU���e ���u=�iu@g��r�������Dx��w6���0ō��h}O]�R��~��b���5���a�	�V"F _o"t�E��G�b)&��v�����OڕJn��yy�J _ X�CƧT��6���o���ξ�)�|$��jB�OK_��j�}�xJ��m�����L����[)�C�Zv�T�+8����&-G˸��w���{������G�p����q�Rc3A�α�~0�4N��-l_S�Z�(��n,�}����Ņ�O-�o�jxz��I�ՒQ_�cm��̗�h��L�2�v��#sY@h��s�u6���:q�
5n>����=�
)�Mb�w��b��d�q�jHX�yE X��q}�:z�+U6x�,lIi@�[�Jw穬=�:S�ؚ>Yr�kˤ�J�ׇ�!���C����^5�����9�����p��m�I�Vذ2��Ѳ����_s[z��	���Wws��+K�Q�}���;E�g.?�*;�h}�����w�8Z�Ŝ���L{B�C+��%d6m.�f�,�8��i[��_eG���v%e�!��ϸU�!Α"�W0��Kx.�l!�;OQ�E��5f"�&Vy~�Qj�-���^M�2�l��V��IZ���E�V9m|��l,#>�����a���zZvlX������U�8��붏"v���ak(c� Ӻq�"HH:8h�;l'a�1��s̨����b�=��|��M�7lL���E� �
{P$���tSUz�U�*�&'p�p�҄�:X7�b�P�ȅ�L���餙��O���g���&�k=�1+i.R����J��fQ�ދ�pE.���ψ�|8	�>c�=�}�P�� �?<Mo�<nm�1_'�\?��F��L�vs/e��S^��j`c������֓�#vŕ��v#�܋�	��gT4bＢ�cӫ����&Q����G���1M^X�JXf�r�Y���oӳ�D��D�,g��bvV1�E���Π���}��o+ %��ʶ��n[�'���u�&t�m̷��W�ֽ=�_����`f����@��)p_��%��׋����v�����0��M�%7��Ij5P�����)7����� ���ëm��f0F?Dׄ�¡��dӘpy���lH����hD��P���U,?��g~��
OSzF2
5?����H�9�{_�Fjo관U�{�hn}���� ��_�h�o�&�,�����3��P�VJ�)�����e�C���� �a˸Ym:��j�A�����r�yq�h��!�3�&'\��nn�y���\r~�\1��
E������tl�R���	e��/O��DpH�ej�TږYsVXGq�K!h\F����RD�1c%���*�>�hۘ%�׽j���J��6���q�^@�*�@�}���_��!�=���ó~�������y��f�=w&�Ǉԃ�#�ӡ9�U�����)ʌuK��\s���2���W�Y�æH#���a�3ϰ?��i���f1>cx?>��BUTq�G���!���B��9?�K�h�׾�?an�}��F)8�M�d���UІ���'�8O<Vɸ_��T�����&��]L�0���se{h�o�������f�V�,������%{�إN}����ř��fS�kζ����N�� �W�eF���()OR���ݓ���*����+p���푋)s���D<�>��~�|E��Zϒ��*6"�Ⱅֵ������n�i2��cV��;9
ȕG-A3��?�pNt��Y+���7�0��ŭ�r$[{���S�T���C��Y���Ԑ�F���0��zr��D�z ��#�eCq��>/��f�S���t�z^ciFB��5�x�S���6x'����_ͩۇ�w������ш�~��S)N��V�7����VO�����W�n�.�^�>�7�K?��S������OB�9�&+�KdZ��7�zF�^���P7�D2�7�LO�m_��^ط��/���L?E�,����@"�ב+����'C�S6.|�R^p+.'�H��̱��I���p!���چO70�A��*�q,�Ts��Sa���� _
p�����w���R��?��0ms�]>���/�j��<Kf|k�~Sɀ<��1���Q z��e�&ۘY�J�J��M���wp�3������M6)���XMp�1.��p��d��ʆ�����~��P�7�xnG� ��H����'� m#��L��(L�*�C�;��r�BZ�`5N��n,em���y�v&r[�G�F�dR��QK�����O��|�`=h.�����.u�����ޥ]
�kK�j�f�a��LU���E�����lZ���g}�j>�J�3�E��1���b��ř�>��g���&
L�� lcV������������ȱ��j��3��?���ql�FR�&�m���7b+~��.�#�@~��Jq7����!��.A���c�V��֩��1��ē�6��-�k<.�`q/�<n����ȩ�(�j�py����g)�&k�7�h�cQ�U�rF����$h~�s�J�F'&$��b]�M;�2s滙��y5�&�mH��<<z�I�C̅>�p_G���� ���Q���E��EL���,V�}���!˧" ��T'_v3�uB &��#�jh���.�&���Y3<�!7��C�a >.p�O)]j�F�99Yl�4��&1	L�N�^}�%���+�y�~�jaQw�M���7��G�y���{��j!��	���M�|����
}���%d�����;����T�}�����SN|@���+ 1�+d��q��v:j�ϐ��������D,o~ϰ���oo����1ʕW7�̝�}��g6Ũ�BY�;�z���Q�'�~�FS����x�(Е〢/�un3m`������0�`,�%k��o4x����wp�W@-C��/����Pq����������D(ҥz2���&w������˶�7�5��Ke��<~\+��e6r�hR�;N=: �o����;��1f��fX?q��,�i��9��>���{!q8`����=������91���cR3Z#���`�V>mt?�N��O�6S��R�~Sd��B�ΰ��k�v�L�{ҟ�WP��W�A�P��a�&ؕNj�#���R��7�ߣ�e#�c祁&Y����WS�K������t�j�d���	�Ҝ�}
{��yz�N��q�H�x��e摖�(.�����)œ��zLw�P�]<�
v�j(�
K����6�k����� ���E?V������b1�S��Y�*B�z�c��e�R�a2#��x��e��D�\��(O=k�Ns_~]�P�>��Z�Ա��l���E��6<���������y䩶E̜s�
�	M��kBn�U{�~����Z��a�k����Y���b۟�*qe�f_qk?vz�֍R�~�^50��g��H������N�K�b�v*Ҁ`A9C����2E������ɜB�%���)^T�n���?��w�*BvNZ�Ԁ��v=o�����ע����n�T�
Ws_�l ��������e�5��9H̓�iv��<�O������q&u��:�v �<���Za�ދWd#�XG�i$�<�9D\��"!~H� y$�ߑ�&�BC5�<XCi3~0���釸��͘�;��[[���1��ڿ�!�¾m��T���<N�~�vXq8����[��z�M��(H�+������ʜ��Q�T�88DZ���m��ܝU�k���Xh+�+z �-��#��ř[㹹�������!�rPR��x�Gq=��
���eh,�!'t��7� 	��qb�X(�|o#��%j��୽"����$�ʍ5i�<&�}0(��a�%����V�a��a��}��,��[+���>;�h�	?s��P��n6u�I,���|��'NO�������ᷰ�>��~&�TO�P%����Q�\W$�=��L����\ǚGJ�n���2��Y��ն�.U)'�fӣ����x��3e/K���|ۼH,��,�+�����"ک��ˆ;Y̄i-��.\3g�M�.�Rz�A[w�V&��@RA	��44���x��)�������=��M�_�)�Y$�2^��d�����afE�<<��i��F�����C�e�\**� �bDHo��h0>�$�G# �f�Ȗ`y���V5�'�	�"�ˤ8�G�6��:��+����'-��>�4�����a3��.ɉM���"�j�n�'�[�9+�pQlb�#�hR�_Av�q=@���h���=�v�k�3�5l��h1�Ԣ�9��ti���\�)��g�_;RO�6$^Ƞ[���4y����6��6JwUa��Fբ����!m`�A�&�ِ��q��'s[��&Иl�{�?�׻�d+OO)\,��P=&}��<sU��F}����#�z5�r��*Q�+���DG̃��<�I�a���kr�"8Xe��hw.�jJA���Y���}�G瓧|��&����*�>P�~����VΆ��M�9[�����E["�+�ӣ�B���w�%T��f���|�B/�����\�rp#P���)������@Y�p�������2Ѿd��u�M�,��t�����3�Y��^�����5�P�\EA���&O'�6��#�Mx��q_Ca�xJ�z� ���"+9�Mf���	���/m�W�%yw�x�I��;*�2�b��#��v2:�u �1��KH�S+GF���I�Ձ.�3���Е�5�y��[D���^��dn��>��d/��oV#�k��jN9f����z���ǢQw��4Gh�a�޳��R�#�&\$Rl�?3I$�*��B��?b:������~����-8{��G7���s��r��%m؅��<S�������aO��!9(�v�i!��r�S��(�B/���N�<*~���ʋʽh��ǝNl�B��9yg'YxN@q�Yi�Xi�w���DȠ:�F�	G��Ϧp�'��Bk�<Ƀ櫠3����?kn��N�Rš���@E��-�JED׊E�0��G�¤NI���*ك���
��)\��t��۵l�y�\���#����>$D�L�5KlH��pأ-f@uB��ط)�����9�|�7v}+���ѱ*�=&�D��k�a����{�*V��1Zr�)����py�B Y��pIzi��3�>36L����R^�$�1[�2e��祌��R�k6�Y4��T�y�