��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]���U���~�̀=�)l�X���!K��_���`���X'�Q�>�3��� �Q�a��-���w��t����$4��y�%���5���i�����Y�87��Bd�F�����Vred�0M��i8{�OK�Q�?��21N69�����o�RD��lK����%}"�����8�z���ٮ��!�q���&1I1eQ�̥��p�oB��.D���V�4W)|C�/ V&�Í�~��S�@����G�N	C�12���q����q��G�����_�ʊ������>#A�����i��^���j�,1n��g� D8p(Ro9$�6�'|Na��`�'�@87%�*�a&E���?�A#�p��W>�W��Nŷ�V�e]58_�����	���uI��L����I��66�O":�fe��oВ���a�Gv�b�Mv�W��p������U�� |�I�#��~B�p��D���I$�9�6��mb�g��hD.��zҐ^?e�Ī`�Z<����I���ɲ�i�w�T�J���d�/k�t-m�o��~������N�xxK�/���� %�8c5��j%:����s'z`P cs��֤�F��e�Y�};"k�:2��� 0Q  ��>T�A��3���jh�|/\`���UU�8�(�3����<+���e!h�ylՖ��apw��J�ܨ~��������yC�dv�Gnѡ3���qY:� ��6�n��!h�ho�-�<���r�Q3�b�6�J3������r�-5�������@�;�d�:�6�[Jm� ����N�����T�(���0Z��ΩP7���h��'�rιN4U�&��w�"� e/�o�x�gG,�����+����3E&M�A�Oy����SS����9�m�
��p|��5^/���4���F��UGn���/����6���j�G��|�X�й�W`JV�5��S�>DH=��g�i�"̿Nּ�n��6���ua�f��3�{��ʔ�O�T����94_4���.�0-!N����|�g?���tK���"���kD3�����ȩ'�8�`Jq�~ܻ�;Tᮄ�r���,�"�zf�f;=S9�gr1�R���f�''l%�)�E���=�QKR	`#|7Z�ݩ,'M�o���7�R��h(�i)��q�MS�r/��\Xu�' ����8S1��[A�6�TݦZ�a!�ᩞr�*�m�(�e����]ar2	�������ii�+[q�?�ͺ��/�9��/�ǰIt �G��=+�UIn��Z6"�
x�1ЪT|�!��i[JV��i���t��ajv�a��S"���H�et���N��N���01ـ��K �����^c�����@�"���XL�F@2�>����R5x�4F�}(A��� RB�P�P��;������i�M"`Th4Y]KF7G����DQ�����C>h�3�F4ſ�Vn���0�T�(��_�խX����X���k�_�Z�a2��U&�?v�r����#Sm����;���-<��N�hJ��{�CG�&����%��v)���˯��%�v CX�K�=�F��W��#>a�G�2 ��/F��J��M� �U�vpD6�N���t�2'��#�S[��u��NZG�����M<��"u �5�X��?�����k�!㾗	B�1Oe2X1��NL;�ن� ���
�ا$�j8\��ή<� �����?�u��D~�"�4V�Ҏ��e�`�y�׈hcR�FQ	��Q�B�b�����^ʌq��;�I���ɟߏ-$�\� 7n7<������-	����%�&���f� x�\���2��ܔ��g둤�]G�Ē
hܱ9�i�q��j�;j���S�}4u�|��`��C��{����HNR|����R�j�vQ��J,��V���3�ҝyw��>r��]��v�p��0 �V;t�G��ܳ�c�)�ãFU)0��WW�Nv����%;�'U���}4��k��.�M+>��'���e�$�U�[ߝ��SZ�oۼ��Ԭ�`�M����cю~}~��Db�[C�2�ݫ��bg��s�A�y_)��ۥ&kb��#L	E�u��A\�*�as����Ef�����R`S�-õ������)�k��(mwA����2-�����}�}Ȝ��C/ߧvC5-!&{>lɼ��|�¡��u#M��q�D�3���)�QA��`�h͢]�����#��q��v��e6�s	��e��%�!6��H�m�@ǆ��t�}*c T�`j�q��<K�\v�ʜ��U�|����%���u�[�X�����2@�Z�l�N}�xUc�喰x��O(Ϸ>��?�7��t�N=�{����7Bu��4�ޗ�=�f��<ȽO�_
�e�}G����V��euu�Ga��I8�����&ň9����!�$m��(>�0�I:<~�K�Չ�&
=�_8�HY=�)�Y�����2&0��_*t����`b�Z4�SA#�z&�/�����S@��>���9���ƭ�i���L	��!Fx����ڱ�!�+_��c����U��S��CeLџ6&��#� 7W[	x���1�d���B6��C��u�	"��Y���Ls�;��~5��/�}�Ԕ�O��'���&�e��R�R�Đ��2?��$��-����*�惨�_E"��)W�,����G�=���ף��.�L�e*"��L�&��i/]�~��dAeP�I��{#j��k�9܀RA��&�5��VUg2�i�s6�\��^?������9x����&�xHi�?�fs�!U�{�D�y9��qC1�o�YEMݤ�+���p�2B�Ó�"���j�Q��
%XW�_�����:����=Xx�2c��`]�+��~&[c$C-w�@��L���|�߈���i�9Y
=�+FS�uYPu�/�t�(3�>�s���]�\2�dg!��;S��R ѐ���5��(��g��t��u��A�- ���Co��rcL� ,�Ѩ]�(p70&+��`�޾�]�~]9J�!̃v�EO?�P�k����:U\v�W���9�{�0�,����y�OG�)�jG�b��Q��D���dk��ϡ&t��Z̙�gl?~��R������!Ċ� 4�8z�Q=��-�])~�1r���/�(�*BU�Ս��B-��p0�� pc;��Q_t����:ѝk��x&��|��-�t��p˚��{$�^�v�Fe�� ���\��h��"V��C���w�b[	�n���O-�ײ��\��W����G�-�,p����O��a��P�1P5%�	C(�~���jC��l>_�jF~`��N4m3m.-~л��"Aq]�%l�K�2�E;�C�
��]`��<	<�C.��D�������ǋdmSVH�_���WPǀ�n���41KZJ~��VL����R�T����3~���=�$u���&�e��k�T��7f��G$�Oo��f
��� q)��J���X��Tyؽ��%�p���g3?8�h�&ݕ�D9�,��P?:�ޞOSN��ƴ|�WK��;��[�?����ۛ�����9�� q�o�<륍�����2Ws��B���;Ba�p�N�( Lϴ�k�4g����_�7zV�+}��.�㧃F,��Ae�<�fp�#����Èc>i{������.�@;�9/ڲ ����p0�9��;���05�g2��Y��n��I��$J�KEa	s�w	�<�bK��0�~E�H�?-��L�4^�� P�������L���-��"a����W��!+aSWRW|7P�Ҽ-ʴ-��<!�V�����F��{.,Fn�g������r�ƾ��}�i�7X�("|��Lr�i����cƀ���0{S�%~���gJch4��C���*a��i#���3I�j�ag�D?>6	�%6�5��9�[�MeȲ|:e�|5R�=��fm�c- �Ԧ�3�˜�]%Jy�W,�-y;����7)E�ė�w'�I�WL�=�8��N]�[O�{���N���;j��j�2��h�'q�dV1�8��տH�����5����!ҍ�ӷN%Eu�#FV�����6��9`F]P�gJ��l?p��O�I���;����gl�H�3*G���yMR�RĜS퐞bV$J�T�	9W����<߉��%Ht���	h�0��Cc�&sw!�$�/�R�����(�J����/�N+ �<�J)�5/%G��� IR� :
'
�~���<TR�NW��|!�f��f �!nT4��~�����#��hD��\i�� e���Z�o��Q�p k��"�'���:M������һ�`��G�uW{�ݪ%1�f�6;�A��p�y�߄����$��ƒ=���9�g������������<��`��ػǍ�9�R��0�)�N��(�q�/����~�!�G5H^�x��׼RX��-�2���̿�s�܆��;�\�X9m����`�C&�ư2\�mB�����qh衟�+�90E�m�3�P�1��P̋�̰��Z���wk�O������^�~�5Fb�L��]|�g�5�-_�6-]`Y�(,��E�о����K*Fk�#jG���ܽah�596A~��0�Wg"0��ٺ�,�yX̊�R�С��#sN��(��&���Zea��Dn�.DQ��E~�R6�6S�xjK��@�����W���
2C"�ďM�B��n�5�<�@$�!Bv�5�r/t0���%�M�����%[�������N�����0�#��F�c~�B� &`�Ղ9U���h$%��o���q�%�V[da�6G�nIw�{jzj}@�����ף.#r�j�k�t7�y6`s��otGTb���ɋA���*�A�w�<o��̨67�_�P�_��g�_�փ�B�<�v�s�u��;-@L`U�k�K����}�ak
����J���������F*g@%�f��9�q}%�o�����z���d�0�t���0�?#G�S�q��\m�Qu�5�.s�ć2��I�K�b��+�~�i���ަ�.����Sv��������M�7��T���B!�n���U�9�dK�<�4`�ͣ+I��	��i{��J���}O�_��?6+���\�ihvt���fH���1ϗR���޷,��bS�%kη:z�'����ڻ=3!�%�
���k�v>���+��u��G�fC�<]�M/� VU�͵Nn��@ �+��-΍=IP�!�%�ґ 
�s'	)�'���i����� ͛�K��\阨�����M��+Y�\�z���;��!*� �B�פy����o�;���Irk|�4�ѷ�K�_oX�t%8�6:���p�k3M�,l.i��F�c���P�zܚK��f�;3�X��Fs[P����Y�H�2TU��*=#��5��Wֶ["�\bhK��
��]���	~y�1����!���; ����*6�PcGk�6��ג��8�!����T��n�n>}O�y���?��ni&�ޙˏ����Nr�]���L.�D|Z���x�����O�%��|�}uR�'����/o� ���S�;���J3��J��ބ�1@t
ov$��0���G�b"88��4�=L�Q�ȍ�/L+�Q����UD��o��G���6�7������13.����AW���c�T�
*b5y�.��%[2�
�i����~����?���}�K1��|�D��ߒ�.緒�B�t���߼�������E�
�(.�%�q�l3<C\bC��
Ė�$Ǟk�\��K�g��C��$�^�kf<č��;������]1n��z�T������,���4����]6��:Y��Q]����V������B ��!CJ�2s������Y��������Z�`���!�%准pbߵ�Z`;(Ou�1&r��LNcx��_�]�ZT>��e��[�E�oR�*�"�r�0������L��Z�X�-7.	Iܾ@j���V�
��M_4a��c0/���2C�(�~��6�v������ �P+U!�����a$��+�ܽ,ۚ(�w��hD��<)���5��}l+�icx��Ǭ}�2��<.���ZM����ڹ32�.�g��S6�K[� �"�6u�e1F_����������`�MB�o�1� �p�C�Y�uqѣ�':�泻%���I���P~��Zxe�M�qũLB��k��y���=σM4k.�EL��ck���TN\�Ӝ��}l}�ͤs)�.E[Ǘp��,�	!A���#�e$�B4��/Y����� U_�r�Ba�� �8��� �@&@��s����(���q�+����������U��\4Q�;P����6)y�{e���)��EO��ej��=1�n4U]P5��S�̉s�~jn�#���FC�t+xPf
iq��~�C�`�8�9����rdP{�L[?M�%h1H���W�����|��v���+�lb�zK�?L��(��D$d�D�f
V����m>�A1K��˛u������ֿ���-80��nO�"-������1}PB�V�B(u��FZ�#Vϒ�2#�Z递�:l�,����u%>���u���0\Aݼ0��x�n��L��+���7C�+Ef���J׍䝊���$ތ4����"����C�`�1�P}�˻�\�`�I���M��R���]��[Źgn�^�z�aY\�A^�	UYp�~��+��R�u���G�����s%%��Պ�|��|�����|�����3-kF܉��	(ŋ��qxV�d��KY���{dm\]_V�&��-_����9a�5M�v&�E�h筞(#�y|������^�,A�t�����R�_��:���g�wf#�e���#.go�|�E�Ӽs�	���B��!�IUԳ[u�VE��^̌���ީ'28�64ɳ�0���R��=��&�9e�b<l��.�ˠ�ąB@O�ׅ�����T�g����p$CVth��	�6�:iS��=�D�{���2+Jfco�v�U��ԋ���%i��� �&��A@h�������7qb%s���r�M��$ᣋ���tM�!�e(�r~�8'�#w\Z����h�������`��a�x;��m�d8�΅M��8�Fb�QS����x���N
,������׉�"�U�%�/�Ӕ�Ō����a�]A!;��(b�-lk�q[����:�۹DZI���N��"�ewU��ǇWUz�w���.u��#�6 $(X�M�ԟ���>9�GK�gɅF�'O�v���?�?	y�By}y�M�$�:�\���@��K���xTG?�&�E��W��<���}]�|Ϊm^��RM�=��;��R�~T<���ʐ:�ۘ�w�v�Ԉ�z4������	��N����&��Ĳ����������?�R}��������@D��f�/����`"^�"3�`{]����^����sNʃ:�+�~䥟S�N�vsꕾl��j��
5Q�UΏ"Ɖ��J]�D�Y�-n6ZG�G=���������X��N�@�M�>�χK�O'nF^���I"�2��y��|�<�u;(�Ʋ7�d�x�����~�N���~ݷB�C�C��N(� �M��B�w��J��]����4�J�hO��#��v�5�����A$E���Q<#�g��!{��51x�~�,�4���=��tF���V�z4��YΗ���2L�2Ϝ(~}`���?��*�&��Z]3	Xl�W1垰��l
:���+Z�%bo,�������%�$r N��vZ^��ˬOkSe
ńd�dS�%�qy���HMY���uj{b������ջq��i蒝��/2��=q���5g�+$�ן��,���O�(4c<r����U8F{܋��E��a�V�9	����d8iU���wy1�!	���&��/�Xa��GQ��
��{�`^��X^�����kw��g�R�{/]��l���'T��E�2.���BË����}Du%1"D�/���m����$Z�W�=@�qc�4+zJ��g�Wf�6����Z|�����=���r��N