��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��V�^�Z��i�hW��1�%:~c�"N��˹�wG��5�H�
�P+����ֈ��Ŀq��5�d�TDe&2��xS�\"� �#D�+N�[�ZU'6��s�ON��� d+Һ�޵\�"�J�б�tz�����vk3�^M��q�T��Pg�=|Y0�1ޫUX(�7�'HuS��Q�{Q8u�$��-|9\����l�5h����}������:�#07�Rp��+ yR�@7�f��uo�P��~���H�w�� �%kN�O���#;���@ѓ�?��[OK��*�Ms\i9�#}A����^3*l�ۛ4-��o��W������E�\��z�yc�n�6,X����ύ�h	����C1����n�������Ɩ�5��S�bv� ~S�m7󯛋��M-8k̄������;u��Fj��K"Gz>�-YZ���^TW`�z����d���"��f��Jy�1Z��{*}�Ut\x�I5��4����t��(���aޅTg��/}$�m�鞩���ZTl�L�f%����Ü[�z*q�WB؜N�3T_ӵP²b˞������f)�����e��ۋZ��E�\r�w�M��ǯ+�(�J�K�{v\z�EҰ]!c��L[5�]cDs�e耔xN�B�9�N���ՒP+)J� 2�/z��mD�5|?5�4��Zs<{-Z�V��nd(4��#�hJ�Bl��&.-A�d1���Åj��\CV찍�J̽p�k,�2����(�z=:�ý��4��Pa0��
RK�՛�L�eNRD��Q.\���M��w[X1@���vנ��^&N��n���i�+�Z����� R��%or��ki<͟�	�I�p�@�l��XȑY]� �d(�L-��h
��˝]������K��h`�/���/]1�n�<�I�yN�L���C��V�r�׀���ۭ�����i��r�T�'Ճ��;+����*kP������i�i���Kk�z���%U�w�a{M��F��VI\��ǵ7����s�I/�I�{�3)�Lv��l�^Ndu䳋��芫���8��G�-��J0�uDf��qas�f�|B�H��@_o���8;3��b$Y�ŧ���C�!�&;��|B�7d�>\Q)���W�����)�6@��A"/���Z"O�	b�zY(JCwv��k�x6�2m,�d�T9<������=��Y���t�00R��������x�U�\�:�{�/�64eUnk�<�仛A*�I�]9���zy���i�?k��en�H�l�g�>@7_��w���j~����A���9�݂�<�>	�əF���j#;]m����wL������G�c8yw���g�;��Љ}����ո��Z.�ח�?����g�$`*ɪ�`V5����ѭ�*KM~R�~^�Ǉ�=�
G������Xx�s��x=9�z7�&n�`�캡B�񴄊Rg�$���� M�
��)�q��{17/�ĬX�
�׉�I�N�����(���7�8_�NL���V.�"�Ru�:tZ稁2Gm��օ�����0/~_�>c��Ӡ���7 ��H�Ku7|��RH���������_,��i��@�����%�"�����k;�^�sOu�aU�$i�U�Z]-�.�47�¶f<�m�y
Z`�H�̩�l~��UM��LɄ �Ɍ_<���*1DFr�Hi͒FL�11��P��'��!`��jT:�p�$�x\����$�y���k����8�������z%�=�׸���x�[�57��W׉����*��� �7�d��^f<��e�Ji���7!9z��+�M{ ��B�P�$�b`W=K��[J@ԙ�9'��+�mT��}�f܈���f�5f������rԃ�}GI��MI����4���~b湲N�N�"�DaQ��R�֒���q�??�m�w^f�)h��KD�vL��o�����?h�~�� 8w��E��i^���O����-�m��J5JK�z�se��l{�䆋��%��w��|�9�G����=��T�4`����mi2ߖ���E�az�.T�L�	��k�{�9��#���(j�ɿ �!��DµG@�l�Vl	i~\���cؔ�&t;݃���C�nqvU/٘��gok��P�S:�f�|���t|����N��`)�4��@mw��y�*����ب|��n�PW�h]{���|I�JQc9 :����5� ���~��xZ���Va8�;K�_`-	{C�"�v^��x7��F��k�U���>���sN�8	�'a����Ϝ�v�Sfټ`������4!���Ί�[�m2[l<j�c�Е���HV}�*�߀��G� q�3�����[��C�qn�K��81��%`�*Z6v�7[��w���Z����}J��c��p૞����c�P���
�po�㺏.[,~CnǢ-�!<C ^��sЋ����Jˮ�<YD��g��]���"N����tq���bc��x��wA|�NJ9#��+�*�q^��-��bh�Z�_x�a�qN�u��dq��K�K+M\�NZi�tR̮���_|g2�p�M��F���W���~�k���O5��7�'y	7Y�����n����f\�ͨ�S�c^ʊ�*���0��n>̛�3F��YO?���[L��JЀC�Ƥ�;.�%lU�_8������ [}���a��_�*e�͑&�+���t����Ӗ��T�#4��)�o3��D�(��]�b3�����>�?U��m��x������st*ծT=N�MVr�6�-�{�B������o0X�?�ГD������f5�CO�1�`�;b,ʵ����o��G���ȉ�t̑ǭF����%��|n4t^;�l�<��LoF �n_;����+���̪|Ǆ���X�zK��� �Y����`?��(fT���Y8��:�E�u�Іz�nA����0�������Q��~N~����_w�$�T��Mv+�T��,��t��)��tϸ����ppz���}����Æ�712N�>��	�f�:�Y�������M��S��F���{[͞+t�B�f�V��J� ��4^3S@8z{cb��J�u�F�'�y ������g��N��pVG�
%-����SKda���^�:���)%���XN� ��w?�8���k��h_鉋�0LD����p�iS����=ƭ�
)�\G�1M=��J,��m��#��{�I.����bu�LA�6p�s�|l��X�G�ׯ�'EUw�9��''|;��%c���'�⚭E0�h��p��}�sâ0x��t��e@K�Z�P	��/�b��Œ�g�D��Ο���G���3~p��&XTr���؎�����5Gв5/.oعt�,�+��$5�	eT��R�%W#�z+=�v���W���m��B���m��n�nT�Zz[�� =�|��'�b=i(��"����L>`{���Ǚ�e-�mr�.I7��ήuH^��վB4���vn��W�4���+���#���g�V
���h�_�ۧ��.`\?<f�9���ȇ��;P��v�Ŋ��7�Zv��U�`�nоs�� J�
��`�xY|�d�u?�K(敃����A9��!t��ٿ:�"hp��{��`�� ��[��ej>��m���qB.DB7���| ��.��i��2�Ig�dUz��iu;��S}b�V}?����I����nN�lК��%4e��[Z�\}K݊�7.�/?��A�q��\��)�N��䄜{�gƙ--�U�Z�ER6j��ע�k�>=����yF��A����T����6��<Z�&<VZ�9�˛��n���va��+�yU��V��x4�Ӡ �3�oBhhm �.l�[�J5C��Rpd)���3��%��{�'X�@֏_�5"��yv�'�A b�����$wA�w�#6պcu���I�����������K�P��C�L���:kU���l�}\�T*���zh�I���냐�$b�@��C{87�S����!�8�������>���
�cy�Y�2�irD�J��{����k�<��]dB�Oi���oƞ�|�UO������d��y�AޔW�.#s{��{֗�{��\w"�@���]%ҍ��o��.3�k��V} ��:��,+d) ie�3���%�AO�/d���짧�� V�L�� ��hxb�;�qHO������c��A�^�W|��^�$��l��
b����a/�f����(;��c�j��=��"��m�KP�a?�MC��%]bg1��z�#�4T�d:�{��!�ALO/̬Ɂ�*��||�<u���MV�.���,�	�X�ō���s�?k�oFl���X-p��+1�/ō!\�L�.#Je��_.W��xfs�(��ݬ��8��V�k��ԍ���Vޅ�������I(�˭��jP䱕�5������Bdu`���e��t���h飈��]����^��%HC�N����ޯ�����.�Rt�;%��Y\�C���N4�M�ɐ�Խ�m��)�*Ʌ���a�ӻor�A�^�����SM�8*i<q��1���:W�F��wѣV�ÖȢ8��]T�]+��������ٖb<{�H^WD���
�S���z�drunjQ�:��+����5���<u��;�RR����8@�l	��p�����!�d�\Z죆yP�\�
�2��XŷW��(�WJ��/��]��B��ѩ��� 6G��uG�kI��N��������F����� j'�����YW�H����Ґϑ�AG�$+��a8@{!�{����({lWl|��~n0�yn���}9��y1�5���T� ��Ƙ"���e�]����1ؾ�O�BU՟�=AG��<+1�F-2Z�����=n���_�G��i��ѐ];:u��]�r���n�!�b��l_��V�;T��9l_�ae/"׸{BYG��'�?���Z��!���y*���(SO������.�fм���l-��8�nn��6��ĀB\����5�i<�䈦:�^G98ZO�c�@X槭��R��冸��c�F��xX��R!^vڳp'βB~�N�Z_�M�(���H��y�Z�2?++J��>^��H�#��;��I%#C�Ohz����VB+e�#W@�U�i�}��;Q��zɋS�Mj�'�����G�%��Ce��q����鶻e5�0������� �=��3�T���΅'�&��{RC�4.-��5}�f�Z�V��!���&��:���+���H��l�L`N4I�x�,Oڵm�I6��o���7�ڵ�b�:Bӓo��7���zzeU��)e,�O������k�����*�M3����Q�i%a��H��{N��t����ie�/�%��:�UpTdw�����^À�=�`S=_n�d_�v�ڴ�?��yݩU��F�1_��P�~+���%�y\�(��n.�AL�edh�mʂ��"=���#�ª%I�����}K�R�I�����ق ��!掞�R����Kb���m�^ñ����!ZTf���p(Y&��[hJc��S�������6���&P�?~|+�.��%x�x����`1a_ �?srB�Yy���K����p3�MT�(����6c��-HSb��<���[g�����~ΐ����b&�]�����rl�N4eA�${�3�	&� Tj Qa��S�<������>Y_�A���	��gD}�e�X��@�M;)%lX�)�/���W����6�p 7�m	'-�#n��x�;Liǿ;�2�����b�h�\��H�WP��M�t�%yy�y�7
,?LZP����d�"�T�m0���Ƕ�8u�������Nl��b6a� ��F�o*��-B�e���������s�`�T���[�jw��;��|
"�:~ ���#r�+!�É���S�6	T��yY]||c:[�G��W�cm����j|aU���ur�=�X��]���e������,;�$i�m�싾�Y�[Oߠ}��������n�vG���VZ�zdzPZy�MU���:ŧ���z��~��`ܩE�/F�@O.��7�e�%�W��]f0R��|��c��D��K�οɩB��5�o��"<�A�S��`�O��~�ր�_�� �Uh��玉�<.�`���nr� 
����|����@�z��>��t]�vc'p$�D���pe�DP'Y��y�/0������$o�����	�`��PY�ٍ�L��&
ol��wH?��9^p7��A��jF�����a0(�H�g&xϊ`WZ��v}�4$�&��/>�]b�	K���P_�&�l�ʦ�8����	:�UQ�a
��*2�e_W�����ݯ(�o�6{K�%ea���OP�R0`��j
�	�)�(U
]�	6�O8�|Y��~p�>�s�����������O��Mg�����r.��J]|c���9s`:��Q��֗�zڈC�b���ҁs޴��#w��r��m�f�K������7���������j�.I�:�3Hˤ�$��sZr�4�i�|׵�����`��Q�V\�����|��}NwҘ�V��E�$� �:�p��>� ������� a�����v�j���p�Ѽ����7��a��\����9�����8��p
����	L����5<���6a8�5��!1B���[}�LE����;���܌ӮC�9�K�s�w�hCS<��x%XbѢAv��	*c���fk����s��|�U�c B����G��Mk7����O �����/!8��p'e��A�� v\8͡�gI��HA�c���B�<��_|+o5�A�1�G��$Qi���bX�͡C��mU[ĪP'ڜ�O�=�&q%N�s^��cv��߾�R?�N�dԟ$����H!psRB�3��p���!X���$*|�"D��� i��\�<�i=�����Ń������Q��-�c��_��M��"g�`A跣��9������f>��1K��"Z(���l�����#_��Y*��t�ujl@�l�~�T��6Z�B�g���K�!�"��R��k{���M�T�*��Ù���(Ys�}�p<0�3��zȹ?{���e:,d��V9�?����*�=ѩ���7�D}���R��EL��O"���5]%)^�q��^A�=��
Z��3�gNP�/�l�˂�Blc�)�x���̍M-2�[*�4�A��FA5(�8h�t�˧K�s�ɼb�|LKCO��]���^��'���¤K�g��ۛ)��qp��F�D�Hǖ��+��5LG��
���Y΍x/K(5=V�?]-�t�Wڌ;a_���$��vK���ad��������*̡�y2��ʺ_>�=ۊj�b��W5%z;�=:'�B�Vc��=p�=�~D�ۂ��!�_$JJ���!�m<���1s;�fCҖċ�B������_�ļp�UOM������:�Ŝlpp��pL*0��8�e)�pz4�����%�s�Q�X��ZF�zh=�pF�������
!�� �h�f}����?��;��nu���p�S݄G�c��^K��fK�絵˄���P��g
B��=)��QXq�n�������Ս��_}]T\x����(��ǹz_v