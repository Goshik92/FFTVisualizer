��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܫk�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�gߎ[�zZ$D�H�=���3�r�-�7�Y��B
6����I?�����k�'aQ=$ X[Mo�o�����o~��P>��]p�]�9��D���M�y�~I�ʘA��l%�T=���溟q|��iN�NL��zH\M�I���u��L
�{��D 0�w��h�g�>%����2��*u��ПmX��)����/�̑蟕�H�����6[_ �oY&�,P~�
�c��~#�	�5���6VCA�F�_/�c�o�9JW�c#�Et&�.�Zv+^l��!����NB��>��92�L�'�ߩ�Wآ'Smf�8LH琝i�iݴ�`")S���먕���N���t,*�e�^�Ҧ�
���9ӌ������O.EE����J��h���~/ 6�û�p�r2���v"��8�V�u>��#{��k$ݺ08Ls���w6�'c����O!�M��:_v��V$�����8	�&N�գ�a�8�^����[\�Y�����־,��ْ�Ҕ#��]��}?
F����@tFB���Cc �V:�����5gPi��CJ�Ҝ]�H��q]�f�n2۶�0B9�qXgPA��I,3Pj���TyK���Ww�Bu|̳ �˱%�_ަ;G�dT�	������S���Q��<��*���_�&����������\�Y�X�� ϕB����9@�<�=������cM�x�����`j����F�j��d�`�gx<�"��C�R6*�^{Ky,2LZ�g�^D�>�~���d�_)h�(�"r�~�4�娓�^@���F��II¸<x�9����[ʹ^OFS��D���ڴ��qR��P�8bG��,3�3qZݡ��j0B�>ݔ {����!�)? r
ť�\�B8�>��W�o2:���D�E�~��#��l)C�yC�S�vS�bR�.]�w����ÿ���Tq�{"5�\��.����Udj������6����?�������L������w:3|oaz#����rkr�2ؖ@����:�hK3R���_W9�i���K��}x��5���ï��+�<փ9``�d�W�[���kjS�����ټ���`4Y�t;��mGG��*�H��� #'��| �EgUp���)�gAu+S=�+nz��O��*4�4b*�|Q��Ls�2��q�n.Wl��!��Q���+f��-ƈ���{���Q�=����Vdl"���XMPoZ�5���������AK�V���'%��x*ʰ��1�Dn���-1�ĽJ�i�l���=���p��o�������&-�"ς������5G�q�	 �A�fs�D7 ��H�<L*�\7�$߆���y���A�c��������l(��fr�$�sw��7L�d��"ֻ�^��uDmQ؃L��V(H�%�l�-ыW�D_�|��*q�_�ie��DK��2��zb0����9�_��YQ�n���5���~Zgc���yO�D3Û�\��)��jR����@c�Ң�[�::O �yyx4�tY�.�^1U��R���i�~�Ƞ�������H������~��6Ъx��A��5�P��~ǀ!ϑ�n���n�/([6�r�+��zqa Y�?M�_Sf$-�6t.��{"h��	e�\�#!�c�:ZR�*k�E1%,5I���N����P��Uj�
�:x�����W0�u�3LJ����Q��)���l��"i��s�jΐ<R�X-#1�)�A3�)�L��=�;����cK��8��&��'�C�Y�+�;ܸ�*G�>���Ϊ�aٱ?�".�����~E�P�ߘU
 �\�)��zAM܇mxc�4�W�2b���ݔt67i���R�D���T	'Ș���Cl�8��EӡoaY�� 9��A6k��N�h�+O�����&���,�D�֢\�� Gz��g��eN? =�!Jm�"F>�34i�J���q,�6�+�w�a��z�A�>�h�v<Z�����VN�\�.���.w��P���!0*in$T�Eg��H 1�)̳O�:������l�x�z|�i�SaBP��W�� N6�Ք �4"-�0�n��J���ö9�# s��sl +�gv-���#�3N�9�Кq�HY6k�*��I��H+˷~I���4��8p�^r�EĪ'�Zkmq,�u�A��͊��<Wb5Ke�q��E��|x�~�pqڎx1�ϭs�+~,�οV�Ɲ�E\h&s)�DE��%�;y̡p�:ݨ�p@�T�����!�W`v�������NR;Ob�i���_O4��2c��ع��6������̌�p�b�,�����O�K�Ӧ�>�EķR�����ie�h�e���Fx�����mJ��Q����[Q�(o1�W����0����#-��O-ВC���V���09f�fBU�)�I������_�D�rRw7�G� c�n�FfNK�8"5Iz�@�d�t��M���<Xw<{ts�{w�B��P���p��PG��n�O_����_ 3t�����y2i?��['�X�Z�\���#��:/�_��H]u�w�Ɣq�ܯh�
Dߟ?�
.|�[��,I���*r��\/p�?���y׹xؼ@������84�)��"��߉����Ҥ�<
r�no7I�F�v�w]���!%�̔�i���?)4
%˅�nȦ���.L���f\��0���3��`��{J��W�@ � ��9е���AJ�����gO��v�0>F�N \�2@!�I��
��ah��m�^�wX�u�˜A�������79���$�@ixxk���ٮ:�3t��3KvZP���f��/"�
a�hJ;t}�<A\L�i������?�z��ʠ�&w���Y7e��1���]�y�<�(U3����;V�(nֹ0`�"� T��ݺ2PtE����
�m�M������eG��dsOY�"%��z�,�������ձg��8N��8n�lt�/:mF�|�*c9�l�Z����ǆn$NK|��1g��}}/��1�X���j���~T ���T%;�ʻI_4h{jE��ɠ���e���ݟ�:e�e���������aX�,X<�Y�5��8�{�:]� �o���F���Ԁ'2L����3�'�~���'�m��q�(��fk[3 �>"��N2^�i�b�g(�����k�����<%=����a���%'2S�b�&A48�DV9Ɛ��N�{�wԉ��=�$�L�豣�e�Ņvi��t@ ����k�AM_�H��7`��f	[1 ��r�d��L��UQ:󜏂]m���`3i���\���y�?�.M����K��˨C�ϫ�*��z	mZxz/]�&�l�$8b���8�-VOۧ����T�j����Ќ,�b��ޙ�>��6�	���yGO����87�B�cthQ(������l��v����D��1	5M.g�z��YT+B��y��8ݤ*1�س3d�i���xC�>�,�W?���nB�г�&pF!�^����e�Xn�0ԀS�Vg{�K����5͑�1Pn���I�N�[O�	u���d�/�":��<Z0������&�IE�"���և�{Ûߩ<*��<���`��|SXl2'�� �ϗ�������y���͆(�&E�_"�v�/����ʐ�n�q��&�َUVuĔnƉ���w7��jQ��)��/P���rK�a��F�#`&a�[x&dNX�V������:���\��s��bMT3��Cy�P^����sm�ti_S' ���$�{h�
�����h2�q������5�@�n�u��޸���Ii�jc��Uo�u�R���Ũ��r�c�!�S��Qa��~|��f�>V�)k0r�1�
�T�9��o�U���X���� Or���6��Q8�'LP�Oc:�;d��1��͍v5��~���%R�@D�t�I����R  {�5�=e�����#���r�d��"'�G�mb+C�6����o��zZ�UM7�n<oa�	U�xۄE��7,2�����fmR�%ښ�%Ʊ�>����'��c�V��f�掟�G�k#�p@�ݚ���C<�1xv�F��������ظU�ƾ��<VP(�5qc)�ɗ���U���� �4m֞�Q�e�f�#\����}�y��A.�ך�G��0ۻ=7r��لC{h��e_m�1���
�H��	O�M o�Du=�s��:�{j�������V碬�%�V�+#p��a�N���+��ƥ�l�(�����+�	�V��F�L�	��L�VǬ
��U��Ϣ��]?�4��?���zH��b�F6o@X-�*!N�d�� ��׃�o2���m��bP�7C��Q����rch�$�)"r���4�+ �6��٦�m97ټ�ϭ��ڊ�����=�n� 8y�G�y�}4��Tp){H��=����G�?՟�����?y�-Q���;�V�wp*��*O�?\ݟ����Z΋D��2>�Ii������#�S������������:��.P��|���Q����8�Z�k��|&c�Κ�\��F>���O��d�uMw~����M�#�_U1��e}iD�iH��^���G��P><�y)/g庙��}�Pd���1X��$�)A�L�w���$��c���.�&�	%0�P�q E��X/�
l��X�jM"�-��x(�[5��I˥�0��,�ͅ8k�������;h�Q1��ր'�[�:�OZ������^h����o��C����M�B�z�>qߵ~�"��[F�H�ͪ�64+3N�y
��m�M��J*��m#hQ9�� ��JRΡGr��7t^��XUհ�O4X�j�l�?f�v���/���e�qpl����hR��V>H���H���wY�Q+pē]�  ������n��%#gYz[���B6r2_G.v���9�+�nPډ�Y�m��⺇�1:���iQ6<��~�el��Ly:ޒ���б�b~��-�6�H����G�-�]x�.ϓ���Kr���(vy%S�S�%��V�F�V�]����R�=����zhL��>�fi�I��%����>���t]e�03���q|�����D��qOhV�:�b�FP�u��!"E����\�kXF�*`�nݾ�S(_d8�ؑY�fY�y��r��egzM�k[��RsH-�k��.1Ho���`%�F�[Ü�2�}ӕ�-U�}o(�+3�.4)������o/>U��f��W��Zgy5���*�]�N�F�$��QHm;NT�/URt՗�\m����$��Z�/M�7�P��ⷞ\�\"�Dt'@��4J�QXd�me�l�s�z�aO�,C�F�� �G!�s�̽y1e/�o�vz�ہ[?3�r�=����*6p�$��ko�j��{��k7L-��}�ɲβ�#�Cݵ�@��sz�B���9T%�l����
��c���.�aΙ��e�X2�HhZP�;g����Zv��]e�f�8�x"|�
XC�>��&Q�K2�o�s���W���V���SY�E}k�G���7{�A3��kʳ���R15��E�,Β�r��q�8��Q
l�~�������WE�EK�r}�e�T��u(=D���R�66�:C��R�i� ����mˇ���+��m��qT���\3�8b���Pq9jń��14`���
���y���F��wa�t�!|_����Ae�b���{L�⯰��Ĉ6Ȓ7�`���e�s(r��I�Ԍ�-��Ef�(���-`�	�
ݜ��9�r�M#3X)-�����v�]�\�1���܏�L�D���HV�"���rl}�7'A���^���h�ؤ�,`�o���VϑDC`jP$��"�_�"���{ޡ��k�J�@�&�U�ެ]xX:���II�j��l��/c׽4�vV��i,v����_W��t��q��<A�ʭ!a�M������?������ϸ��נMZ]r���
��Wtx�M��ȷ5J��aٰ�� sVm6&&E� ��H.���I�)�䪒�dY>طM��0�����&�L`�	E�qJ��{�ѻR[�<	j�G�7��ݔ1\a���J{�����4��;��ɥ�!!����D*vFH��-��Lr?\��}E����q�]3Z����vj��鞽�]�����3��V]��8;%��(z�HL�Ҹ}�s~��w�e���������6�X#����Z�-���=skF���_�!�4�/��Ʃ*q�J�+G��K�Ƴ*�Ju񎪏���gwmK���px��<�w�`�<�C�렟��h6]�a��VU0Sm�e *=�sf3#z;e>�.;� ���G��tc������I:v�vxV���dS��'���!(T�Z/=��M���V��=�^0���<��s?&-EE��z�<{�3uGŜA>�CA���l���~qM���%{�_LVa����߭�Ʌ�<&��e�L��U�RF���B� ��x4��8@�Or䧇If*��
G����0G�L�n�-"lۀ,Cޚ�Ě��r�zj4����^w���"2�/�s���%);Xs�o�]V��E��̹&NK����0��+u3� /�NF��Db���ܬ}��N���S̓!�R�4s�IC�2��
k/j�\oX�J� ��٢y~���ުb<#?��}뢓��n&|� ����Ks�Fc:�M�n��t��:�	�A���>�WV��`�� �:�8��-~��`$Jh�g�5i~)="gү�J���)�}�KFJ����/�[�h���*̍0���@�l�M5}N�H0�M�k���o�.{�L�-	����X��>S��� �*kr_�{���Ig��.}-�>O6�O`~�A�(6y��qf-KR���ϊA�bhduE�r�0�����L�(�G� cHI�U�g��|k-	!����ے����K%��4�l�-z�W��*k<�.��o���7�_RP�Ѿ�ۜq�h���8%8��xy�}�a����b)3���W��8%��x���%I~䏂�����-/^�
�DF�o�����]����w�e�i�0��BL�Ҁ�Wֱvڸz���j�4!-+���J�M���'q����GP�E��=l`�Ɣi�t�BKЖb�ޝWlt������6�y���h���a<r匷Og���eU<=K�#e�mɘ��:@��w�#��2=Oxb���h�e���kq%�2_�7ҪV�`E�Z͉�vbi���ze+D�4WekƗ/�����u}}R�����~�ά��9��Ʉ�z�"��z*+�P�����'�bP�f���R`�
H��쐄��a�4+���=��^�Q���Nz���𬩣1��Dٿ%�H��ަ����4&����Jn�e�	�3* t[E��،,�����)����1�nz�p�h5��-�ޤd�xOl�fՉ1b��|)%�4�5�F�\ݧ�ץ���W�)8T���2�I�G���f���7�4wW[>��[�I�ڹF��%?���B�嚇�����??M
}��q$>&�W�p��G ��A!o����{;��q���1�>�f����B�]=���o����4n|a�y����xA{̞yDt6�=�S�%G�v2U_��xo��$�q�����2i��zN"�)���Ci��o� ��l_�9�3��az>V�s}��8��ӝ�ө��i	1�f�a�6����p���E��ǈcU˄>I�B�u�E�ɬc���|+�8�c
wr_ך}��#ӓҫX�(jdV�X`Km����=ߛL!��=�_g���z��ʌV�H�]֗�l�Qu������[�Dג6�c����2�� :-�+�Kx��ipv��;��CV��X{�ѹ�m�<�Q�(gf���Ś���1��(C��|u�O��>������4%�lLz]|LO�z5-�&��R�d6��^�h�ݾ�V<�� 眇C�����Q���뢶���a��ސ�jx6f;��J�W��FT�	[q�GPb����	|��^�����i�)n�eNZ-V��.��	��d뭝�9l�����������R�m9�4@D=;��$!7���r^F��L�s���ԅ^,�<�)��)2E��Z0<��p�U��X����ɵ��Q����&,�N��C��vwv��`���Pq��������C	�ּ����v��s1u�(���bA�7y��3ec�9�d5�gb=ӏ�5F+���_�S�)y��7�='�t�9�r�v���&z�����	�(��;��s��w��p�/;J���O�ӝ.-�ZEy�S���[�q�@W
�5�4 $�E�9�ճ��K@��ҎwPʸN㑄��-{�����\&~x���\m$n�vԡ�]9�Ü��s���D��ވ�
GZ ��	E��_�&� �Yyi�����S",������prK Eg�� �������@L
�mҴ�MK����2<��S�F[	����6���'��^��F�C�y����ߢ�a���w鍼��+0L#ލ�)���}}�ڭ!�����oA��[Փ�d��{�ՒH|&(	|�VU�P��,�Sw�]��g��:7y�C���V��vƍj���is�u\P�����<�w66�G]��fi�Pn�@]"D����j��H�J���y�-=J�����啨�������5����;� ���T[{V�Z�1�.��R\�����t���Viؼ?j4�F�
��a��"+�Ѽ�/�����ePU.�l4SJ�LٟsS[,������B�?p/9Y��v�
�=Aָ]FC$Z�6�F+6���_��J��s���@�l�!:�󤿌qFrr��=>l�Q��W,	�d#wa����歃���,��N4�4���	�XJW%��P��|Rá*������#��R���?UB�?���rw(+��ԡɑr�6���XYkhK���P<L7^�i9�f�J_p����+S�c����a��M�LE�ي6O%OK�_h��
�f�-wO���� u7��r�
,�+���sO[�	og�ͫ�aL��ɯ����G{��r�7����7q"0�,j�-�VhP�i���3~�C�2ƪ�{�ApYI����V���HFT~5�
���9n2���/k�VT�իH�kpy�Nb�Z����X��ߘ�L�;,�0��<%��b��"W�:�>�C�x�6����d$�,����;F�Y��U ���� ^�9���v#�1���e�	^t�c�+�mzZ�5�r��qƼ����2CB�)^H�d)%���Bϻ;�m���|��]w�z��s���M+j��m}�ƫ���YLs���}FU���YL?�4g���m�/�D'Ҋ�:4�)EP����zܳ%I
��7�X�n�> ;*�q��Q;��;*VpŤ]�y����k�1��� ���`A�ˠC.7��ťT��iC���G�bTҮ�+��d��D�oZL���@əwE$#řP�)N�:k��4Vk����/�y������p[|Rd�ږ^�^����fʷ��/n��i��g�^툫��Z\�au�p?��9�9Dd_��H�S����.	��x�Xܻ��<9��2���E��d<��n$W!��u�W�AH~�[�X���7��=T��r( 1h���~6�ٽ����Wv��qޚW	�6p�7H����,&�N �9��|���f��=G��`�@͕����k#�:�#�/Fp�<�?��mG���\��s�S4�� �'}�1̥�x���pJ��sG� ��2?GY,�?!�&��Sp�̞�<���z#��-�
&�4b���'K9G�ͻ�����aC�3���)۞�r�i]8w^$�hgU��h���n�h�]M���"�*j�dyw��z{]�1A�e�%n���X �Ģ����))�+����������B�l��7�0�'���7"Ț���08�q}�����YS
Y��Xo.K奴F����ua9I!��oqR:kl�����ɲm\���oƕG;�K�>��
eH!}p��	v�8J��
]e�=�V�gL��z~+�������Aj�A͂�@vt-H���߾
�g�1-sU��E6g����0�֙gq��� ����=�rfcƧO�4�,�M� �1U~O�B��b��]�h5
%���{7=&��)��஻�=A��7���.ˬM�q�щ��*Y<D_Դ�k�aF��lwʟR[�K��q����C�6����BIZ����b��+�0;}2�53���m��w#B�|/c�S��j�f;XxH358��bR����.I����=����@�s��h~-��˒j�*"-��L�K\*zbћ���@�v���W\�Yh�(��J$
@��1jx�P�2TA�8B����1p+�0�����Ł5)�R5���AL�h��+�n�N��P-XM0'�X@�=��K���۽�~���H��1y_B#c�<�6tݳU��~����㰞�ʖ�>����>ƓQ�[�ӷ �V��h�-&ݷK8�D��!��4�!p�V>l,�-s������ꃭxz9��#;G�i$=ODժxPwP@$�I��J9fT�����ol�3T�`�[O�9��	t�!Rתg�4�d���T�,&��h`�W_=����'��^��w�g�VV�2�Ø$%z��(�Z��!9y�SK�=�|�%�x��8C}p=è]v��"5�^E�Ζ>h>Q��>�����I>��w-Z�q\�i�D�\G�भ<�6�5e�;�d�����å��6ܤx��ݒ۷Ѥ�.�I�0��g@q���7v���q�S��~xs6���l��H�ma�rk:�}Ϡ����mNU����˪y�# E*�N� ��¶�:<H��k��/��*/a�J�YXI5�`؊�6j{��N���a)�{&7!���d?�M6�f0tk�)ÎF�����C=�2G���x��t`����<x5��<�$ל�iжt׀�<�Z�?0�����o-��"��:�?���CD'��"2�G��hc��-����I;.�p�vR�Kc�x��g��Zx�-�� �9��6���z ĥ��r Pnծ�ݲs ��	��f �� ��#��c�Z�Br�v#b ��X"��5bJ)�or�j�AC�@�:�x��(A�ց4��\a]9���.Ã'McP����@Q���熍�|,����)�ɱ�D��9j֐���&'n�Iy�B?�\e�c���LM���������H*�*D�|\��<)��8é�mY�[ȼ��Q�?�1�%���������Mc�^�]�g��(��nt���4rRt\I_�Hu����;I���p��˿�r�Ypy�p?x}3����.���ꌙ�_G�U
^�ަ�ѝ ����p�	 6�QlO�ٷ�TeG��j-��p���`u�7��cJ�F�n��c��s�J��(P��Egd	̽B��6�z0������=�T���#2~I�My֮K�/�r�g�X��j�)#��34�3�i^�yy�<���F_�-@vܯJ�������p�.͍ݠ;���5,nÇ�HoI�OMY�a,l���{�R���{�\�����	uɋVϙ� �:Yn(4�ܲ4+6�5��[(�^�gߩ. 2-���	�6++k�G��d��	����K�ݜ�[,rɳp#�>��o$r����`ۜ��x��p�s�Cs�q%�������9���QFz�?6����{q�{9�������T~��ƍz�T�F%���Ǘ�
̶!MY�&Y�2��6�MQ�&��۝��-�����V1?�� b�ʴ&���'