��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��I�ɖw����$�OkA����.�⍁�cWg�J���>�eI
/��%��G�~�g&ØtW����t⿞.��� ˙!�q���Ch;�IF�N.��.I�u9*����㱽�q����6�c(*;q^XՉ�n@F�FM�Y9Ȩ���u��:����K�qUFArF���B�Rz>�n��~3Q��=���i�47��e�)w�YI{�ӝ����M�A1�F%t�U'�}�P�*m �!���<�� �*V�Uݮ ZP�S�dv��{�5����e���M�I�&u�7,�1��44l�}:�F�T���7�{Ԛiÿr�pm~=	ne��Xs���������X��w�KV��S�La��8���)��l=�*�Vʲ����R=-K<�҆�� m��>N����
iv+�є�L M��:�-�.D�'y���R(��0�|^y珢��D�ł~9Kr��ZN��!�\����n�P�e�ݕ��Jn˲|���7�37!v��B��]���ajN�Ŵ�e�k`ji�I}����'l:�6����/�s@�C;�2�э�g 7i��"�a��I�@$��	B*y">Ǹf@�y�TF�p�$�͝�ϝj:���@��{g~�^P���p��Y��q�4b��Rj�ͻē�Lj���)��$&+��89�pDF������J~�lc�~�t���G��{��*���d����!���)z�ɚ����*��s��G3㇖ے����J&aO��_p/�]P1��.[����4����4�C9�zo$T=����l��oܔp�v�'1LQ)N,H0��F��,�b|�U<�����&�v3��ĐE�ܧu��F{�\�1�: w���ͨ��������/, ��[:��RE��mgX������;�ȣw2FωJ:ց�����z.���Rт�>�tNq�e�.ۥ�ǈ����/q��>�m�f��C��e%�Ώ����:�[h���CN����|ZjTo<6�ZL�%2�� ��F��.���2.��g�%ޤy��F�;�4�g��QF��P��t�)?�c��r�=ha%������F�B-��/��%-�&U���܊``�+!ƚFϮ�R��1s��F���6�rA�R<��fɁQw�Bb@vOa�/==i��K�G�4)��FҖAoEL1	�+�I�|�U]�U�wͳ����P��J�8	�v�.F�p�����Q����
f@D{u�4Y�L�{�����C�Lc����o2�}�h6_$�}��?�iy�$rT����Yh���֛�ȉj5�(Ǻdg.O�� ��y��޻����9�`4�w���B��Z�� �@���_�$�3avW����M,(��n��~P.5��Χ�;�ϧ�U>��K��]�KS��0rd��#�+�n=����T�?������V�b���X8��W�q���Z�0��'�K|�Q\4ͮ�>��sP-�R&�J�=���\��xS���_d�숇u�)�H�x���qai��x��B�w�xcI�y�݅�W�um���	�.5���ǐg��E4��j4#�_��f��[�7ZK�萠������]|b#Ke��yW�M�ix��ƃjrk:?ң���p��2b@Aު���-�_��THM^,��!��~կ����V�) .%���.9Z�䌆:�,��4����9~�����'��؈�G�T�_�ڳ�0�_��=���3ED��!��ir�[�+:KM@�""�ɴOKǧ����j�ɓ�"uR�"pr��Դ���[ܙ��9%�^7Qa��S��@��i�#��-W�w�ZKXU`�)�B	K/����:�a��,��ؼI$~с��|O���:�@��}_�W�

U�X���Z������q�;R2���;$�WF���۝F��� `�+�eڽI�������K��E��~F;���eS$��"ƴHЄ�m^ξ��:_̩������C@���Z�/��9���y��a5r���$B��OA݉�2�rOs"nS���,��Lҝ{_R�{�0mA32Ih���ֲa'i�ZT����;qI��x�xކ&ܵTh�sZ2��<F����(ݍ�0�I̯�{@\F�v�2�^B���+�=�*�<��js�c6+�(�嚂�z��]K-�y���$Z�mv�:�\�p'q`*G��8�0���ػ�>i�滙!����NB־��*�	�A�̠-��E���j�����+8�u�}�HH �}i �]̰��>�M������qk�l�[�&E�{�ӵIB�F�?Y������:���R�=��fp&zf��PS��)}ix��c�F;���=��X�7�t����ɽY�ѹ���Cy)Mrx���'z�udD��z�u曨�=�ǭ|l����)} ��,��
�������˺O�$��6�����K��˃$(G~Y�`&-���|�s~:Im���޸�g�Хd��H�@�U�:.��L\����
��y�>ˮ�FPj�6��1��mЈ?\���a3j��^N�Eٚ`J��q��Vb���#lA��������u��[1����� ^�o��[D�!��5�uad��:=��.���]e[o"�]�w�	�%��?�[ܳ��K��!!��zlF�W7�v�Z�jn]9M�7���xa.��I��~lH0U�t��嗹��u�2���ڣY)I�DEG{ѕ�rw��YRO��d���@� ��൮e!���N��ٳi�@���.O�i��D�Y!�-6�:�Wkz���Y�4C^��v�.g1�)�?u�	H+ޅ'�r����?j�Dp^�D�5������^h���NT*��Z��0L������=�OK�oN�)���k�����GU��X5I�3�(g;�|�����>�`� �Uz��F���3���M^�!aR�gJ��t��U��,�����	�uԫ�֦�@̘�\����B)*uCP5D<��g�`�@V";=���!9�T�H�����C�'R�I)�V������j��X	۴�^�b�"��AO�4!:�qgΆ��5�ɬu��!_H[hOǅ�JLV�"#�� �F�Nԩ���폲���/k���@�6�x�ڸ����3�`�f��3ڤсB�&R(Gdk�h����5�'\�};B^Y���w��/f�h�W=e��P98�7����`�O�<Ww�x(����n�)�y���^�?S}��k5����p��R�i�3��)-o��cl�ba,<b	GX�*+K��)�q�X��zǉ��}����
�@�W_΢s�@)�HX�����q1���^������ CD�eu��T�O(�KO���SȬ�'��`D��7��{�rR�L��,�o���+��ZZՎ�J6Ỳ�<��,-]P�\�.-6]��b�@�o�3��j�p��/����bެ�x|�QBp_�!20�By�Ы��x�vZ�/5ƠK,tl*1&�U�ԫ$S{��h紳����/J-�M�#ll�)�\]���  Oצ2~��p.� ��f{�*T���\!M��:c{P�	� �r%DX����=�~��������ݏ��d^��ڄ�C��ؓ@�I��Q��3�9�x��<�>Ū2��˘��m:"_C/�[��뿥 �����}SV���-����bb�,m������6�R�A���m���`�������:�F/(�qA���ޡ=��т���L[~�)G�f)��Mݳ<,��<�Vrə���zp�����Ŝ�t��v�M�i�q�SRQ�^���!,��o{���@_�����@��c��7c�}�q��
��Ϳ�N�