��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��)sZtYzѦ�#����������^{���f����@,�B���ul@k�"T�z-��0��{�oQU�<cM i��CV��Ǣ���j*��>3���B��1����ݿGi�b�2g��8��H�2m��@�}
�G%�p���.�x�T$X�v
��;�b$C����f$����D�j����+���DM�#��k/��|�S��p�k�ҘMw�����t���3��	�ΆLww���LG�\��*B/qR�n�d�"O��
���<�[�ٮ<��?^�+�#�����\`2Y�Ϗ�cR�W�G���	@oU�z%�� �˗�#�fŪx��>��1=��&��mErc��ϿY>g#d����WQ��Q��h�.�8� {J��=}�17=E-�挴ە&0�3HFq���F�W]E:ń�{�B:�(��=Y��َ�o5qxE�~�4 %te���s�6cܮu_�b+�K�s�_H��м����-�]�Ô9s���f�Y�5@�(�:Fl���t�����"���s,*�D|�ޝ�'/J���v5�������n���4��>� W����� ��驣�֢�7]�DÚ�\�y-DӢr�X��5����}'�E3c�j��6�۫�����0D>��Tf�G3�>�~�0e� ��d'ɔl�GP�j0d�S�T@|�;�'���t�C����K�j������E��n1�$b9��z��!��o��1V��%��xh�Xy�����B"�u����hk-)���7�b�ψ�V�*�㿓M�}0K���.��"����6�4�yjᔌ �a�o��������6�1s���S��.��j9��;�;��|K��Z�n�>���^�T>�6�b���W��J����͆6}��;�"����W[��i<�_gP+Q���m���+|�G�G{��%7XF��y�QL�u����,�+�_f�4����9�.W�-��DFW�tڛv~_1��0r5�[�V��9���K�H����4���Y"d���s�,�ڣ��}�_��<1#e쁛�̍c~���y&�ꮀ��$j[��G�-lc���ǲ����?F�	@8���C���l�;�d\�V�hq�_sg�>&��4�n؎b������s���d&�e�)�^��3O%>I`^J�f�0�m��i^�¼�w�f�=�b�R�^��d�Ҏ�n�5f��$�ܞ���4S�&'����&�ra����zD"�I�J+�%�	oz�M��rM\G�(������<.3�{�l��Lݐ�&-���\j�F��U��0�%���{��-�K�� ⲵ2���6���:�~��8�n	&�BH��ah-��kx׈M�'�W�
qj����LK�]�`���@�)�d^��� N}�t5�B
�:�8��J��x1�����c�W�2�tի��x�.	)�A�Yh̊�9�B��=qY�o��s,��F$5�M�iԭr�ٵ����W� �n ��IQe��"~��L�<Ծ�}D�[�̻P�|
9��%?��$�Ѥ���G&|��}o7��__z����ޙC�K�U@�L�,e����T<��{��Cr="�����}�ZSB�鷺r�K���C�f��~���WP�j空����d����y�K������U��AP�Ff������	��P%������&��ƋqQߋ��yv:��I�*��$���`��-B����Y�J���B_(-R�;4�W�\�|b4>�r4/����;<?7c]��&n�iu �)�CޯoZ��j~���b���߷<�@�u|D�2 /Bw���:�yՖRI�I���Q���JB��vre�Gx��wj��9_;���i�9hBZ�}Ҽ#3<��;�N&Z��P���ʃ�D���YaH@����`�J*���)�K����%Z9�!�iBJ�x8��6�(�w�v�yﴸ~T��pH��W6R���7W�ʵ�PO�)��-5�kFg���#�	.=,���taT��D�ZY���u��l����ҜS�����zIy3��og
�!NӅ��j!s%��dM���`S���j���\ikw�sh���ҩ"��Ag
J�::-nWJ �q�߉���ɒaQ�A6��SR�j��K�^�B-�7�i��r�!$�&BT{e���=2s��q�;+���`�@4�t�9�����������2�T�UAiDՙ([��=+���G����H�.dYͳ��-RҮ!�}N���R45�s�p%��74���L���=)wP�ʭ�v�]t��g�Cl�Ei3�­�-��|VЃ�ʠ���^�&+���1��/����V��j3ctV����Zw��z��zD��h2�u�����wB�Ww:���j�jj�f���~tdu�h�wX��u��Hj���I�����P�h�ɑ�S� �:�)�叫������ �,jf�I�����ZX��y��%^ 3���[�s�b0|ڹZ����̕ʐ�.���V��Ȉ^r�Y/<l�W���`>���H����dtc�P�Txc���}�D'KF�/`�}��I�-�	�M3��ۨ4�b򨎹]Ms9�8�Z�n�j��ϙ@A��/j��f�/�kX��a��<T �d8���t�|�_��N���7�&\m�D�q����!���RxV�$?\{' G���F��-d	T1��P8D�f��	��K6.�SV���|y�����$��R�	�|��ni�M�Gv,�p���?��џ���ʄ����?J�g@�t������CI���M�:�M��e��� �L�=����w�	�X�����(�3|��[��գ���X�<�"}��#h�g�Jg����="	�@e%������M��=a�S�.S������� �]�,7���G���{�Z{uc�!+���4LpagG�L�m��w*���T�%�A��£u��>�5� 'Y���-̓�� Ӗc�t�Ä6_H>�:gW�l����V�g�Z��^v9
\�i����j�����X������E �(o��c0!��Z�<r�	��(OC�x��d鏶�R���=����9eC����O���9�f�J��-?��^S��,?���"������(Q��谝������X|�|�	�%W	D�N$�Sj�ӧw���)��hWΧ��0�,&�Ź��e#a�F�]Or�5����ۢ�$�o��9���kR(��Y�����7�)��o̐4������_q�o��INE�	t)��Km�f-�C�{���`^'��!�;�MQ r����$���3Yσ!��Z ,�j���8[!f��+��8�0.cz�Dҹ5�F}�o?P
��ӑ��E��������O�p��<�Ul)!غ��K>�%��6h���j��|���7�au4:��^:ӛ��՟s*#�������s�+F��P�o�6|eg���m��}��_ƶ�$FCƣ�(����Tߪд��J/��h[�ޚ=��rZ�{t�ޅ��3����ƛ��F
�0K�3��BЄJ��Mߞ���h�xulFSU�!�~���G�%77�����xN��j^�9H� ��_E�C]��ov��w���r���mLuĤdf]
_s�}��"�E��y_�&ԡ�� fcue��<�m"ɓ��8��a�0�����G�W���:sQ�u�������Ar4�)4Rb�_��n�