��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�fL���2��C�W�7M�̰Gt�6�����Ŝ`x&P,�"�ABha�ǁv����Y�?J���~���} �]�	��x�9���|h��*v�!�H�/S�l�����
�MTW��'==5b������z]���-���t�H��A��nI��_�����T6�Mv�X	[$��G�M�_��ܗA��?�4Q��F�h��Ō�c�dEt9�`�?xG�^�S�E[A
߻a�����C��+ۙ��lǅn.�.���
It�rƛv���c�{�u�?�[�XY��O�}rC]qE85��'$O&����M�J������A8�Z0��Kf�6Hd�J����s\%����� �,xnp��o'�6Cԇ�n��L��2b{8�����K��+�q�
�ͷ�<]%�<<X$�8)��\�`�A�l���+Z�yG&1iC��M�u�#�ƫemia^�Tb����#�d��2�L�in��K��zgL/�np,
��;�G6�MO�"΃�ُ� �lh�́�-��bNш�&����#��p�bdP��k���m��ΝE:F�6ލ`���tx�P��>�p���/`+��IOuJ�S��[�mQ+i�܎6��� �ѷ��޿�����Jq���������t�K[��4���f���Wd���G8*[`��PM8X�����M��K�'q�``���.�u�#C�1�s������pDpE����Ίq�zPhK$7�	�A.*@�\XM��~?4��C�3wVN[��l������4�`��`得���&F�B#�	�sY(UY��f���݄`��~�c��ٷA�7aʁ>ޠ�0|qcI�f���s@V�sCY6�Re4aX�2�����
��p��n��+Nc�dA�g��[��a�߉��7V��Qnb@� &8�H���&���$䯚^�W��\O�-k���k4`�5�Ǧ�3 f��C>:,�ND�A��<����*�������X�|��8��~'��������:���K��%O�[K��j�����,����P�q�L�	|�P�n�!��؍��6[�ï>����?2s8Z[y�8�����5������VR��Rm��KVL�M:֒n�i�5�U�M�p�Cd}��k��pH
TP�1�Lx�Lf�1q��i�D�w�	/<����9)�4l�o���} ��䑁ɓ�<>t��G0�~���t�@�|6sc���-���;H���� "O�󈭃�-4�C�a���2~�e�7�Ķj�6#
X�ɣb�Ke���;�a�3���p1��{ ���,��T�b��W��_K���R�� ^{%���VD���5��&�)�)��l���vb'#��u_=��~N*�5����@�lLycpb�� 1�!M=����T]�ޤ�&�wY_,.�
l_�y�$�Gl�סX�&Y4�D��,�NE�Wȷ��0^Vt������T���_[������RL.U���C�&èN�&ka�0�Xw���{�7��z��%�L��@��Y0{�����#ˉ�ç�FK����M�0Z�b�``��F@0� �@V�j�l ?�a��P����m4@��Q�)e'� �Z��x�Rj�C�����X
�_yG�5 7�m�M�'��N,�ħlhVE���㮥�1&�VF������J�j��o9<R���q��q�UH�|_pt�I�=���p ���ӭ �f�,�f2����L%z���D�ds�ߊf���;���<����WL��:Aˍ��^���$Vc���i::f<F������~���&wƌP�^H���0:F������cy��a�/~aqP�A����&߸Vܮ� ��C�	!���)�����W"$)�Q&�mqވ��7`��Rϧ���$��M�gɣ�]���e`ȟ��).���y���A���i��x�lT9tL�6y��G��i�.��k�������6������l�5�����S��wMQ�QԤo����*�e)�M�����o91��]h�|��Oj�00r��[�	���R�2v�d�(C*>�>�<����E��d���X�dA�>FtΩ��Ĩ�I���#->��!�w�݁�p�f�avv	��aA"�~��Ro��kV�`l�#(�����3"���>v-�ՒK4�ˌS�Y�;�fuH]O
_��!�aV�?�-�����6p؋z�ŉ�4�4��\���t�?���A/���o���z���b�N���S��z��܌��î�AA�S48�Á��2Rռ���@���3�?��!.��X�)1'���\�K�c�r�W�T[3�=&b�Qje_dN>6l��������יM�+1����$�2!*�Ь�`��I�K���2�l�VOb�Jf��ۜ�T�Eer�$%ƪ��jAjgg���zп�����D�������,[��/G��ӷ�Y?�}�J��DB�_d'�|�
��D��`�x}@:�FV�A�H}@j���@DYU@�K����۶X��N	��<�bd���v�w�O�U�]�%8��H_|bw�c����q`&|�BZ!�>���,�{D��{<�T�*�t��7���C&#W9�g��*/�����w]6v㟝�aPh�T���ϫ�$JAz�]�A*��p��(v���T�����s��ܧ�A��e�U����'�,@A�gk��y�it�����U��Xu����mQrAV�ȸ[�}�����.��K�K2����Ħ�e���h5���hR�F���J���4�J�ď�{\¾��*�l#3�]w�K�\�:0l�wz�@�lJ���_o�V�Q�s,������*A���l�eז&���d���`���u�"j*m�����m�&�����l�<�ȉy�ݍl!jH�����[������l���ͧb��|uK��P�����=N�b�lֳ	Yas�nX�C��9�J�����6 -�إv���^�������~��������o��j��oT0��K��I#�ۡ��m�g����ke�p���T��{����hx�u -ͨ������l�o�X��� �GK�@�Q�5�)B����t�S��˚8�>t������nB��?�qq��F(����:NC���!oE����,��u.Ӏ�)ۄ;o6��2�$�S��|���Z�:�v�1�A)���O����B2]?-�WUyHW��2å3���y�։�<Q�:�F����э�C'��� �"����ԃ��y�Y� U���[�Z���3����s}�/�	!�]ʍ*׆��8�K���0-�mn,�k=sl\���%a �z5^��"�����߃����´��<f�F��^����,�cE�FŪcy���#ڈ���	*�d㐭��j�=�w��ن�ƤI[ϸY=P�2|����G<�	Q�� W��Xw�'�Ӌv� 4�L�Ē����c^������Q��l#����'
�&I`%�G���ܝ�K�½󱯷���ǎ|��~#���Dj�9�8]�ڣs���c!\��Q-?xHk�#X�|��sJʣ�P�r�|Wm/�v��U�6��+ĕ3��z��.o������D9$'�M���\X�3t?��
]0��K6��ZBu�;,����4S�ꤓ؃�A���;����
B�aX �1�y8�JgM3e�����U���@e�
a�8H��o߾^�Nʺ�#�3����5��?���r���.�I�ژ�T^U�?d-U�Y��x���w��֛�A�Z����XC�ז̨<�pc3���j�t��uuf[���,��g}!J���CfC������,I~���a�S;]�xZ&��K>�o�	k搂(�ϱ[���O�uC�w��1%ŇЉUN���q�͛�	��ѥϻ��뻃�B�s����bL	؛��
Q��s�楻p�a�5i;��p�E`b���J<���^�?��"�M����gJ7��W��}��dʺ�_t�5�<k9��UL��_��@j47�ؙS�C�ȇ/b>�I��i�~�~��]�Y���	��`���b!᥉�>�3	�X�Bg��\Y��a��ơ��t��q��Ę_�Q냽;痕d�T�2|�nPڼY�r��y%�K�R"K�`�k��P��=>��E�D50���Z����n%�x}S�D{�rP.�ܞwD�PW��2�T��հ�)�^_�e��튃7b���/����o��=&�#6����Heb�a��iA~�Ð�T�h���@��/�O�e�k��_8P[� ����?���b
,c�`���J�-��X:��7�ԇ��KM,���2�T~�s=�4��C��*hc��y���$ 0[�# [���a���D�THQw�gA�ĺ��Gu*o��"��	��x��"ސ,�f�H�|��ʁY���Ԁ��
�m��_�kʲ�֛|Oj�0��]0���k�y�������z)՟%�-��M��Z�,�?/R!����9 ���0�ђg��V%f�T�s��sQ^�A����f����0"�5$�g>�o�2(ߧ���S���ȍ�1�m�cN�[�5��I�%���'������o:�X��l�\»��9��D���tV��_	P���^�v����zL�Z�6.���U�6�q��'��00s�<��v���gn�E�U��X�@Ri`>6w9I�/���7U�ۘ��=���N��OZ�Ar��%��֗N it�>��F��m"���2+��>;��c**�cD`�#��!x������z�<K��sN�>[�%+����k\9k�`�3��68��z�N�y�o���Ξ8�e�X��#΃=�-�����M��=
�T�j��.$�ƈ^��gs���>@����N��V���܌ҕ g���D�������ɿ�XC���_�����N��d�������\ej��!�{��|}Zp3}��W�֎�������:2�b�g_�I��F��ф˂�+��	J*�1S�J�/�Q�X����^�R�&�Ec9��.8 �0ì�Mwd�;Rq��KZ}��ۿU4-����3Y��YM��������ܞ`q�g��<[�	���c�Z�Q�P,Mi���>�'�ǣ��I��"��ypś�yi�����$	Ww����	����q�1�hIXE�C��Lm-��ӵ7�?qfK=�]��X�	c���C�a_Wނ���;D+�]�����ɇK�e���ڠ�g�u��eo���,h�)���F�}�'�|��Xs��s�M�8��	��pͶ<�5�^�]�}�$��%�\�+��P���X���|��?�DL}�ǽE�&<�-<#�d��E�lڠ�xP�]H�bFC9'U!�{���R@�������U8]��z�L)�E��
H9�j
6.���Ϥ�^yiH�O�Z0��?�|!}��kz9��/�����4�KOd�n��d3�m�FH�ǎ�=�\9�f�w���a9ǌ۽��)$F���y���a���z"��n'?���� ���22���o���Z�W�����;��
p2,��O$���K�+�n�2_;b��i��y�'	�H~u��_:���j!1;1�$��JY_�殳[�<��c�5�6���v�%��~׷�pKn�*i�������G7_�w�C��X�m#)-Z����P��(=�J�+H@Z��̩i�b�<z�'$��V!|�4��Y��Ǉ�2'�+�I���D��������6IS�ga���v��o��7}{ش1���dX_%��쳍TP��	���J(]��F�/����Ӡ�
�tRV��x��X�����uJ,�=�X��Г�,I��5��-��w��T������."M$7�l{��>�1��v���˜<U{*���H�g7�����y}S����NA\��wү��XA�����!`�2�X
�]�6V�j؜�QƸ��ض�
�Wff�U~}�T4����{��)0�urek���'jWpԌbR7#P�݀E�x�|���u�{�`���,ם��ɿ��6��9��Mw+-�G��5E�J+W#T������n���;oS���,�U1��j��_Z�F��)�4#6	Ŀ�ȏm��W�P*p���gѱ~{��4�	O��n�v��a�]"QԚ�fdԒ��mL���I���+v�cI��T�^[諁�i��#e	�� @��3=����e�F�!�!fZ����]"
n����$��_$��4���3}�g4M��x�8��~6C䥝S��[�h|�ҧݜ��d�k��J�W�%�*]�UE����z!Aqt>`�ed�/�)gК}�+�!��$���ĝWN����K�b6ĩ�z�z�\�=�[�q��|u�;Q,J�Z��+�}SҘF��l|������{�0(�E����ULZ��HA��6�	�)�L������!���`}���,t�&��":ۧ�
V�iE��W���D��1K���D�'A��8h۳�
<��
%�����ܭ�
a��a�<��E�Q@�D�2W]���;�wϬVc��ɰ��C�ݭ5�?����'�q���>A�8�$������s�D3��Yy��h^�#�X2(,�D�j1 a�Ʈ!7f������om��O�˜�V�!� ��oJ�F�&Y���®���ʏZ�T�L�8�IW�M�g!Ԓ�U"]7$�yŨ�j3=�!��4�C���.�Μl�u,1���s�GA O%�xQ�����J�)\D�����|<?_m��>��4�8rP���N[nm�=�<~�.ǼR]����ef�Չo	�\{�i��P�E�fF��[^��6��Z��\�m z��ZJ����b�ræ���uEHI��ѤP�TDR�K����Z��;��Օ������P��%U�Q�Рf��p���?�萯�1��d����l����tq�DUf\�6G�m�h�%��[����'�Ǆ�z���1
���vG�����:o0�;�x%2mˠE��'U��Ƶ���q�qtC�\He���G�+^�V��F]����s-؄��|�7�$*sL�x���"�����������	�+�_9�;�|�2#�����-`>X����)�<�ć�������r��]��\��9�����щ*�-���-�E��`1��P�Em�Kp��#�9���Y��k)(8�߸�7�`Ӑ/r���:C���q����;��v��H��9�!(�-�w�����`x���1��#dO��Zo]S5�:�`��)[ �]S��������=��
ip��-×�}��H�y�����F>
�0	� �Al�P]���!��;��q���m��9���S�l@p�q���7І��@��Q�ʧxҩ��b�u�rO}ĸ(��N�����ka��,l��N��/�+*p'{e�5�v|��!�X�R��涡(�{�hT�a�EO� ����C�1�œ��2� tg�CI����`t�]��b��]z�����ngj��_�٦�D#�@8�i��a� n��=��՘�Y�[I!����yf�?��~���&��n0���[=���=��=rE0���?D>���.�|�5|��L�:���˔��dv����%}8��)��/�J�[���g$�Ź] n�c����ү
�\Q���r�r�R�6^�W�����ti*��\I+�?l�V���E��v�J�}�Wo��J�#D�1�M����9��U�e�(2;
��z��f����b��h|�qp����ӕ,a����3�K�֛�G+�߉���I�:�[${T��X;d?f�(����O�&Q�4�뿍��2I��ՙ����- �A|K�S��xm��_�@�?��%���p����t`8�Y�uOok7�{-)���*=�(o��U?�M%��$�O/	"���%��XW��l+���f�'7�B�I��R����y$�ȸ)�B|�j~%0l�we{n�B��tņ>!}���jK��R��?���tఇTi�C�e�x���h���up���fe{W��b?����_ق�=�����ؒ��A�ц��kΣ;WЬ���N�}ѿ�ϝ�U-e��C��TX��ȩ��g�%���;���#�]G\�k��O���
�`�5�J^r��g����R��iM49��r�����7Ƣ]�Ԝ+�f9�u���4U���՘�����i�J�i���i�)�O:���&�ˮ�֎�����8�ˀ��>�H>��jӔi���e6%�_*P�r@�f
M�п�EM9������X�pA"��a�(O�r}q�=w4(���	~}���9����������U��Q-y��-̆�ș ��VvA�G`���|.��~�
f)�Q}Pa�n�������OP>B"� ���A�c��0��`����3'BW���b���aVF4�~K\��u���1��H��n��@�+��r !·�6X�8�/�w����;�|��f�����5*W��/��)y�w>U���t6��ri��aPn��Г�\= ��ճ