��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]����'ԈO��J��m�:]����@�G�,ɛS�_e��zY bZ�el�2�s����^O.�����zi�z-�g�~�j �ZA��9��8B��t#d�IP�?=���/��E	���A�26��xM��v�wm��(��2&�*�|�ӁV����T����Uv'����+ɰ`a�a���{�?�����}��1mk�oy��[��2F�M���K�Y�(���;���=�qv��@2�=~�(�L�O�-FSq�3�~��9r��!w�Oô�MRR���0"v=�΢�,�hq/0��!�Z�d���%T��JL���@�O�׈*�:�E�O�Z��+z��=/E '�����je�g="1�P{����h�{���F����%Y%Bq�{U�����nw�F�5����:}%�
�#oOx�P��Mo^.��	�[]�f��������oQi�ހ U�\q�D~��C�d�A'�{�>��Y��0�y.�k�g'�s�>�d�Fbk<U��S�}�\s��rYl��=�,�䍈��;���fgh���h&��*��[����˪u�F�V]PpM�oǚC� �t�f�{#iQ��\����l#���u���6���L[CG��;��hAV��N��0��h��f�>)�1
�π�-�fpy�d%8����Vsפ�~wR<jp��o�dh�pD��c�;��\T�/z�?�Z��R۠f]�3W鄗d3�SԪ|Ϩ�J�]߸I-� ���se�\R�G��n��r�I�W��o0���[0�3̋ce~��@>j�f�D�WY쀙nz����ۏ.h���|��l�:�+�6�4�3gF��8�V�qt_�=���rJ`�|�LL��a����+�̆,�+��)���=��!޳�l�t9!-E� "�	�n�M��u��oq������;�nJ�ͦ��Ɂ4��lF�'$��^=+㣥�x�==�b�8�ǑZ�Ac��`�.�A#@Z�����x�.�}ARH��X��h.�f�5'��ޑ�$�R��H�T�7|IV�P�)d��8$�@7_�tuQ�F�s�5�<'�:�=1�9�SU�����Պtfk�����gX[�׬���hh��	�hB�}6�ɯ{5+l ؙE���>*��:�Cjq��ea��	�O�.�$��V����;.��Po�L�1��^[	�qUvm���D�뿢^�ɼt�:d=*�z�x砛�7p�5��F@�N�Ď�����9w��֦���ά��d:_�����m�²����L'�0���T��㏕��4"!���?�0(ܚ"x�Ő����=w6�V}!.��Eyvި��`�b!����B�	mX��^�ى��ͽ��I���"8DGd̊a>·������/;љW4�;�R̶�V�j�.D�q�A}�RW�.��?�9�4������ m�6���3�wb=��bAI'���:�M��wU���,�D ٭_QV������r͉.��AHӻ���?�`X�f��q��0�h�l��W�S�V�)��2��S�hB�
#�e�kwn����p^=���[
������j3�6�ez`4��?����j�"3���ၱ-a�]������A�XH��پˏh��P�5�D��7/8^�0J�����D��#�aO�M\�`>�%����}�K����l��h�ҍ��L��&�]+^�{�G�MHǭ�M�51*D���~���P&��	+L���"����Et���%�W��7�=��{�a���Pwߌ]1�M�up�Dw30z�>I���7���C�n�^���S9���}rL:���#���nuB�� B����2��i�$IҊm�$7���>5��x{gg%a�h����P��?(C����d	9Ğ��6��{f����T��(<��&%F̆%G6�c	��w5��_���r � �G�h9�X��l�]�h�J;ɵ�6��İ�&��3��v�*�*�	�RR����_�
��[���J�l�Z����I;�"�=��Z�S���3���r�FZ���o�kp��rJͤ�`��Z�@��J���;�|�����c��mH��3���$���7<t�A+�]�;L&4��ܒ,~��cŶu9"���5��BLS�Ń�^&�v#��E�:y��c����V0E~<��B�fM��b�B�~|�7�=���g����( H�� ��"i.@?\SI�B�w�wX��+�m#� >�_B�MU��aQ,ԍP���u�� O-��5�~4�f�X�u#`e��c��^�����:���y^g3G�7��qZ+S����?.��L읝��\j��+�C��a)���,kq�z�P���@A��Y�����n��j�V�t�l��1���Ǻ�+NV
��J�Rj���Grwຐ%U��|H�������X|��7�����ඨb��,;�ޗ/6iS�w)NnD,��O�i�h�-A����7s���$<y%�X�����(�D3��Q�rF�3zG������5(�wa�?���S�L�V��׷�N�H��ڂ�LZ�r}�����-�h�O�w/�U�̅+��I2�t��f�]���뷖sQ|��ٵ~���~�7Z֧qS:��b'B�sM.H2�VB��]����q��W����?���Ѱ���H�7}��K�qj9XVu����$����E�˟�hU�{��0�f[-	N���&�*9q#Ҝ���� ��:%N�g�/4�F;<)"z/���vn=Ջ����|��x�\�����.���,��jIIy�nqp��PLh���]⩷Po�J�$8�x���$���{ơ0�/���uN�d���W�=�FNZ����S���98I��$R��KtV�JIٯ�u����R��3LV"�n�)QKፄ�SĲ����7bz<�UJ�=��1�7�������iN�8�:3�	Š(���0���t�/��eLl_�N|��2p�;%e��;,�ڥLw�t&~�A>������<����@
�q���~/L�֩�����o+Sgy1�\?�&��:��
�����X�ai�[��W ��/ɛ_ϑ`Q���ߟ% �H��5\����c"1V��u�:>�#��;��j	�v�X)�>��ɦ%�s�+?�9�r�P�V�?-\�^N����'���ej֒����� p~+lrL��\P���F�C~Yj���!�^z[�w�����O�E��A�\^+m[|���Q^>D��&��.;����/r ���%��ۯ��y>7�8рG#H���TW� m^����	s�qx�oeL�ʻ�¸m�,����a5��~�Z����A]���o�!�q������NH��l^~�E�	��4W�A�髶e��}�2;[�ZJB`6�p�)lD�Ho�;�@���}'�hҸk�D�6�$d���v��3���F��������a�O��ʏ���B��E��p�Ǐ(l��3���ɵ�#���"�o_��ύ�L��Z�b��(;�|���p�kL�T�j�[��1d)X��Qޔ�i��p����u�iy~�HwU�R��P�=���"앪~���� ���|>��@R\-N3#�G7Z�H����A� PU�BSͽd'���X3E+a��}	�
�7�� 8O�,�����-�w����3���ϓ	�3Z���_N�����Ϭ����	�l�b?�ڜ,I��xgfd>��4?���Hʧ1�a�5�F��P�b��519�C�
��@��*Da<3"!�]]�$]���hĮz��6���S���gp�,n�"�"��-��A/��IW�=I��O�6~���tn��a<�u�[�6��  Sŵn�%��$�X.���r�p����~_f��=�&���{�G^�lw��Y�����_�9��~�����t�j���-��)�	ו�	�zޑ�s�ɱo�+�B�KWY�"����C%f�×S󕩓ۅXZԕ�.�Q!�ʼ3�7��E'��tS���4߮5c5�����u+�n��~v{�/y�x肁�����7�Rk%�ı�+�0P���k�MYOS���<4�$1E5 b_���J]��T���w���A��ze���y����;
��M���O]5��C�w5��b�9lZ��!8_�8�Zn
���0^6fd�aI\��� �yD��t�[��^^��'���_�d�O�2Í��� �� �C6��1`�x��K)�Yp0nrx�QK�aE�#�!+��Ѭq���sZ�-X���}�~�T�i}V��./V�Q��
(��R��m������oqO�	z��K	�]!P�Ӟ�s�ׄ3���>�K��Ϭ4؟�Y��d�%-9켌�A%��6�8��k��k��>�%�d�4I,Q��ΪrG bxm�%>��RwL�&�%������b� �U�V49�ē<aF�@O�)�?F\a���<GD���rm'���0@�7Ĉ�V�u\2kH`����"Ki�����Mg�R�s���2�*�	�4�������ˉ�D���@N��|�>|�
 Z��H_˘�o��0�K&�~NZuq(s�?���g�D��$Gs��3I��f��`����L9}�X� ���쓚Z[s�C��J����wmI->�� R�����NV�昃}��7��)%��V&�H&v��lw+��f=���t�;-U�?s?��"��M�4�h�O�%�(b�ێ�ri�J��r����S��/�Go�K�=�0�;��'���/��uWn�/��b�=Ku>��L.���#n����1Jm׏f��^�=��v�����z���M��+��^;~#�B/��
�h�J8��!�Ҩ��j\�d �.j�R{�=d�fz0t!ڸ��,}r��w�c���OE�3"��"�h����D�y5�0&�C��_��&Gݑr�AK9�0�^���H��1�n�Ɨ����q�����7��k����Q6���\r�W�屯��`��/*�vʘ�s���$����PL�q@�X�)ﵡ�����F(uw�ULu�y��#\��~��9�]�񥾆:�*�܎ר`��	�f����������we�FHqX�_�sެʏu7�)�Ԅ����Δ#�%Z�,ct7�@::����KW������m� ї��A�����#;	� S�?Y.��T#��E6��Tԙ6���a� ���-s���W��d<����Fp�H>$	���*����v��|]�XgK$��l�6�K�a�S�|1ڕ�ig�fw"ZW��bɺpKZ�Tl����%WI5��P�9�7YF;j�zW8zlb�bk2�N_>�lO�9��(�E �Y?.����(��h�S���]H�j����^�&�o��6Iv�)�t��$��ڦ>�_���N����f�Pր��@[~���sz�uU$ƝB�
{��]�ի.��j��l��U��L�\�c�|���|�'=	�e��O-��&�M+\Q���N��/��֩�j����j��yp�x��zQ�mS���k9'g�iU�B�8޲���L�la�G�l�J\�М���l�?@�&ɻ��м�J_�w8�hUipfW�p�F3�
���H:�	����^�%GTA��_,�Qߠ���,����YA�������la���œyM�tJŨ�0%�h�Ix��M���,��Ϯ�
�u�*f���=  �n�v��glyUӔ)�Dr�}��s4@��}�0���
�0�r���r�uզ�9M1t0��K�pC�����6!GB�a@j�����>��G��"�y[y�{7-�bc�U���o>A\�����E�3ѹh��Oo�xy|��+�Ǡ��Nw�R��|QRM<���%����<��� ׀
 ��K�;5SA�_�I�;C�����8�h/F����4����8vy%�2��|r��Dl��R���_�-^�2Ax���,@egă77����u=Ghؕ/�L%����x��v��Nq��18�Xn"!jE�Ϗhօ3i�&Bo�Z�\w߽wE(��ˉ��
v�+Ӷ���P2W)U��MndΊJs�V���[�^�%1��+����Qu`��aw���A�:=y�n򱸫M�gn��Db2:�ا���R�ڄ���n�|}�^!0�4�_fR�� �n��@)5u�����OŶ�1g����^w��O���4��5� T&%aL^�M��&bj�[��r�BFLIչ��x�:���+��oc��Ť���\�j��-(B�~F��T޴)g�J�9^��<���vؐDv(�I"%^��
E/ �F�Y�c��j�r8����Gu��,:�0�\t�����wm$d���<��̵� �&���1R��؋?����\��Ц��'T�Zh-�uH�7lp�@�"��WBw\Z�^��ƹ�%T�w��p#IZ݅�U���I  BǠE��j�~��k�	˛"m���c�W7�҉}ɳ  ��&7)�g��m^gŅ倖�`��n�f����H���:|�Q��1�1����{�d`���p+-���
n_��Kg�J��<>Ȁ[v�m�֧oV��[1a"Ha2�L&H���0��P�P2P^ -��d
���u_��!�ޤ�P�;��פ+�lvh(Z��-Ldr�[]�_:-ʈi�^(��7���`7�vE���d����Vh� ���/״Ť.m��Z�����g�%H���H�X+9��ӥ�����5�/Z|s?��3<�+���7�IC�!�XX]hv/o6�KB鱂��qӻJv�d�,�*/؅iO)���7ސ�� ���"�F�bj$��d��Boy��O%3��P�O�ñ~�5�@��d�8��VQ�2�Mno�Q{I�PK�	T����s?����� �&7}�ۙ����>z����jtڍK�]�����(����հ�SM��iJ؀8�ދ����b��q�C�M�7Fz-�S���f��@�o�n���
*���#��k,�⺛n���5�Zz��9�=�Y�B�6�Vˉ���D�uМ���͕b[�&��I�~Z��;(��E�KB�4R�i���+�8W�(���Q�֐P�;��}9����w	�{6�!޲�H�BM�n�K���2nHV���牲�"�z	9��f�~2��;ؾ�8+Q��66 ]?��ͬ�[�Q���(>erA|,�Y�r����d��,{� �l�E�.�C��g�g丼���Xft���s��:b%Ousls5�X*���%R��u��k�ki>9�@�O{��_-��^鿤�z�����#��8���1��d�R�q���1�$ߤ�Φq�?�������s2mi,���Ξ�N��']��i'��!��M��?�ޮ��і�U���3����#U����!�0�&tp#����/��`*����u�PY���%�0�9�x+�"m����$��Ή��b�.��l�g�� TB�b�gT[2턢�XD��V�* ��i���J_*��P8�G�Z�[
��u�v[npZ-�Z��p��������r�ٹ�!Iui>�3�e�@)�j�Nu�D���%z1ğH/�̚5`a옢�P�����ope�VX��!�k�J���.*1a�;m��'ȅ�����V)������x�5`�Ĳr؂ozT�C������N;�L���>������r��d&�G�q�-�䢧�l2�������|�F��[t����Ԛb��m�O�!gt�8#����v-I��ofu���RL0rqC�7�j���o�3d���L,�hw��Ղ"���zS�:�~M���/��<Ux|���=�[�I�*Ke�K�{.wR���W����Ҽ*�м�+�"���(B5i�(/�r酃N̴�^�l����,h�|�谙�ɸu��!����}奘 O�7~s_M؝�i�ۖ]��30�z�eD�쇠$u_�a)�-�gjooNd�g"%YV�-e�	�ֲ���m�ݣ�H�o�<���e˄|Pښ�'H�1�&�G6YyjN,C�®�˅NͶ�e�NN����oʋ�P�l�u��,�IBm*�.�e�O�}���]�A�^"p��Z�q2�tϤ3b�x9��5c�ؤ��N'��}�,�+���d`U�����#��J��x��鉂����������0ŧ����@�1���ʵ�����!�@0�?��"��/wJW�,�/�P�L��7��ӸU0j�\#|���~�q�Ǌ���Ы�4��!B}$��vm���4x6N���U�>�ʩ�}saت^]e�T"xd�2R6~U팍O�8e�t#o"����3R��da��:��=p���n��;t&gzY�����M�f�o�q��D�n��&�/ȵ�J��M?�	/�*��!��$ ��� @߀d郌Π�^�K�KNx�� Z��+�Uc�a�YkA���a��F���~����i�B� ���.�#���fW�D�������|k�騮:R²�����G��(	��&m���>q�?/�/Q�>OE��t��z�_���RL�CgA��Hs�aDVL��,��ͦa��l\4�n���:��`��p�9����Q�MW�/�A1�����|t�s0߱O:�'8��l�i@-�G�9T^ᙰ~�X��,+�,ݛ7��N(w�,��)آ����/�K%R��iGH"Ul�t�Q���v�/�*�*Z<K��|�,]����ģsl#"Jg�P�q�Nh<m0R(�����c(w.�=�d��������7m��^sy�е,�&f��K�=}'�z*n4�kЎ�Xm4")��H��'=E�^�~�ҵ�l 9�����Z^���G����ע��]��
�~�9�L
v���Wd�!�A�̸���j�Ѷ�aoG�X�f��8c��MT
FD�7|A��-��t���H�SaT��m� m�z��u֥���}2e~�O�j&��my�Ou��݂�g��~�RWB�2�m0�_e!�R���>���A��d���I
/g�r����0��,��Q1��Drxw��;�V�����&�^�9`u����e�9�w�!���2���i����u���b�of��v�ƩU���sˣ�i�وX���gO����<b~��eD��e��KC;y��P�L�3���ȣk��t������R�Ф�`&3$3(��]"v���ɏ o�KW�-��V�v�~7�a���`�g����˺�a����^�
~�LO 3���E����908��9�V���	��|>��TQw�Ï6f�64�������� �v�eKa���o_GM�U%���!�,)���bX�y&�J���R��˜ˢO�L��f�h\@v��aa��J[��u_gp���G}As�;g�0]�{!׺'�E�v�I�J����vW{2R�e5v��<3Cη�7a?�H���c�Y �75&ꍋ�a�����Q$b���Sv�Dz@��Oe#L��� `h��s-I�UZ�Ԣݞ�-��|� ����N
�D%�3�~6�{���4��Ey�-*��֓�Q4����w�T���rœB��֭�2��t֗2hһ�V��E&��Pf��ǋj�
C�m1����)�0�d�z\�l˜�[d��vӞ[�Oc��6h7s��^/�1���kp�'�|`������n�;�K6������ J�%�%Tɠ�eA��6�G	�/�����%���3�<��j��L���J&fm.?�����[)���e�`|�Ǘ��g�_
ܬgZ������ ��
f*�zυw����y�k�^�%�d��Y`�v�HP!I��?t�:,$�m�'���̕��ߵF���,ꁟg�T�=6��A�L<��:��+�9�3N��U����S�-���=��$�NU:nJ����S��5�E�ZӜ�*�2��q|JPH���z��Xȕ��?M�hG��|�WEf�|ǛS�;�#��e��En��'��Ś��t��37t� �i�$i7ߑ��Q��>	��^>%��8on��ד��!������q�O�,S+X�@۬��Y�x��$Y�����/�f�mf�{.0C��>�U9rV�.b�-Q� #���eț�t�S��hK�e�����?~k���{y_l#�ƾ��Dz���&<e b(� mӢp�#���}���AR�ܣ�y?ԥ�)U�;�w1ߑe�b0�ڄ�N�oSE�a����1b$G��+܁�AL���Ӊ�IhHi$
�$T9��U��g�#@o|��Qg�H�æ��Y��:p�(Q9uN�*�e6E�i�j�������g[�٦-c�;]�`���*�ͦ#�hNj9H*6�@k}�/����h������..r�s��+�d�e[�l��PP���W:�M��C��=��w��A�:c���J4��y�5|�:���6&�����:m�MZ���Pg��9ZA{���ɔv=o���Z8��%�^p���T���e����n(n�{ T�	x%G��C���!1Ok�ȋ���:�<+ѝ�钌n'q ;sŝ*��#)b��v�����}����p�<�@e��Lh8���$&t?��	��F�V�Q
l�7���0?���;6*�h٧���RL���{��r��ib`ߟ�Wޒu�Q�R��j��+$�X�M:��t��!AXOr���Yt@)�-��f�^�Uư�:&��:/�wXԞ��-��
��t��*�����\:z�A����������E]�A��2�b[~�He��3/x���̙L��Q�B�VD��$-�ט�?]�ĈzA�5���4�$jN�n�ew�)?)�/�h�g�c�71�9O��Eakl�E��G�������8l�۔]�;����1?��֜��v�y�&���!����5�[���AMD�t��+w��z�Ώ �2�J>̗>�Õ�7bJ���ˏ���Y?��[�+;v]ծ����~�@cN�����쀐���K�o�2�5$�.#�3x1׈���ۧ�]gfF�)&�.��ڔ���p�gQ}臹 (s	H_�Z�5C�Z�$k,��ᵒ� 0����E¯��<*rpі��`�#�T�_�Q_��0L�B�����BlF��v��ԗ��|�������!�6s�^T*���e���;�·f�}�u���.@;�,{H�m�H^�]-�M1���g�
!K0Rp����Kz��6����K�^8C���O�pX� eF����p�6";��$M��U�w�[�K\squ�zVs�d�v� c8���|1I��$��H#+L"��S������� %܀���lK֏F_�pJ
C�h���nr,�-/cut�nJ�_۾�
���Q��]]�Iu\8F�r���H�%x��k{��EHa'Ճ�ʡ?��ࡾ6mA�l�^���q�7P2|�x!I���K8�*��>��e"8�	0C���& �a�j�2¬����?>�]c�#��lF�ݱ�A$�S��O4�&}�ѫ2Wf~ߟ��.�
�:v����1Jd�+��;k�i���դ�L���Z��@��/\0������9g�aA�4"��t����*u0�=�h-��Cj�
=[�C�/`&���nʩ��YO�4�fܥ�U�1Ȟ����!����o�PS����r�����:��3��7������T%Z��.��tC[�<Ra\Fz�����`�9u�
0Y���{l����E[�M��;�$�	�ٖ���f	@4Z��ǥ�n�x�誎�k��#�Z�kE��qhU�{aC�-2�G��;ɥ�a�2i�#���R��oQi��|Qy��dZ�=�د��V�kk�Cٚ��ڍ`pp*���C�b3L$e�����"�a�E	
��H7�_��=�.Jx��f��z=��#F#4�(�Ľ���X��Q��7���<�<���f�|��Jq��bKHZN0��4�`�2I��*^�����]�9N!ioƛ�Żc�Y�@�0kl�	�>�@c8|���NU����A�����(�`��t*a?�M��Ĉ�xi��>,�����I�ߞ���.-�/5���Чk���x#ĖuZV��JEb`��	��%���Q8�) ���?7����G�w=�����&�O�y�;��c�ز,�c�ǵu�Z��v�Dk]��E2����6��2�n��y���8l�?0S��P��d�J#���M���g� ��2��M}�f8GƵ[@��Y�'gVf2渝4��I:��3H� Мg��g��a�P�RE��ւLd ����˝?���4��5!��>`�.�\�9���z�����Ќ��L+e%m'�t�@*XE)�=�x~o��:\Y��"U�/3�wΧ�{�ٜi[m�|����I�a�Z�]x�SE��,�Vq�������AU>�?��~J�XP^U���՛����"iv��l\�N[!��݊�발)d˲}m�Ɠ�I�fۭ����[����j��tl69
��ـdI�k�L���x<�V�,J]n����惤K!S��m��4"�������ߵ���7^��
o����.���$�	n^1F�sR���n��Zt�UV*`!��,	%�A�*�:��/5B�ڢ�����C�A}�n��P�>mV�v坰L�C��x�I���������EH� ���D����o�G��D����%s!2�*6���'Ѡi��>�@ه��d�8������c�ϴ��[Zb�8�YR^V3�ٖ�u䷒��$��m����ym�5�QC��v%��R��W��U���#�jZmD4~؆WeAy6���gD��[�'����_\rJL��d�H�}{f�Ty'!T����7��f�Q�7`P �xmЅW� ��o;��*I.�H�x�4M����A>
�z���K��W@��+�VMG�����`%��7b�r��M��QV;�7�`@^Q>w�8�r)OAj'.��\�>Hb��o.`ui�q13JF�m5�SBnHC���	j��J'��k�Txy<�vS:[lf2�s*$чsQ�AR�?蹮y����1��9&���Q����{A��� 2t`��� sȸ*����}2��dE.�k�w�Pw.I�4��_�Lc�h���DP,�0(#�k�ί�~ǣ9��Ÿ�`�c��y]�c�S	7�xLxr^�6�>���i7�g	�Yr&��pd�{1�X
]�C��d_������t��0XN�1x`+$��ƀ�����v`���U���*����I`����-������[Iɶ�ba4i���e�/@$��Q�]���N�v+����6T��t�$�VZ�H��[naPM��d�{*�:�ާ�X�b�dP��,w�`k�}�r;
�6(ڨy_}�H����)HZz�o;W�fv_�<s,�H�U�.6�W���!{�]�z�)C��=��3�-�R���/��9�fm1���&�770؉�|3zf�Yf̼��Oi�������Nʡ��9���O8z �E�{L Z!��lUē�Bn+SH���8!T�NC����U�����}�Z,|]b���iP[c-�}f����~? ���7Q��b�{� c��xigY��o�C���k�咿�T�Gvʁ�����l�!�3^�i��$�[2cJ������g(L��p]!5}�p�.�Wj������{]�,���>SN�|��Cp����rJP4�*2�����.I{Y��z�yķ�] ��Uؼ�F~���=�Lt�����y���4<ku<WG��GL��iJ��&���=IM�q[�
��H�.�1p��|�0o78�tֽY��7���&���iX5=�=ŗ���}�>|`F"��gf�,<5�$�p��%������5��Xb�����K�η0ް`��y����������y!�_!As���}9����]�����(���+R�>hh�6(�J�	��b�@n�5;>���z��C����:ܲx��m0��!}za,�
;%.|��͚4��v)c$,wۭ8�V%�J��Ǝ f�W@����6-$L�ת�~���y��#x��?�O��<�j1 �G	Œ���ٜ�Q�S�1o�����ғN�R��}h^m�8U��)�KCu�|�ʆN��8���%ߒ��:�� ����� �@�����9�l���zf`��pJ�%r{4�x�q��zTd(��&mQ�u1��6�Y��LOA��aPo�Z�(<�������&�⓸�X�{g
��������w�����Q���q9]2���or�;� �1m�}Tz�ѥ(�d#�e����	G�AߒE�rj��cwɐr�z�u���!�S��!������p?�w���Q��}�;9���WZ������C�P�ʥW��	R�E�X4�)i�Z�z{ӳ�E���e�ױ#�-OhS��h�C�є�`3�����1�)8D\X�]O�Oh�U���VO�~��f]j�?�!B��`��ڋ�D�x�0�K�������O������m�ꫢQL�F;br�d�K��W�^ �ɜ��xҝ�yV�E>R��>��鼊�.ō@�Ÿ1�{����^t�)�7�[3�y�h9�kg��I׶�Ϣ�P�_B��H!Bnġ��> �������z���ٲ�P��nd��2�S
p\Q�J,T2��1�����2)'W�9�@�H�z�3P*�xf��]J��xa0�h�H1toI�Q^C�'�fZ2�e'�#b��҂=�
��f3�/O�������,��F��#4���F��Ap��z�l�#�S����Nz�GH�6����>���.��ΰ��3��Bl�(Qo�ZU�fO��.Vw����nU�Q�s]�H�b'e�j�qT