��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_ �c��2)�}ma�dظ��v}�b"@@�c�
l�bx���,���M�4A<�r���w�$�S߇��`w���~p�lV8���
��%�4�0Q�Hj������8�Wnwx�5|%�B4|y��<���C�bA��T�N���Ζ�:U���J�::��;��B��O����k�q��Q'�O"�h$ZrgtI���IB�Q��s��P=�=�F��Q�4d�mM���v�#��D����)0 G<��^� �_�\�y(����¬.��	�y�* ���Ob$�}h��@y��y���ѫ��A�".R�]�hڳ��2��}Έ:�g�wQ� ��)��E�w��V9w{cJ�d��(�	0b�9k�X�� mKٺf�רZ�[4D��<0p?���T�4)G��L[7[�4�l+-
X�tv{Z����N�8O��B�埑{�	"�=%����Q�FF��bi@7��J�5V��n��fo��; ���Cn��m�s`%s�*�+u+��p�m�|:��d�%Oʴg�6�A� i��8��tK�K@k�W��'��X�@�0���K?n{ץ4Ej����=��l�=
q̤��+'<�-AOU^uO�����h��E�!A�M�]������w�l��C�h�a+�����?���{��}e��_����9�O�н1���8����J����j�H�R��T��f��ڛ�.}��դe��;rJz~ل!���̽v�Q(����O�i:
I>{��d��Q��r�D~;�������wB� �����AP��rB`�\$�Bg�E��Xzy#0-IA~2���A�K6Q,��z������JX��	�����%ӟ�ݙL�?��f"S���s��w0e(s1<aj����!Ԁ�D�0���U;{�<�棇j�2��k� �/.�uנ�J�P�eR(�H�`M<bA�����"هh�d�J���՗�]1��h۪��ﲒ-)_lu&MW�x�F���S��W��4�9���{�����<���ɂ��b�Wu�jF�ɞ SX�,F��ypLH�WȨ�%Ÿd\yd�%�lJ��VΕ7?�����Mg�ܗ?��BTDr���M���W��:�$���2S�����w~͔ڴ��hӳ=�AʜE�`�/���+��S*�K������[{�o�m��2_�������[�2a���\ܟ|,`�.ޗ��+J�bD_K��`���
�q��Amٝ]�%����]���H��r���+�jj���Ә�x	�A�q���LM"����H��6a��#�$2e�3�Q@T|}�>2KO`&�1�f-��PU�G�n�z���6�5���k;x1�)�Е[����˯����[٦�.���?��%
���e�V\-�@��[ד̣Z�ٴ� c������6�O�\�ȳ&z�{N��.�ǥ�`��#*zz� (ٴc~�`�n��6��m|S9��<���bYG2�ѿ,S��c[ [k�Ea����b	��xv�?X���פ����n���ZM��7�p�
�)�����⟒ѩI��v��f�i�)�۩\�������j�����)���:�i."9L\���m���RQ:0���+ 7����pHL���8-Y�S��*�o�k��S��6��E�zm[pKE;�ߖy�> ��:�X	O�_�� �YZ�i�Y �ajM��GC) �ЉVV���)ݝg�8&U���u��v��p�C��R5�z�/����r�*����}�%״���a�A��6�����GN鱻A���1�ؖ.GD����,?��S��`V�d`�ǵj�i5ʗ'2�6�?��sg	&��R��k�Ò*/���ː6�g�i�����j&7i4��8\��Q-��y���H�Ҋ	�i�}��d�oH�(���HI���(�4^gLd���@?����W������	<΂<Wr�$��{��&X�&����H�����#��1�R������Ɍ�s�!ƈ�a$���m`�.WuUL(��ϗ6�y�34Q�/^�z���d�I��Z�t_7��|���y�ͳ�-��_J�
4y�ŏ���&Yo�V�#�^�Vs�p��2�2�V�e��Z�RlyҺ�Nw(�)3uJӆ�o��iJc�2_ w�';"�F3#t�i�S���T�WF��V�>d��d%%,v��r��+�l#i�p��",��{˶:iW�o�q.g|Q<�
&���~=�����)���,l�A3���)��s���� ɽ*a��Z��ϳ]�Yz�)������a�ߩh��xf���s����]s��K��ĩdl�1�ض�O��G���C���T�u��ǲ;`�	f�z�A�`�p�B��]��\G���4��l��M�D�m�1�<Jz�*�h�d��h-��ݗ��c]a�d�m 3�i2h>|j�C�aG���+�iİau��=Cr�S����H��L�j#�-�V����5��K��/Aq����v� �E�����K'�  �K��nG��ӌ��R��O�@ A ��N�ܵ{H�P��_@v�����\�]�gh-\�G��ui��Q��_ff���BeSˏ�R������24�$#�s�4���O���p�bS=�^�Cg��P���f��ŧ��Ur�R)߆X>�Z��F�S,Hz�8$5���Ա=X	�`IW�\\S�k�ߕ�'B{npq-}k�p��ÿV�K��C���u�4�Ĥ�������}s�v��HT8�*���UV(X��8L�,Iu�q��E���uRg�����򁆄.T|���B���T�Ԫ��32F�A�L�?E͈�-�V7��2d���r�C�ձ��\ y�ƓerP���*Xf��}�1�Br��C4F�|3.��IK�G���kN�I����=g_o.���s�����bQ���h�u�F��F?iO�=??P�]���9BJ���h����}��0���)������u�	:���)��W]<�Z�Q}{�Gj�;6P���3	R�[a�������n��Bb'Ȋt;aN��02Kw�H���Y�;���`��,a�!��J{+���jY�/��8?I����(�թ0퇐j0��S|h:��ǖïb� �u��mDcx�t��}z���L���~/���><sAo�G%)�>{[ק#X�S5�}�emE�5oxq@A?�&|Ǖ&g8׾2PZ��I����Í��P����h�S�����3#�M��aCg�G���X'<Ǫ���� �uu5w���f�΍5�W.4mm��1���l;ƕA�1A��1j�N��D��ُJ7n��I%��.���Ǩ��E����n�듯<��*L[?�E
EC`��H�[P�-�~��тx���R�=�9�q�)"U�˯�,o����봎�<�����K%,�����E�lg���k%+ʨ�B /�x����
����'A��=��w��j���H6�@�����I��9�
�L�(���U���X�1����:�~�Z�d�Da4���8A�E�*B�^>����^��$�z�{�U����6>d�wm���-�ӯ���=���M�6��ܢ�SK�Sp��>ݽ��H�W�g�Y;�Z׷�of�Eb��+�Ӑ�1��g��K�'8���I��.l�M��aױ�{o�!	�X!ϡ�;M^`V�z�'�8 ��������m��T�,������͉�M�P��{��U��M��}�	��T�3�w��""t�t��m������'�O�2ds%��'����I�N7�e�:ʍC��v+�`h�2�|z�6j2�.N���Ԩ�*��Ė;%P��怎� ��_A����[�z����۳3��>��(�wr�'�m���?뺁5�n���Ǧm�o�O�kD��;���dD�@������ 4��
�Ӗ�K�'�F�]�b��d<x�!3#��d�b,D	W����3w[�i�H9ƜH��`�~�$�fט�h�x�I�:�U�]���n�x�bz��ձ�v	i����òd!�y���)�/�do⽎=�k]�XuΫ��dM������A�����Lm`P�A�`�