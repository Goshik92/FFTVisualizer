��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn+�b<�ਞ�~L�\��I����5��<���5�
6�@c�_�Yk_�I�'��Ns���m��S�s�|G0h8/��ż-� L7b�_�ʁS�k��ĕ c��U�d�� ����w��	�g����H�ˀ��ͱ�ez�aL��q�������$�|��,%�_N��\gQ==k��mOR ��1�p��nн��D�D��vVn��B�*A�k~�d�� w�N��e�XUE��g�LJ�I�&-M��:�՜�Ʊ<����V��Ld�М?��ʊ�Dˉ�C������ꎘ߻>�=�#V����πk��8n
�P���I9��f�����R�\F<�]y�C֔�� ���qt���0#�]j�C^*��/��$㣿k��z.�cLl����RWO@�nm�%3
�Đ�"A��/�z�M��H�ȱK���3����dci�Ҳ1�=�m���7h�,?PIT$$��_>�R�O�O�w�	gƸS����B������-46^<�ce�2a�>��?6\�����D)D�V�n����'Q�d=���-�㙂^S�|5����W�\:�>�s�d��-I�\&��_iW�/˝鲍oխGr�])��
��MV���F/@��] �(Fy/�{��)�]ai�vo�d�'�
E�@�鞽	Z<�������cNn�>����>|����Kt�@q\ٰZ��Ü�q4�y9%9�jT'�����>r�� �j�IK��j<����x<�w�h�����=��H�k&,6ޓ�9!��A�+Sc�Jr_]k,�xw��R�ߝ��t�p~p=�+�fl%ıh�G�%�[U�_K�.c'�C�l��_fX5¨[~Fi�.�B�Rs:�M�#�h)'��I����)�\_���Z:������4� P�
a�Ί�D�n�#w�ƅ1V}�)���m53p\>̓�荢�:�­),�������Oj�3Me�ZW���������w��
iM�3�<�`�a.w���7�����ϐ�7�5��1���K��35y�0w�B�}J��1
�Q�i�c��/�r�5r��u�`�~7�=�$:��#�p" �n)��(rZdz/�%�����-u��$�lB���/y`/EeRJ.|��xq�U��J��� GZ�UW��M����:����o=�~k��V!�:�%��(���ic�9�o@U�����Ɩ#ȼ�8�V��n�'��(�k���N��s��L$̧ TW9��C�}�]&��B�u��|�9S'��?������.X��)JLo'c(PX�{�_0���bck�V0T{�&����·�/�n����Q�lu�U��[��&PS�Ρ�9�$AX�]��~F�"1z������z�|MJ�J�ޯ��?���8��6�J>�b�v�&u3椦��8/��<gJ�����g��ͤ�&1o�OI��Y�t�\/�M��}��
ޢ˘�32o�f�OÍ=Y�s��ЫD[+�=-�4�)�3�s��B���b����@h�">L�x�|(���R�_Z����1��
36Au �����X��RR��<���\��˂bS'�]���\���씜 �
2>v��)Y�!Ӭ�g�jW����!�I�pA�����y��*��0V�>YȌ����Q�[�l�TqŮ��472H�&{�I��yW��O�ҟ��������ڰ1RF겍�������>y�=�m�-'uiu�ᱞ�t%�ơ���Hc/��p`�Ht~l=L�53��&�K0x�/���ن�j���s�F֩�E�N!ӧ�3y+)�����ُ�$/�B�N>�rA�G��ңz��,ԑ�2��������Еmm��j��e�9�G՝����0���vpA��>�V��Q �o��tmc烣<�pdq/*hn�ϖ�[��i��lpM�I�Ɓ�2�Ψ	��XT�{���:ꄐ�=�|"KS��4l��'x�8U���a1St��|� &E>�V��������=�!�ͼ�)�2�K�T�x���A9ꐗ|��D^AD>Y����_� /9g�P��Su��~[&��Z0t���KRj_��Ia�>�lCg���U����o�Ȱ�t�B�vv�b��B"0C�e�F����z�� �ǈ5�{D��'�1Oԥ���C�jC#QB�lſ�=���*��i�����ﯧkh��;�6����D�����a�]<#�t���k���b��l��niq��#�#��  ��_�ބ���E@��~���z�j��6WLa���vaZ��)�������y��GN*xs���z��Y7~ީ��d	S.l�A^��b��-�3�@
S������1ls�Za�O�6k�:#�l�Wׄ���RXk��4����g�+��� �6qu�� �鎯�����MQ��f�Zj��U,�-7�i�bN)��nፈ��>j�;n�e`��l��n�L��J^�hN`�o������ʶzY9�x��yB �
�82��Hx��;yFH+%:!cn��X\����+�Yx�%wQTFk����-��Co���n>��mu��P��3��!�	 B-Q�j���lt<������s�>��P�(;���*牿yW�~��W�/W15\MB�J�WM��ԇ�p��&�0s�)G���� ��X���h�ٱ�ze�0O�#sb4}����љ�Uҹḃ8b�06�sj2���r��䈪�x��l~�@]u�)��O�G ��'6����Kh�-��pN��t�|��N���9ܹ����d��ݤ�A_�r~�tS#é�wmL�R���i1A:��T%-2/�$�&
�l��ņ��h]ď���6<_�/�+E�I��u��a���Ұ�,�Wz8J����/��卂�1`�Q@Ss��&bY!/ه�nglUٟ��
�D�!��~=���DP�r��;�ƕ�w0�*�}%hQ�j�3�L�ث&����G(NRNT�N:)'���{5M����ukWm�(��<M�6���'56<#Eb3}��d��E�$��5Mŭ!9F[�Q������l��5��y��Uߚ��PѪ ȴw��f�$������s:�=� ��rW\�-���@U��J�
���
��[A�l�$����K�N'��Xk�q2��Gto�w���/7d���C��:Ne��IV�GW�ui��3~qS�J�k�׭r8?l���]IHO�1U2{#�GN������FJ
}�YN��-�ΐ�ѭN����rl��R>C�O�4d׉��ͨ���,��:�g�^xz�W���x$i��ȗ�5`� g�!(x���?�s�*9��;_m]6�)���8��>�W_ڥ�R6���y&�(T�qA���B �u�'HB�U$�D�B5�le��.eis��k?v�Mg.ҘZ��Tpr� ��c��.6B�$�x����)2�ty��Fs��Ps���,"=88��X���ŗo#Z.��tK��菜ӊh�w�mj���=B� ���Tl����
z���9�ˋ��V�:4ay���c-л�S��m#B�l�mOjsJ]����ӆZ�rA��b>#��Fu��Nˎ��c-�c"���޿e���~{N�%6��7D\�
-u�,c�*�M�b}�ik��7�"�Ԛ��{��F@���Jn
�����~V1\����<EK#l�f�ؑ��eK���g@�� �Wׄk��|k'�݇G�g�a�X��f�1)���ێXhml?W�`w�f�c\[2�;�~�-�g8F����Ѫj�M6.x���j�U���U�Q��>��b�����w�]|��"����uތ����@5�����xwf�nP|�S���'`[�=�v�ʽh�[�n���G|��h̿��R�䃑!�����ɇL(]T[wi�\��3���]�x!-ݫ��{n7�RJ�\U���*����1��z,T���_�2OM�Y�LX�3Ԅ�B	�)�΍�V0Z�Qy#<~�J�Ns�v�L��0���VB�[�He��¡��7�&����cg�XF$$c�x�� �ܢ�������W@})?�j�yۺ�>��
>���tq��"Ųrq?��+����6�q�G��θN�^מ�qL�'[W�ʱL�u�����C������m���������`���E ;W����®�MŤ%�>A�*ȣ���<R���z�͢��ƝS{�|�D�%��/?i��*2�5����;lP)a���&�O�����T#t���D��T*�[Z>@PP�|��H��O(�z�i���,yG<5���6D�."sǍ��)����0	�p�W�>��z��w���NT�JBءw�{�v����r^|1U�-c�N�$�s�pu��z�%ڛ��O�1[�,w9��u�'` R�ƴ/��$�����fh#�|���)AZ�q�8��7A���{����;!��gʌf)�2��c��;��mVc�7�����낑'*:��̾��*(�37�����bx!/\1F�����&2��2h��3.珅������&q�4V~f��D�!���r$���y�e�N�N#A�lwi�H��P���y���9(Ip�7� ;īS�Ĭ�z�� F�ߝ�}��J*�R,�I6��b�����~@}d��:v�)?���@�/ZwGB�m�����7g{�cӹ�%|��"�A�(H�86m���鈝�dX��{��>�'
!�k|�kE��.ߡ?�G��S��re�;ٗ�l��d]�c�%�F���b�G�����K���ܬ\�m/�k~����y�qd���̎�\����H^����� �����LZ��~rcn�(��?\�:9����a^�!U5���B���y?"8�/%ļT��iK����_��㷈H�;*��S1��
�E�'h:��Q3��8�d"fڊ��31T�ֿ�w�oùQ����T�-�g�/"_'�P��S2p�*	z<fi�s	D�Y��������OD���[��.�A���R�Nd^1�gY�$�B�sl��d�g�;͔(�ܟ�$%�.i�xW4��
 �at�J��Ƈ�����r��R8�:�0Y�n�u��l�\�k�"S6)���r�6wnz�R(>�}E#������H�ud�s_�3���F3�'���F�����i��O�)W
�m��ږ�c�PX��6�mxm%ڐ��X�:����\ɓK�;\k��VB_?����b�`~�.��_�;�id@��S3|/�����O�i�s����3c�c�X���̙��Q�&���
]��������b�U#��V<U��? :��Y5q�$�ɥ�Ǻw�R�۱}�-m^�}��bq����[���[,z~7Fd����획�D�'���9�� *R��k0����L�g��yu���3�C�V�Q�v�f�0ϯ��ME������2�	X��&��~ː�8�����`I�!�B�Hl��Jc#���A�n������q�ץm�z8.�����+5�]}c��4}���\#:�\.
�뙄���{P�+]�T-_��<gC��'��':�g�c�s�,�3�'��$}'h&�^W6�䖢Zo��szB32���da�[�Eb�%X��r	DkЪ+W�(�bc�E��ѐ�����+��M���MU�4��Ĝ6oOKs"�Ĭ�"5��η��m?x
_�����zJ�In?�OMz�<m�^nU�R͞�/�Sˉ&�&g�I���=;5�vtC�����7�U�7Q�j�=�Crqn�{pq�ᖛ���&<�n�?!�̾m_ز8��#� ��1S�埍˦X R���:�j�W03��!&�Y�NJ�/���}��)I��h�T��J/I\�����m�`�i�֝�X(?�L����Ty87߾��1e��}����+j��w�I��ֱ�'�لF�.
{���64���ˑ��H�]�����ʦ 2�HQmj$�|"���G��.��j��$�I�@�<�����g��:��@zi�q���tݱB�E���]��hѕ(�}?��:��ժ76O5$Ck��i�V�a�>�\"t�n(���Dف����c@en���t���7��3I��ճ���>x��}#���R�e~�})�+y�߷�d$�E"M���n��c0lu�)"g�������ש�4��.YO��iJ�7��1��|��b.�5E�9DW��#U��p7/qaz7ǆR?��9��4j���z4�\kv+�|_X�v|���֤Ä����:�N@��JIOT��Y �h��
��7�Ta����
�)_�F�lPXb�
�K�/Wr��[hz৛� 0��!8p�@�(U��T�;q�PEy1H���Ph���("�8�����弬��N�կ)��SFg��U-�X����N�>D��a�0�^�̃�3���_�`-�=|��wĹN�g�ZX>�_�a�*w5x�,Iw�@���E�|ƺ���
�Xd����S�O�),Li~�X��O���g�.��婽�y��~����#jL4R1v��]#+i��$-�}�r�m���c��k��o�l0�����!.�(&�
��4�2�����Ӗ�:}&��j�*�gPp�| �2�3�m��8zu�،�/�Cc,$ېf������&���E%�GS�]�R��@�!Q�tkS%$}�D�����}�-n�vDb���Ǔ�S��7O�%�6�*��W�P���y�%�v}�|I��eb��B1��GM�kjӹh�k�S�z�J#Kњꙮ���k�����^�	r��{,˥�l"��j���YG_����z=�����w��2 �t$���;�}!fo\��X�j�v��P�E���h�|="`��`k8�&��H�vFٵ����a�!��%E�E�:D�R�r����R3s�(s
!˛wa*�1!EК�*뿃�u�������u�p�Z�0��8���Tw"ǆ~3��Ό���Sq�ը�@�Ej'9�m�v�ݬ��-�������P9�Q��㺨��3���8���h[�0��FS�C������K\~(H�_qA��P�qJ9I{��mY���?��7�Oɛ���s^�~�v\���"c�$����ϡ�o�ЧX�D���^C����*�:�����:���F��{_�!�Ƌ�0qX�]�P����y{�k$�q�Q��bI=�q��w틬��M�{����:��,����Ȱa�N����C��/�i/Y�q���C��UE��5����=U��5�
$����R�6�	7T&��SF�y�@����o?������(,�2�#f(�}�|�M��LG\.@<��pg���wf����a^!�x��0ca���7y
�Bz��O��ά������u|���T꧞!����o)��."��z�,� r2��A.�S����;����ΒHu�� ���>oa@�L:Λ�4<�?�|yõ���h�a	�s9pN��9!���W��A�a��T������6Ƚs~j��Y���FǥŉgxMD���*��SZS�)=�G]X<�_���b��B]̜��
r��<vUV(mC�q{\�[�����3v���ρ�+����x��[b�%AN�y�E�Zi�]�yr�p����
���\�VleǾ���~�C�Bqc�v&w��?|��d���[�6[l��:�Yח�Ԉ�U"jEii�maN ��K��	f�*먂�
��h��O����c����g��d%̈́'�W���eӶR�� ���i
�V�w�o��(g�B�
:qOC���\�v��+��,U�Qvs#��˻�?!�u�;V�5H�.~��yNs���䜌��=#�'��8h-�M�q�'n��T~j�̋o̠/K����?B٩QQ���%M",�f�����U[�]%���l��~�gr�hc���  ������k�)L��)���ќ�If(8Nq���޼t^�F��w̑���$!���fj��ݿ�����)�C�GR���Ϫtm��-^s'҉.(^<B9�^�V%빧����ޞ���jC?/so���'����\YZ�<
��=��V\���΂(U�P�ܘſ�.�{pB����!^a����\髈��-il;�u@����RV�b݄B�0�BeL�{��b�H��-��;�Hw�W��r 
�*Sb��7mL�DHV�����KxnZ�5�>"q5'��[�A>�Ñ��x費�	&��W��6i��]��w�,�:�o*oq�8c ��+�f^�|C� �rR�������Iv_��Ot��%�x�Ş�y�j1}��x���lOR��g!NP<�ʁ)���L�'�� ���c����S��ޙ���(���d�UMh�I���}g2�c����(	�V'�i��d�p�s����?#"�3�F;��f܊,GZ��a���=4]���P}��Z18ď�b����[������mm�P����j8�j ��*-�[w(B���s����=)
 C��{XT�䶇�0�֝�ܰ<��5�L�Ɇ5���{9(C�	Oj�P�i�dN�̬�y�P�--ɍw�ks|
�D�؈?Z�u�`��d�e����#�3k���+ֽ�w�J]s�#��.�3=lO.�'y{�)�/�S.~�i���|��m,�a�/�\��p��*��`]\]L�B7��J\�riD d�|�n��V�3x�,>�z�z���(���\���#>N�}�^Qٖ�l��:`���s#�-���r{%�P����a�e>�JU�0���%�2 Y�цN�
6��0V'�Xt�A��k���^m�6z�����r�'�eMY�i��\�GF+x<H2G$�g8�粻"�Dά�G�~�>���
4A�#���$����r��x��̘k���S>�fZTCD����� ��|��0�˼�{��X.EH�~�!�+d(�n��X1%܈�,2�0��5@FWl[��X��qA�=iQb�[:��R�yOD����O�>�N�iؑ̓Դ�"�n�7tZ��0f/�aIM���S�b1��X(j��jIT�l���6�:����-�ܚ�,��m`���Z��(����z�xZ�� ;�t^��y����K�}Q��;O��A�Hg�y�0�N�H��*��8�o�Ȭ��3(���Zp�zJ�I�2v+��*���@R��q+T��3$��k#@Ek(����A���HY�k��2%�Z�<ѭL�`JQ���e/�yù9H��v�U0iO��bW?b��0J�U�H���6��βgul��;�N�߸f�x�J��6����k�� z�A�I)�����^N�c�yX�p��b�{�V��C,�(7��N��\k*4g��ZwrT
������d��0:eZI3!�\�\���V,yQ���K�\�7E���Fܻ<����}����51�R7�,C�r_P���Tl)���޾ԅ!��]�i����g�u0e8ܵ��8��rM��\j=�K��e4�L�������F5b�:��Y`:�+��&��)���V(�����c���Ar8[Lb�����E	 z+bסo݋��I��jet�
��&��Ԧ�^1p�;6�|��(�?�j��sB%�9�JD�-���L��/M%���G���\�Y;��Qi���!�E�A�/�w�a�k��_�a5��?�]���6��Ú�
AB����[�i%H��W�����|�>���UY��f�A0���˝���H������K#�MW?'�If�=�D�xE���BB7���n�K1M��ܫ*��C(J�4c	�Q���?�<�{�/:�\��79�K
�ߔ�5u�d �9��VS%x���X^۞)6����r�7��P�Ie;�H����HPϤ�"i�"e�h�g<�%D���&KF�YZ�h�qr6]��h\�]���*�#3C��.=(�=��]�c 漴=��%�k���#�����rxN��$㬥�v緒��	 �څ��m5hudW���A�Ozj�5 ٟ�ހ���ϔ���?�n�u�J������d
c3��	Ӫ���k=�AנX�|Y^VJ�ji�5���e�/&��ي�MN��E{�J��<��IW�	�����ˤ��Q6���*�BP�n��x��k���e~r@��<�]����)U%��S(g�b�Ypk=�C74e��o��3Ԙ�N��Is��/����n�v�>�Z~�,�Q@��.S�l�Au��v�2K�5�>�pj�Ԛ�IhhGi9!F� ��[���_�9�����T@��<�]4�z=)��ȍ�v�A����;����?@ 
�)�fx�"f�V
��"7V���aL{
Q	�vuD>��W�q��C+]�U1�a���=���vѭQt"	�y\�H�`����v��e����8*��L`�ED�|0�X*�!W���8��^?.��e-�� �S��oQv��9����Yk��j�"���vz�21Ӗ��pJ�
 �[�������#ŬďU��˗�nDذp�L�;�a�4v����;��qkԖn�z���԰<�v�o�i�z\�����
��*�����Q�Z��M5��ޏ��X��M>�Q�~�y'sC-&KW(�~��)i����7a=��B� ����މ!W�F⢧�Z�
�7��˲����R���{�J�2�K��C��M����z���xyU���=���~�ǭL=�����6�xY�<�kf`%[ѯ���[&����T4�L�(���@�	������wGQ�/j�F��M�!1۪�#�R���C��F5��h��g���������z��@���MP?�OǊڞD��=�8k+�ơ��pc��S*�� ơ��Ը�3#�d�������c9�J�H�A�{�;3�R󁧃��ڃu����\\|�:�Xߥ��4 Q��%|���s����5جo�L}�_���ڥ.#����1'@�čJn�7![(s�J�G�#7������a�3՘H̓y��קS�V��j[�����j�<�f�ς���_HY�~����Ѻƪ�9h�%E]9��x�Zk_T �k�3����:`6�
���T�}��L@��c{�>�]3��YW!\��eh��P8J��[F&梕M�����r�������7%B.Z 1�JaPs����HM�4�G���EY�2��d��
��wRĭ
,&�=m�%����)���t��I�t�m�t;�Ay�Co��<��9�`"?r��x��3	R���v�S�,:�*���<M� U���K�c�O�,��q`��ڍ8	)
��m�Y)+*�u�	J��{� �.ٗ�Pxp����-q��ŦY�Q�%g1�tN'�%���x	<bY���0�
�g�۳��ڳ�M������ie��oL9r���HB?F��sU(�|Z�y���]'��P�g�>������dr>��ul}�f�,< N�r:�W�b�Sf��q�B���|9�j�|����� rٛ���h=e-�	�N�ѥi:�#E~���[6��9��
=�92\��f���ٗ�4�:j�eS3�	ՈI���@w��;]ik. F�{��U�\�X{`�O����W�
Ɗ73��Z�<}C�%v�� fvX��A8�m�~�&j��o�S�/���0�T^��'\G?]����A)�)������~��J�n��#l��t�CEJ�^@)��y���M��0q]�̕=��ĭ����t�o$�N4���"܀���A#�ںʽ�Wj�G=��^�h���8n�	Su��uy������5U�ʎ"���9��u~G������w����{�$������8��kd9��D����uX�vY�4��wVT�W������x.�H��}w(](�IM��Pz�wߎ���0(����5˟`ɒO��� ��u��g� �˅��*�C�v�����<�ʐb�pі9)�s�v�ԗ��e�vy�y(�l'_���vh�b���V��+���� ]V���j�+�E���-�&��q(i��u�p��h�fD�*6�ˏ�*�T .U>�̈��H��~[(6���y�.�kG� �\	+tV�����2�y�EI*z�4M� ����Z�~_���w����$�����r��n��T���X@�~)�`͘��6��N�բgj�Δ�!��Pb�2����DB��8�p�"ly���Ъ9�~�:zw�*N��wT�s=�D��6B�_O��h4��_R'�&�y��n8�>��"��M��3rD=J���(��-�\5��L��0)`�-`ӽA�n�����%Ӏ�;���w����W�(���M���1�����e$�zӶ��TDѝ�#|��R�f�^������G��_j�=���'yh��!�ݓE�F��[��¢�)�G�W�Z�G�����rOQ����]׾�{E�պmtl��_��0�:=q*�,�;nbZ�P�	v-�0�^��?ܓ�|�D)f�[�6��A_�<��y�5,u*a���R���*h���G�"7 X]�U�㘤9�k(�x���5�������L��LȖ	���Y����g ��7�@��c	H�})1��׭���&@�����y�ʃM;;L�hJ�P�uP4d�[�8�)/��-�Xp;Yů
v��\W�M��S=0y<	6 Ciz���l*�od��=<��,;�\���m��{��a�̋/u$Y��҂�8R��|�O���8R��V�ȑ�-t���'[)]�'��e���}�0#�e���=>|��k��t$�(��B�K\i��0Q��A�@�2��3��yV١�= ��'���%L;�1�SG����^�ӫ#�F\��z���F��2>cX(��0Si%~����(�Q丣cߐY������� �(��֙N���2�Ru�2sRE��^�a	v&1GQj�:\=),�E�����+��.�tѥ 72^�h���~�-�=��A(G����T���'����f ;�Q �y)�ަ�b�o4TU6n$����[d�U��\;`��ΐ�J`F% �ɋ�d�5�S��l�A}�ʡ�[�
�WK>�4c�\���C ~�$�1WI�M9u��M����Wg��_g��BO�� �H��υ!�"�0�	�p/�ذB��Ø��+%�/Y����_n���u{4mn=��_���l`W��a��EP���^�G�0��[w1ņSP����pw�-��[ls�8y�FnD,hw�ׇ�v��Z�Q)q�j�A�"cX�^�X)�HL峗�qQ��"^�%��'���<�n�_�L��F׳S����̯T΋T7�s(^�vK��c4	�nR�)4�伙��7c��#���jw1nY눍\l-���0�J���0�Ty�c|�orK�ּ�3�z�r�$���f!�H{��!tJW���j�Stl����?lV���ѥ�{��Y�bP��fg' [������}-$��>R�wx�tHLc���N���Z05����,�cdI��%Vңb�a�`1Z���vyu~J�>Q,O����9�����q�x2Շ>��X�T8U��l�Z�G�68O*��i���I��c;N��xW:ܟy]�H~̴+��ѥvS�[�bI/X�>��m�knЪO�w
��\E�҄sج)�J�q&J�	i�Rn��	��lİ;)/��$-� {N�UEg��\V�[�6l"i5������I�"�KH"����$*�9�����,�-"R���ȍ�G]Q�#��	xƖ l�-wP�;�#�ܨID�W�f>]�6-p�4�à]Pա���>�F)(�%a�f���'S7��i ���b뻄3�j-6�|�c�c����n�UO�!�Wm��c�=�׿E�?z��Y���*�w��ڦ�4�2B�v,�H"[���+����L���C&��`�~��S�г(����#���dz.�>׉�'�i�M<��2S�LS�E(W�8$�D�ž���4#�c6���D�<)M����B+9�U���ž5m�R��sf����!!O$���[��s^��њx�N�(13�OE&`������ZS�v)���~Vd���33��}���*fd������� Z4�=�#�o7n� ���>v���9��]��Q�$����Zj�O	�k2�5X�d��4b6�������7�KK�#<����2��\�M'JB
y��ś�T�U�/_���+ǐT���Y����L�y3kBΙG|R;H��"F	����j�����q���mD����8}���oA#���du�Ψ`U�xdR���TK鑉C ��z�{�Y킶�(Q����W�-ai��$�!�ř�����Y0��9�Pf����_"�!��ϊ��,b��T^4URcL�<�z��&�oOq�8�xlY��^��Y�����ͅ&Kb�^�2��:1���mv��{�B>t&G4�)斁1�+��-V��U����;��v�|1�,���?���:�.,\ng �Lb`#�I�1?�n��ab�'���΄Q,:�ڎ��jk�C@��be�����Ȼ��C�J��
�:��M#4VY��M1b!v'��%��ϓ]���7��m@�D��&1�����;�n7ު�"���1"P'=7ɉ��2�ѓ	�39��8s��0�8�o��j�%���&�~�[�c%j��}�7�T�+n�h�4���8�BY�
���K��ÁrB�C�@���U'[��읷��07$�Se4w�:1�ݥ,������|[��
8s��3Y�uA�4�8���H>��H��p���d�un��䖝�$����ҕ��q�4����i�{ڜp=G�Q���zs	+"���|��+?|����"Al^i�<'l�E�q��$�񱐇��b������u��l����:��;�)���w�<�,��_��o���N`*1�!�����+'�+�!G��UY��MB��aĪ��}���J�����C�]8 �?�	M7 D�Et�J]'3-�S/�kC���5�?ֳ��
��C�ߨ\��mk�?sx��Q��s%x>0��|g�3����q򼽈[��$*&�Bv[�@���N5e�	�J՝�=��ۿޮ�B��G0�*͗4m�������h�q1?��rdn����o0L;W1R�6�f�^[J�G14��̀��࠰(�_PTo�}�Cp"HQ����&�n���HѦ>=a�u�C��ƀ��n<�4��ů��NF� �t1�Tj[�ļ�ѩ_�Qr:@��s���<���o:~��ښ���h&��)$tCɵ��@��U��p�
t�d���34�����ڌ�I���5	 J��-ݓ6|ԙ�|R͎�p��==*�WWŎ;X��R���Q77� �=6^�OB ���w!�x��Eӑ/�����UP��.�]���`m����A|��gΛ"���O�A6��Wx�_�ۧ����p*K�{��'�*fc&�n�S9:�X�;W����fZ,�y급�%=ҾNZ�b�[�"���|E=�A�wY�%�7��):#F������Tv����޷�a����Έ��#&
+rU�۝2�4��EX��d/2�`�y��em?Q�$��b��G��Z�'�f���]�R��*��t����	������N}H6L�����a���&�����% ?/�o&�O(������=x��}��n��[H�m0@����V ����>.Ku���w�U��ALW��|������3&�fW�/��г��Wb�GUn�=���O��a��s:;��T^�2\�f>+8�N�/�B* ��!h1kZ֟B&6k�xhG���0��U�����MQ�Tg|M{l�jS�u�2�V�܅�������?d;M=/�SRIt. ���kQ>P���0�j��Rv�n9�НJO��4M�Ӆ0%��:!�����W��j�}m�'�(,���jt0D�j�T��Q,Kn�:ot!��^���#�7��E��4j]��/�"�,Hd��	�l�[�#)FA>�S��^�(G�Ғ����:*�r��y˽�gs�U�ġ��L�T7���� �T�9�k��S;д ��v��k�$*Dgy��\`��.g,��A��E���8���]�a���2`�VhMg��Hq�?]�O�)��_Ƕ1�f�CR3�ñ����iJ�%�pu.{uQ�x9Jɲ7��Dq��)[����F�9C�A�����Px������cQ.����Iٌ)J�r}�N#�"�����O�3��+��-�������e3�f��
�U��Ў�)t���𩂞�����⥨J�l�[�gTO����y����?7ܬ�R��6�1
�+bz�X�y+��K�(���آ$_�[���D:�%�ģhgD�ی	M��U�������Z�*�{�P�	qco�Xw'sȓxZ�L��Ӡ�~����m�Q�|��Ŧ����jKL �([T��oy�څɀP��(�6��T�x�j	���.����1��&JЗ"��d��Ə]ѹ�nD�^XU�0Bv[��jm~��]�X,���9�nτO�6�G� f�!�-M��h���"�LEL�Ss��,E8�qz���ũO^�jX9I����n�`��E�v(���0x��"뎣O��/���Ru��;�O�{��͵�Z��* ��o'`�::�ֺ��H�������Xɮ�J�ݙwF�n)��%�Yv�ޭy��?��c��	��W���2��T�/� U�����M���=9�u]�#\�g`�}�H�c=RV�r�C$���Yg?��d }���t�5$t�� t���wO�5i�~�1��!�2�Gr�����P����y��m�hA'鈘��m9EyYZe��<ҥl��4t��"�kn�1>��F��M�{�sd$��������O����Gj��}J����� y����Ƀ�D��yy� ���C~�1W0��;�sJ'[ԢV5�n(!J$�}&T�(�e5��kA�� T5A*��D��3u�|�n�<��X��˖��w{t/�tr?N��5�F;�'Qs��WQ����I|]\��JE���r�W4��*�� [���Muc�-�����3Q�!��%��0?�<˕ ps���8d�֒����E��OEV�-���Ǚ%�����<��0�)��dw^��a/��A�gH��AQ�dm���
��,\Q�+53��o3�
���N��g�;t*���ϩ'xr1���b3�īRR� Gd<�U��@���i���j~�5#͚���w���]�e�Lf36��`��^zQ�e]����\eA��e�0����T���x�`Mu�f�t���@�[�<3&����e~���~��H��q�^��D"����Y&u���2P�$�	��`�p���FJ H�����ך٠�M#�|�Mׅ&C-�Ξ��+�N_�s^PJx�̙[q�
8��*�F���yS�K�h�K�=D���20�3�a�O�����*��P��o�J��S��	^����k��1��f��p��BML�������Z��r>`��VnI�� � ��U,Q�fh�R	��Dmش�����Ir6Ec�j�����6�5 ������oQE�����2�&��Y|�&��'�zp�&�J�K�,[�R�G�)��D����-6x 3>��"U
q��K�}*Z�۾�=S'�V�
|���~�]���$��m$|���u�ڃ��s6�Հj"P@�&]񊓺
wR�\!��@�i��d�+���%m 7�;�uJ	���h�,���k"<���e�6[��i0������:�o�x�����Z���g@� �Pq�n\���ש}uN�3�P�-���a��/f��`����.f!�
�@I��Ƙ#����]:�Q'��a�&���SC��Ľ8)�얹r�q˒>��1\e�V�n�ŗ�Ӭ�L�n�>P³���C*��k�:�#��"4):�X�-$�x�/~k&�Μw�����ER��Ո�Z��s��+�+eҮ������݁,��Ml��y��a<k�lL���Es������O���d=J/qxD~aϣ"��8�|���p؂��<��+ȨXG)߱�Q�e��1V����8��1���Q0��q,��hQZ߃D"r���P&s#A��d� &�%�;0��m��T���T�d(Y���_7������B���\b(�b�r�f����7w���o�"g�(y�ܙ�;$�
u*�[�V_�]~( �6��X��|�岋hϯ|��3��&�
�."���C[�~	����fӂ�EڀS3QA�=H�؟<�#���4E�+=I�tF����/�<w7���9~���/����9�6��!<h<�%��c��L4D%��$(?"	pol c6�"�X�?�̋<�nF�wl�,�x�b�Z�$#-�G|��n�U'��W�W�����9O��O�����j��pDc��TS�؞U"=�����iU`Z8�f���I�jl=�\,�[�B���
M�Ϝ2�U�
«A��B1;��XJ�S�$Z{��B��_!80P�S�+�_V���-������6��ic��Lv!;�Z����HKF��'�H]�(�^�L0���4r��X���ƽL}ɓsG�H��ڀ���FL�:��ikX��9�C��K�j���W��I�����0'�w�Y�*��̏��y����cOT`�FRR��S~�)�#�^�F��������!�0<4N�d���Q�|��ո諲C"�ۘ��q�aG"?T�l�� ��ӥ<��\�Y��fC��߽:dB%�yub�B�4�x��k�](�6��
s�� u� -x��&H�!�N��*A+���|bJ��S�6��(GL\�e�t$	TK�A�WK}�������K6V/,n�R{bx�շ���ք�[0�O�=a��k�-*�m���H�z���D�h����7h��$�<�S�)s�-�x��mV'9'��{�
z�:`���C����gt۞w�c񁌘�KoA��|�Md�t�z�.�0�����c#z��>e4���ך��էY�����C�C�B�pWNΚ����c7�ۗB�L)��OqB�+Xׅ�O���3�s/�N��[(E�-�e6gi�I(�����+,��1#�H�	������!q}f+�v�J.�i�`�?��$
9��g�� �P�������=���+w���u*�,@��A0s��y5�#����K���&յ���'�!VT��5�a��7���#��p1�N�XK���c ����\܆@sL|:e�XE$y4�Ab��6zK;/�	.��p=�
k������q�+�'�";[��H��`tϾm֚:�<R����Yc��}�e��ćJ�b��Yl?;ekP��l(�.PsR'^��`pn�<�į�,Ak�~l��������9t'���O3����� t��	o�����
tO<��I�1C�Kc����كVߤ嶋�p ��a*t"�h�K#Af�#n��� ��I�l�p&:��= ���x�<N �±�	��63=�t0���������^�J�P�
S~��A:�`�M0�#�4y}���vJ�L� ��@��7�0썛~u�An���ߗZ#$lS����tQA�T��4��%�]�*n��$��sg����\D�CV1�Xv�ٞ�>.��Kz�X���o ��9���;h��d���6/e��:֮���7h9^h9�N�b?�a����☩]tʚ,Y�cM�[�Ze�D)M�U������|f_!9��%�7q9�́,�����-����1�)��6 ��z�uv���֪&��/�%�p%�㣹>����`kş����ߵQ����ճ���0�R�������B� ߋ���0{�5�Ah����%Ľ���yk�W
�mc����k��O�����U��Fa�����fV+�u�"�D
X	�ݟ�Ǒ�`�f�f���c������]2;F�4k<�AK����x���k�,J�I���
�7�[�%�ߝ��5ܣ����{灁͉)�E�̕9p�q���YY<�ϊ
߅V�0�`�^����!�B�6����%v���qM_�������DS�v|3�b��>��C�gG�?me�m��0����1��b��r���Lj$�%!YF��/��_F�+`B��N�DR��� ��he�Ώ&��[a�  j5��-�e�,��p��E��0x	Q���s���E(���|�ur�V�ߍrM�ATj�wRo�0r� ��=��L�	W�� U?����0yU�U���H�P̿��
��)ѦV�(��_��Y���&��Ԓ�,����d���G�~v�)�yz�x�j�N�_A��������F0������B��ޔB\��6��������>�"������vs}��P��h�k���m���|ymGC2��)�"_yJC�M����v��@S�����es>��GT��lF�2�6GI��T��p�w�`�~��
i�M�\i�ԵD	�S޶7�B��3H�GN\���4��7#0A�Q7��X�J���rpD��*})�uV24L��'�}�Qz�[9���~
��o����Hƅ�?�����9�*R1�1*�$f�&��@M�>��t��;G�녱~v:��д�Yy�O[+�NVx-�6�6�C<*]�;�=�6tϘJ,�		:
Zn����닪���M�=6� �ŻCe������vX�:���8��\�C�Z���m�޾@͆�9���m��X�sRsA�-F�^H~�\�@�i/Z���|~�H�Oϭ�V�\��p�UyMp�(w[��U���k��>����\ 4ں,�M����iP:� '��]O�~ �˭�'�S����V�
=7���k4Et�G�����g��1!��tT����Y@�4��Sf&b��3�(���mC���j��'u8�L]�\�ֲ�@kZF�����呵;�U5�W���#�;j-�K^,���Q���	�t��9�c�fsko�b������i�,N�5"����(0hI�v��d{��&qc�, �#���( ����A�X�~���k'U�7�b�E RK%��;x�xˍ
cm���Ӏ����9( snA�r�K�er_o.�e��u�l�V�B��>�C,�F�سsk:.6����|.z��mcA}QZc2��u.��(���D������ߞ^�;�і���ˇCHJ�f�s�T�����Z��3����@�r3M_�z�Z�`�A�����%�B��6<���0�U�������3���!�g[�J����sV1w=c����Bc���w��^c�
b��SNT,j9ODϼEt#́�hR$+$�l��y����`:籸��)^�E(�������JbMI�,����&i�Ʊp�=��t�$Di���:� �7Û}�r)r|�9��5>pj7�T`���̏S(�ٸW����g���[����!��{�R�'�p�+�.#vg�`��B)_EZ-ݓ�Zw3b�J.�Ŀ�!�s��MPd`)�tm+zVE�ˉ����_��g^�����Q�*�yb��S�r���BS�:�T��`L,��)��q����V�/]��Ք�M�@{����7�M�t�#Q����k��g��Q�M��fE�2�<hQ�c��M@Kl�%�a*̆����m~�H�ch]�@fȶ�C3��z�Wt��~A.�ʥ�[�C����r��G�N.b�Y-dl��c�&�o�	������ss?"$�j��@c�xod٤.i�bp�S@n�������
h��=j�g��!��u]3���:ř�_<��v�Bi9�Ԇ�&^�����gj2<A��1�<`QL�&��䙉'�<J&��J����ǐY�b�"�H�P����+��bw���@�]�e��WR��T#�P��&iL_􇖄sic/�Z�=�!��^!���-�1�|�@��v�q�׺戒�^��ut3�r����bU�A�c
��5xbo���Ғr�na#<V�\����Χ�]z���P_x��`qJ�m6��aQZ_A���� ��5��ċTw���PAC���/22��ɘ��M5�s�s��͔��8�&ݯ���מDS?�=�TED��EM�"q��"�$�aRn'eU��̒<���X�}P���eW���S��OO?Q���;xz[X&���*N\��������M�x3��ڈ�����<<�i ���-�D���2��i���F�^�������rW4 �1�^�WF�s�u���f�C��M��"?�8�"Pa���n�!LS�������#*�87����EJW���=�21/�܅�l
��-!\ձ+m�и��b��G{a���U���ʶ"5tj:��:��Ѝk�#\�w�mx�����bײ�Ę�HN~l��D1�Cm��重��_z�қR깿'���@�&����5hrl�2����Ѩ9*�A�����}�U�'H��y|\R��Y4J���F���/\!��f��Z���s"'L�ŗ���dz��F��I�Ps�[cJ�¸/?��	���}�!}ry��ȏ�<��abL�gZ�D~b��v����(Kuo�l��IJ���g#��+��Z5���0���K{�Qp-�bgV$��7��b�	�ư?K�z��F������E��g-|�b��l���
�[�Ԧ�#*)ܖ�y���e�FKzv��� %r�U��sN�b�g9?��M<��X���#O�*����F���E��jd��A���F�d��������W���ҰX��֫��e�V�ݠ��J�φ/Zn�>�pjX+�.a�3Ie�Z'pܽ�Ch��}��ۿ$�|)\O�gd��ízW��=�p+��$AJ�n�)F�m#������,G�$���+�����
h]�Ǔ6���ÙA�y'�lnq����9gڗ�-a���R�"v��A�I^�Gv_^�d��Av]�PTSV���1��o�T��V�Z>����BI%�T����ҊL��\�.݁QB���蔵�3�D�ٛsq'����6X���>a^(,@�AC�n��&�1����i=��"���"whySJQ���! �y��"[�<�7��V�v
��B�`�3�s�r:gxͅ>�я����d:<R����VF�2�EqY�[\Gd�o�ك$�nD����Q�ګ3�t�n�k��fJe)�E���61�zL��h:𔃴�DLc�?$�F(�=0��G���Kj�y1�Tac����dl^M�ű�_�h)ͱ�Z�d�!K��\��<�=s�U���U�;}{ �&��3?���۸��|`Og��BMTD��3��#q&�G��]�q��-�V�Ck��-礋��m�e��D��y�R)�)��^2���iOk�]�0�FJ�ʷ(*k>@�@a �?C$��uͻ�#����g0���3jх�¤W�	c��]��dy?�����**WZ��	�O*M�M���G����-de̀�L�����P\�_Zuz��`#�N�1��5����n�0*�Ң]�� �opJ_i�|�셤�-`�5��]_:�#��Ay!�÷���T������fk/�?B�l�lxm�,*��~�J6��TÜ
Cʲv8lQ_W5'3%��(D׆��k�D�9|b�|�o�g�]�5c��[G;�[��%Xu���k��̑2j��k.�C�Y%`�������8���-���<��*����\~���m�w�"��h~��� ����gץ�����u��컹��|*�;"��]:U�K�fJLL�̑�t����� =���B��)Y�}L4\<��Y�tʪe)�a�G��L\��'9N�����|݂��ۣ1Z�2BTٍu�:�T:΃ܓeX�*��[�ko1H�'@V ��� ��v�x�aU~f��Jo�K4.�+<�݅�,�܃�P�O��� /�
��`�<�^�E2��\�m�Ȕ!`�׍���8����Ms�0�6��gx����M}�,Ci=���9�9���7|8Iu� �Vj���y��-��J�`=��YNԺ���������-�)�5�W������tp��Y�A��~��˒2֕������2x��&q=�4�ז7� �����_=��OO-���pdY�L& -p���?�|�]�Z�f��p�$��kh7�M?n��g�L_�({��"K���d$�a�cF�pa�3��Q�$�٨�����6��1��
(����\@�	�pU�X�t����L�B�h�3��G:�x�?g���x��� WN��za�E�J�P�M��L0� 3����^ɘ�2S��2��W3!opD"���줧��#-j�ݩ�kx��LJ��O������R
���VD��A��PWh
c;�͜'�-��q|��DT���^��gk����P�P�BW��}�NX�h�i7T� q�u��N�73�#t#�ĥ�ٳ�6�p�X�W%q��q\>����$A�׀���{�g�n�ΖF�S��XB>^�*��B��� ,A�����z� v�7�ge�#s h>c;/���nd�ߵ};�p5��{{Դ�;d� ��2���@4��l�0�)�M�m�?����i���A��{�ػ!Ց|$\t=��J�J�z�f%��@�h�G��(�H�J�8��5�N�"��%�B]XE�WRPt�P8�-ل���=_���?םyna_Yu�S\-��MU�l��G�(�,�	�J�!����>\)�|ާb4�u����G�N��0�:=J*�_������O�, �֑�0#�"���HB�)��7p$yMh�.�5�S	��x��
Y�׹� p����;jr��z��mD�Y�P}�~+�C��9��kך�ĕ�?��\p�7�[�s�o�������1ďdј	V��{��P0�v���d�E�tN�:ɏ�pF~��q/�`Ļ��S>�T�tNN@�J�(XZ� �r��k� �tp������2��פPGb�A�7�_KC��d���dX�Ѭ��+���6��R������O�2��,���v<��Xq�=G��Ga����N�M�O�c��w%���Ôa��)ݑ�m���J��9�8�4��d.�m�[qQj��Q�瑽b�3����ˎbB�;4�]jE����h�������xzo�\G��C���JAE`�.%�q����xv�>wQ�b�?�����Bĵ?����P����!�@��x_mB��[���W*b������V�&�F3�%����d�%ȴ�2F�AJUxY ?��k��9��;��BL��B��ܬ�r_����(i�ͽ�&p;7@�Õ�e��E}�ָ��^|hyq��T��k�Q�F�`R��4�a҂[p�nVa�HP��l�(+;����*���d��o�-Ь���՚5�j���Y��i\��Z-xG�����sq�\Zn�N-f��p�f�Z���U��F )���F-$��I��#Uҭn�zK�����[�@E���i��vD�`S���J��e�|�@lNR��}���c����.A�l�����)-�ާ�H��VH`fG��j���*�9��Y6%}�m�A���ZޛJ��>�����h��'�'��ilF3�� �Ϸy�,�bi�t�j�+�:�Ш�Y��T
��ơ
�ϓ�d5)D*1���EHm�4x���@��S�����+�y�(Qc��,K��k���
��;�����.AF�**�JL�+�<�M����,����I��脾S߈��MP��;�����RC�D{��SSX	��Z�hl���Ѷ�P$Zp��%��N.�&K"~m��x5	V�W���A���֑�\�R�^Ⱥ��W��5��9+���2{�P��X6��������/v��F%;��c��ߨ�����v:!�,����;`ވLm8�$�����(Ъ�i�1`��
[&��;(�V������]�^�O�_H�ҷ4�7�t�*�*q��Q�v�� ]?Z?3�V�.�2݁s����L^�� �W�~U��"��oJQȁ��(���F;�V�hi� /!G��%�r)9g��P,ya0�h/}��*�ܿ�9G�x�&���F���8p5U)������UT�tf��������p�.שܥ�"�ǀG|�3��.�~0ȳ��Í�fӅCv��C{�co�h�$q��d��!�NQ���u���e���s�X�46��CWq�(x�\J�m3���8AzJt��檛:��2������{�ׄ;.fÅ��q�	냄D�{ �Sן�ʎl*S:QA�!�J�#:��r����U��`)��u�@���a�(]l���؁"<"��c�����������+PY[�emH5��:��%��M_���1�9�[u��׳/,iЀ��'�^�l3�0���?�!���i3�a���D���Egs�c`w4e7�����V@х�{��) �C�,F�fe��?{+�"�88)���4�9Я�e������xoq�R�;���L��|��u�)у8h0s������>X�����u�V��C*�$)�y�`Ig�hֽ����%��z�"$��Fz����>�{u��RW�������;��>���ح�$�B+Ϙ���U�7�����ߵ��Z��=liװDm�!ɀ�
�7 q�鼆�}u!�I�O��-9�Z%��N�~�0�m���8��#��M���8`�wB-J1�I����pu(�fO��vk¤uc<�9��u1,\k�_�<)�K��!z+8�qc���,L@bj�g8p��a�1�s�ҷb����>N ��l�eFM�8���(�O�3-�t���6�F�X�f���<���HC؜��oa5�볧�!�R�$�H�A�B����6�����D��j¼��/�|�`~���`vP�0�y@^$�����>����'	���-h�E^�*�!#��Fu��;�qx���^.9Tq�0o��Ό68R���$���! Z�x�.s�~��-(�=6���7�^���G�h�^M���߰���ߘqy�>9��㮦�ܐZ��	P_M���x�9���Ѷa��%u����V�	�ZדP��Uּ�|�a����y:���L|�Wи�"�v둬��b�^6-_�]�3��K�l�����#���ﯵ%�'*�i��p����u�E<g�[�3��E@��C��TA���2�in���[�4X;�duZ7��q�F0x����/]1҄�{�/�`�T��Э�@x��&�m����I���15-[Bv�K�lݟ����N�k�t�O�m��8Z�W$1cYK��=��fC�j��F����YE%�/�y��byNW1㓓�9�F�Jq���x�g�P/`�ҥn�A_���|W�D �j�\T�S������+�@*;q	�@E�[hUsP*�7 �V�
I��aߙ���O�+�H5��3�΋ǵ��?�혲���{rӥz��2,R�"�e�T��	�rj�u��s�A7�ᚉ�?b��*�c��M���Y}���H��L䕟�n/�������T�H�=å,'�T7�tgKr�n��^H�A�#(�������˴��R ����,�O�ôu�6�i�TY i��C;L$�z1i[Ϸ��#e� ��+���X��i��Eڌ��������T,J?��y���8��Y(�W���6�UNY�h5�Hh�J!�z�R��V�p�»�hw�:.�CX4t�1�d�Ϋ~أ괄����ur��$�Id�1�)�ܳ>�#�f��E��CF�홝f	J�2�Q�NE�kܨA������wL�MDpM
����9^۰c�\G�~��.�J�)�nx�&���y?yųlꚺ�'Z��+��o�+��%�0�R�c�6�s�Kt6$-�������eHM�	�V	DA�H�����v���F�~��õ��58'������"��V+A�bP�y�uαS7�*���JU)8S���i��,��9����ǩ�� �=g$AA"�K���F�Z�����S�����<�R�},��h0���ʠ]g��5
	Mn�����賟9G���q�1?�o��� ���\���V��I)q���[���D`��&��w�8�vJdK�6%�Y�w1r&L5�U��&�[�z"�Z,�)�8��H`j�)󧳡)�F�Y�/|�]���tk������^��m���÷L�?����9����Ֆ/�o�	gE�M���Dς�$��ζ�8H�K�+[C|i�fo����4���u��3�N�a{}͟m�CI�`�����m�H	'��8m�
��jv�ǣp�Zd]�׍mJ�m�1Liܱ�2F�_��5�Cpf 1A�C�z�0ڮ����v�J�}��,W�������J��'ޮe�x��r�;��Z}F&򑜱�T�x��}6B����ȷ�JW���{��Bj>G�,�D�.�]�\�,��I���-��,���65��L�yM9t�_�:G��V�6y�X��ەʰۓ��3��(���\�M(	] �)Vl��!	yc�wT��)7rC��xo�ս���:��41��J��2��2���3m�u�3�iȑf�̴o�����b.��%�#w����1�� ����|o�$Ҟ�/~΀�Q��͜yǧ=�(�$p#�L5Pj0ɵ���e�� w�)�FMl����C�-�R���W��7�6X��`����<���cN	+�$<@ff�V�&O��X[�S��Xl��� *�i���$"�83)	Z�{C"@&�a�1v�t�C�Q+[va�q3��l�V0���-0:�sA��o�}����;��ܣ~t�����M?E�xO��uN���4���ˉ?YŠ
 �
s{��a�Y��ϟHM
��앩j�_��-���,]�Z}X��Rz�9?|ƨՈ?	��i⇘�����w?�П�?�8�8֦=��ʯ�Ӄ�/�j�]���j"���}��\�����_�����?9]yp��&���a�b��-[f\e��;A:M��hР�>�Ts�����N�_��Y�$�g&i� Lo�ǅ��}�����D�Z��Zr��P$��b~��Sr+�I�POI�e;	���{j��D}�@��y���	�/Bvr��dfqR�j:�	�2٧Q>%��W�s��hsL��x~Fjg�	DoH�f� n�YŸ���l��H�L��584L�u�TA��ԕ;Ӿ7Iʋs(Ӱ��p(��+u�{�rG������U���9�V��Z�$u�A:#�}������9v��Ǒ얗�i�;6�h�j��<�41F�X�AQ�k>P����a�Ew!�u��	E�8iVf���91dVσ�����W.��*4����&E>&w�3��b�Kz�����֙q�C�I�\�?Ӝ��+����l�*��@���I��\�+��������ޢb�exv򡂳�H\������G�}A��������ۇ����s�}�'�HD��nA�1n��z�dm��
b��9P�^�S�n��]�����:��A*<�y�>ţ1VTD���Ȝ=K��t�F�'=1l����✸DtG�Ͱ{Z��x�ѐ��|���Ɏa��� �2�+~�Ƨl1Y���]�'MjU����v/m�cڊF�d���;��Y���^�.���&i��z,㾼j��#��!��t�?�UB7�>�v���>a��~���a�dg��Lƥ�㨮�5`<��B�T���Ôl�g͟;�J	Jk)��=�05�`��up�,ߎ5*�c���)tTx�h�·t`Y75� ��� ����c0c��X�g ��E�ԩ��ݙ�`�����5��G�+���Ҁ��Jl�8&�L�ܰp.Zfʓ��Q��)�7V;MV��c,�[�:]ˤ��z�1�XJfx���۲��r��{�%�)��� {������×8�-ܔq0W�9l�C��d�3�
c����&S�r�1�t9"��v�5ئ|X����J=S���C��y�HiR�����6�|���i��hq�)�~V��Ȯoм����G��P�dӻ���5�틩}n�Z�uHG':i��wہ�!����*����!� ����or����>��|H�g��
�x���/�Tl��f�:����A^�����)馟��b�A��
�]�s9�q\�D��F�����eMJ�{٭�ƃYg��z�K�`�^$�4��?�H 4nP^5=s��d�(3y���@�ZZ^�i��[���Q��	F�P��#�����Z�	t_�#�/���z Nf�h(L��Ё?�9QI;���{i*7AWo�p~��Π�w�{�h��p�f��f�k8C�!Ō�G�7(�03�2�-�Ȝ$h��X��E�z4(&�C-oQ�w".����9�3���_�o�)���/$%ŧ
A���^>�	9ԯ|��x�����[��r~�
���cTw�l��DC��K�9V���T�����w�e�,�O��P�R.�JV�XԆ ?���<��/�`���] �,Xp�Q]k�&V�8f�˘�'y� 4�C\�4���ז�����k�����m�m���I�G�u��ZNCX�`d��c�\!�����"y��e���gnA�Q�&�5W�5�!�u�6���R�bo�����~����6�s��B(��t-]΀�i1��t� &�Bs�ø96���$˲_�/����9˻�w>eS� =W�_so�S�&iQuSW��͇�t3}��\"��6y���e���5G/�w�ښlL#CU7�u� ��)�%!h`��/PN���.��Y��o�拝����	�O@�F�:�^6�ƹ�[�*T����D0���L��1� �Zq-�x�W�J�uf��j���6F��C��-C{61�oN�N�s������ނ�u},�ǈ�ǖ������ ��c$ʞ��z�Cc2^���@l��/�8
5p��=�8�k�,KZg�m�jcE��(��^��~ Qj��*�v�@���.��>�H(�=��$]����U+^_�
<��b�7��^���XV`pg�Ҭ��V*��H��R3�|Ҧ�c�X�F��q�V�b�d�SL=�\��;�W4� ��T�XT*"�|m�Q��c��:�z��^��~R�Ug����`�^�>�Uw`J��X��kL��imԊ�O��J��	�#��l�����K��0�O�J�j���
��%��NU	��B���]�V��[�NFOv>OU�+�������Mû���B?�9�Z���nV����*2�� B�v��ڧ;��A3������'	��3���<��;5�+l�+��p�mh�W)�0�"Ј�+)<<|@�A���Z�4�lv㗏���:�cu��?���':jJ��CEd�^l2&����xp��q��l4V���'M��в&%�g;n����|��vF�Pj򠿻�_�+"f���n^6b^���`6���@(,�ff�!f�韵�fg5���6�����������9�JhL�}K\��h��$�����-���%�CuU���uT��b��B�������I���x��S�~2B�����aX���V)?��.�hEŔ�����x��-SO�Kж����O�(H��R�OQy�ne�T��l4)�őW�n�:�d�A���0{�:��=��h#X�?���k�ATƣ�+�!w�Oӌ.D-`d���������Y�A��6&���V��U7l�rX���.m$yy��M��85]$QNDV���D~�8[
m����E�"1�u�6�����v�]tv�x��1p���y܇��p�H=5i�Q"����H�����X{��׼���V��Z����雚Og�O����sg/�j����|��h��2�SP:MW���]R��z�?<��!N,��7�tq��,�֏d�R��7���Ğ�Ŝ�����}��jSr��a������ui=3�w�1�}�g�t��WE��w�wZ��=�P��xu��}�օp��F��'��m[T!Y�����xZȸ��\��@pnǙusi���aa��m�A؈��4-n�[�;�y�L#����������2xa\Nob�G�\fOԺU�\i>�P�^ȃ�|_Ac]н����NS�^�L�����&>�?��E�0�ORxD�	R�A{uD�#��:���|�aU���`�W+ʮ��n�${^�8� {��X�D�V��u�E]Hrϫx��}Un�
WV@^p\�9�q\��u���Ta�U�>��AdV"k!Ȅ4Һ=Ѵs��Hkm���|���UD����;6%�Lr�[k4Z�F��q;lB�5MY<���@��\*w�E j����K�a��iq���T����u?��{hK���KU��-úR�1����\a|/�qj��bfW�Ę�%\2@	��l�E��L�n^�j����7c��heC�,u�b��
3�pv����m���6I%va*�`ތ�I�j���z��;���g T~D��X��R�ŉ:����Ϧ�묖#�R�Ls��<�Mt�Tb���Hk�j���P�<�ge��]��
��)�Ԕ�\�����U:X�W%�p�Mthbφ��9��x,V �v��ʎ�{��y^qI[{G�/<�Y��Q�xdrYl��Rs+��������o�?���xE�X"M0Xส��p\p4�7�EB!�$)��x�7I�?H1�kui/���Ȭ�0�� ��!��_&��e!�����/��[�8Ȃ�(��`�x"p=R!��O�^b<��1�.�{�q��7%���

���Nw�Hy��Ah�h�^N �`��#�`�m?�ب����¬)��Y�ud� �q�����-�`[���'S�9�i�P��-��ӽ��:v��TX��E����|��5��D��l�y���ׯ�p�~
�
,�������BA$�k%߃�gi|.�i#����^e�tB2Ru�p})um�����Q��YT�o!�*�ܷ�������)İ�V' �s�v���B<4:Ï�3��e �U��z�g�DB1�@F6����� sPRE8�$�Ȧ�C��M؞X�v��E�Nv(C�^1	�r2EKZ���ITm���7K��/�� ���`�M8�u=s��9��	��s��Q�^�xI�O+*xk�R�۳���hE,�h<�bօo�5B��N݀�89A�V4�%R#��5¿��I����^l�\s
*ij'/�hכ�>���#!�g����qyv���`����>�m�=�vjӥ#N�V&:����G��L��Q�#�50"] ?t@��p����H/vTĦu��Y��ZӚ���3Q��S�f�k.vͽ�}�Y<S�� Te{�����M@N�#F��}��r\��,�\�K�a>���(����	�oˢV��Ya,�W�j.=\���~v4d�Nܪb�0a�W��(O�Z�cx��Ք��RhK0<����m�B���GU��k�T�շP�8�"a�C.+��Uh�!�Q��;F̯=�0���)â��ڤ���A�t�};0n�*̒_D)q���՚Ȼ����sE��:":D�Q6OZx�K?�b�%��^C�ߊE��Xe��Y����'��<@����;H:���.��)ƿp[�B�;cMF�5!>����
�޹J����@ޢY�t�\��ҽ/��DUQlG�I�Ң�?��2z�X�T��m�����+��`9�+5���ܪ�L���c1�n:Db�n�y��+���n�M�#��V �я���B[T�V�/�&���k�1���$K�l� �jPl���IY��ݫC'���[(~�]�y'���JF*&^qm���W2~�!4� �}�[���H>����^���]��n�)�U~�P��P *Z����n�f��%�r3�L
/U��������:.j{�@�~f�\�.+r�x0��	{К���j�-h鑝x,>�w�&����<��4�CcW(MU�ы���,�F��_T���H�:�+` [Y�r�NA�j��kobws�����ڳy(��P��Y�2���X#�t�D�Bu��E�#'N�mTV�nSx*���P�V #/\u��+��iK%�C)���?&��?�}rb�Cu$���ˤ9L���PAZ�ʏr�|SL>᫳&�Ю��=+��c���y�cȾ�|�aOg����XV��|_,�����T��x�Q���?�Z|���׊��~ZmO�W���I��Y���c�y1cA]�c�)��� ЍV� fȹ��$�^O�&�9Q�b�pߖ
��4�*嫫����H[�� Xɾ���/�CD����tiD��2��G�\S�v�y����1�qh����I�=�s����<��R�V!'�>|{b���u$o�c��R�|i��kњ�� c�¿�D2����P_B�D��覙:�����.օLk�3h�J�=#�y�p_Z �#D�lS�r0�f��ٹ����-��_��y��Tt�Րo0W'� �Gw�hI%eJ�����pj��m�s+ocU��o@_�J��8XTR9
=ˤi��1i�=D�h��	 6��zF�ɳ�N�Z���q���W�P;�x��WS�p�?�aշ�)�z<��V^_᭱�O:
�\{N��jܔ��rw� ���X�����B�|2Ѐ����Db�Y�5?��X���#
#����ilz<9:Eu�_�����<�[!4��_�֘7%��M�����Rm����8ӽ-7q&L�P8y���|��Eٕ��ݟ���N�%~�n��[s�^���.j�7{�����R�z0��n`���6؃�G�����M��\����=���W���~��.�VB����x�٠t���(��4'Oz�R�Lf���eW�	���������R�ֹ�׌*�B{�Ɏ���}�~	f�<�T9<W��"�ؤ��i��Uh����D^̛�z���e+�$�����+W����?uyFۢ���N#R�l��<;����g}D����!�s�CacrP�=�rlr0L�:~����.	���_Ƌ���^t X��.�А�v�l�.N=�!J)R��1�r��;������� �4�r�q�ɽ=𘍙F0+[�j�����	)Q�F�-!*�t�w�ILə⫻�£�V��t�d���ذǑ������W�U[�����ʕ` 2^w"�f�+��$�h����ZھflTdz�KT���v���'�~ݷ�+��B1���b<�fW�딠|���Q�EMMS�Գ���Ś��W��j�3�NbpE��_б#l�BjW�1��>G�}'#w Uk��oZ�(4R�.$n��̢�������̟@�3���1�8�A, ��>���@�3���oג;�A�}{1��tzx��	¶L�G��1|Ik��Vg3�K���m�,���N�h�^�Aޘ"V���, �"��,�9����Ð�+N8�:$Bi�r��f�H�{�W�v�;�V����;�k+d-��� C���s�Ó^�f�K%�7�g�N�5u���׊(vV>aԛhkOt��T��8��Q�Y�g̊�*���B��5�;�?{�'�I�kdo !���\|��~��+>�|�q<���S��<���7�6vu*[Щ��i�M��[g�u��;o~�le�N�ڳ�s�Z+��Nh��3hhV~N�b���-+���:q����(���f��Ƣ>��3�SR�&����	��[��.Dl] �yۊZ�:ǣۃ�Xu��cB��^��+�A��la���bK����tX��g	7
���OX�bn��*t���@�у����>Y�ڃK�$�2s����d�H���,��W:9#�u��������S�#� ���*2��Gr���p��@9$�&|��ͺ���{�"(��Ӟ�/�)ԅ�ED�v�*��-L��8��w��^M�̒���gt���.���og'H�k���*�y����G��d��#\�r B k,��j1��	��zc��ʃ���N[iyM�4)��ǹ&Ҥ����'������0���_�k����֔��2�G{���\�,���f�
�ҳܬ�i��ZC����og����^ɝ���>��
��V[8g�̽�����J�uG�ˋS�Hۯn'�p�n�������bl�LY�%�-�&�����w-�c��1 gh�=r��z���7Jَ}�c�"c]u:����o:��co `�a�`�%aBF%� �*�Z����'��kf2�Ll){Ja����d\��kbk*� �D!��ye��sF��>�_�~N����{��RD���ެ�\���f���l+)�G遉���Ej9R1��X��L-2 <+������:n^�70D�]2�K@H�#~\�����Ty��X=N{��dG;��}ͫ��=�������J�-ȨP�J	L8����,
��t������׾w��+���,��Tc�4|3��~,e�,@�<5�1�^9K3k�����'L�xR���B�m����b3�d�˶~_8	�Zq�}9�t$/b� )����^� �F��Q0�-o�	LC4	��"��W.�4�1"71�B��=�$*~���O���'.�$9vě�����F)�/�f.��9�r��9���p�=kǿ�rບx1޿i-�m:�q"�d8pڵP��	p��X��2�A?�]�/�4�j��)(������9�x����Yم�!P�̜7�8�b&\�W��',����ؘ��H�5y8.f��Zҁ(��\��t�td����GY(1	�5/q#�ء�@5��XX7>��l��T����R��Mj؞^��]�"�h	�)�`7a($���B��z���-��;+]��No�c�tԡ	9�&���>*�2f<��#�qx��Ë��%0�ȆeWk��!G�+�S�A�C��I�wN�q��Ϻs�r0q8���g1m`�59��;m���6+�'v�(#J	���Z���-Q#���!��L�{���n�̞eoq���##�Ʒ,��0O���3�m=�U`Yv�0bG��샗�\�b��d�[^�����>�Akl���k�OU�@i��q��j�w�=���1���X��OJVҨ���<~r%��![���s"]C<�s���1��~�/��l, �Vu��e20��h1Ɨ�����o��G�ƜK�V�3���r��8�拾(�����'��+�i�������@uu��m��ڷO츹�N��	΄k�B[%@�C��a��f�w�{*����1��TH15���*[�����/AhJ!68ܟ_6�[	X�tB���k����v�RЈ�����[�@~�1�+Xr7�ط$�2}���*C2I��m��S.�:Yǯeo��Z�R��{�@O�yJ���#~�e����g7䖶Te�rY3����Ho�M�� tA��c���r�� A�˾%&I`t�Ô�I�:",)-�|�0��u����P'�X�*?P}�9�D�(�u���;��g5�f�+b�P�:��~_��>	�@�-�g��ܤSn����궇�"�ǫ9%�,�-g�\�)�^��Ɋ�ѐ�@���7�x����bK���V��$�4K���7-���"���3����]ݜ����$�q��
���~1�R�g�kw�����
<#Z���%��,ؒڠ�]��+��y����t���vxB���i�%�-h��>��1�(H��p��:�h�d�x>:���c:�= m��||Zva�Y)7轐��i�A E�[�'VZ�mp>���T�H����!ĭ�Y��^�o"G-*� ;ua�ք�_��5"6UJҷ	�XG�nm�.���1�q��x�Y���9kj�S�:��a �Ѱ_�[u�MS~��f��,�r������Q��BA�����8W����W�Q�����E���#O6k�8[S�O��Eb}��D�A�����da9z��+�}����Y��R����v!���#�o�̚l��#c>`��*�qh����������|u9�0�	н�*A�).�F=y��s��%&E���᫢wX�q�u�C��w�uTRf��}��\L5/�M_�F�"�]yF�������+耜f�,v���n�$E謹�Y\	٢
Ċ{/"��2+���`h�9͟�	D_�Nj�^5�ǁ��8�k�Y�͊J:�R��8�8��w�	�1+7�/�")�$�`G��g!Iִ`�X�6��4�]�̰�P,xh��_|a�d�t�&�V��T]~Q2�H�MW8��^���s��_��y�?�:l����ؘ
��\�Q�vd\ f���"�F���T���rW^���
>�'O��Y����]w��}/{�4b\�\�m|������_KƳo��V�#'�T�H7i�{I�ˢ�4b��a98��˸���u@%�����K�#Q�-U�z�����ϴzo�iD�X �yg.��<`ݩ�|i>��HdwGcA>ܪ���,���ds-G"7aS5\wd��X.�r�_o,jn��B����� �Dg;���^�u����<�/����ψ�#�3�_V� ��o����b��fLˠ`��(�`1A>��G��Lz_6||D�-���j�%C�!YȤ��5��v�6D(�?��V.�rg��Y\�ۭ��hd;�c�%-�Ͷ����r�N>���[�F�[������&��΅�?�����ΘCz�]
�1�&BK�^�!��O����ɑ�I��)�js�R�%D��o����a��ly����3�L���c�	>s6�t�1���J�m�=����q�ċ���Z�$SwU��}�_�h~���y�	�^;���>]Y|�O�G�@�j�V���N�4jj�>+���-p�r�v�.�5\0U
`��q�7�O�W�*p�3*n��S9\�V���z�K~���-r}i�i����/n*��k�t��EB$ƻ���;g-�#�������C-@^�ɠ��6�b̬R�������'��� �����wΊ��3� �`�n7�����I-q�2���U7��O�Y��b�[vȷA��RS��-���xN�����T<� �L�tp�B�/�Y.�޵�v�f#��afG^֗;�z�|�Wh�g�h���Z+G���YύM��T�2DD�A���7k̟_���p�rV5�,��XJkX�"i(�񶻮i�-��@~�A��a�T8�ik�X�����N�éG��nG��q��ֶ��03e�4�s>�i߬G�Ýk���M�>Fk��֥�_]>�H�ȑ���\���,C�����}�\������Z/]6gGgg�VuVn����e	Պ�L*�v_<��,�+%���9݇��X�3���c�PP��[���:sZ�w�.~n�m?���u�azk�1�i�3t�vBA��i�v5��X��?jvk�U9^��}��g5������gө��ND$�o3gK�\B_��{�*�K�������#�Ƴ`��O��#B7V���w�@�YA���1S��"��>ߑt��J�ݬP�ن��x�ƽzA�ʉ�v�e���=�)�⿯s�"�yi�R��{-`���q�JW��EzO</�[��?�$�a�#�;g��uw�1#$�N�гm��FJ��JO#[N7����7��{��i�x��UynF󂼽W@�η��ɨ_5��)���
v��ڠnv��9�e��dn�G��c���Ī�ֳ�y'��H�MҪ�^�7C(�eWum3,-B�yl �w�rW(����H!*���|9�@���5���>�]Eo�v�-���6�E��>l�K�ez�PkһcW���kf��io�%��c�EIx}�;U$�Ƙ;+��D�a+�L@����D}���A�,���<�ȒKY��^tc�{ܼ	�î�u>��#G��T0�8Hߺ}VUћi��'I5m":xX>�HSN��ۢ��S(��>�y�v)tLFi��v=~��*6���U&�.މ3�~���U��`�_��	�(��p	�g3�]�=��5'_��3�L����Wd�� �G~i�3��'��ZUL1wEE����<ڇ����PY�&�J̎�`� �rU}i���̍϶(C��C$V��.�F]��ȁ�R�'zb��Sa��b�B�M�����xx[�+1%��N��i3�QPph����q�[70I����"-�f��^�c.�j����ğ�̡��<������ѡ�i�܈���2�7�m�m��KYHEp�)z�#�k	_�Z#�3��t��}�ڡH�!�+�Q�>��観4"P���
�(� �B�&��ݴi��N4�24Ëd����gɜ���[������("��3����R��R-�p���	�L-�����L��E�[mIj^������>m���
��%�w��Uh�>R�5'�&R���u�PBb�f	�͖����{n▪���*�Q�.�Cمi^D<E�Z8�h�$VϏ�v��Jr��O�'�"��S�Ԋ8c�ˡ?��1��:�|d��z�,A7����."4ZߕvI������B���π�k�}'??l���N�Gf�a0�)O%ɇ̫9|1� ֛ˇ����������;��- 4vu�H��p�f��4AD���!I�il-G��'�����KJ�����]��r��+�T�|�t��qL�L)��w��p`&�G�C�]�xA����}5�&r�.�S�QQ��a
���>�L?�&��Ͼ��Sܸ&=:�pgoJ\E7+�sl����2�Z�p_�gB8DJ���3)��)�Ҿ�:�иu�(E˩E_X�T�P�4�[�a��1�F�R9�4Ģ�&,'���-���0������p|���,��p>`�U�_�m��c�����չ��@&|9�cŗ`�݄ߨ�-Ў��q{|��zJ������o"�5��ĹoN4
��A���c:W�38����0�:ᦧ{��,�X��U����V�=������ KvS�B���rg3�����{��ו��vI�)�dgf����[�c��EV��kt��ih�_F�	)o��w_Z�6����cN��F�̍�́6�̆���|�@Tn�L�u��0:�=ݣj�Ըe�(>�&�e���5�����dW�&���G�{���э���=����wL���2��#��37�򙗁�W���,�z�G��1�	�_��4��6sI,|hK��sA��#Z�[I}4šư�=-bտU���#�L��Ϗ�H�_�R�cI�y�+-�q@��/�����F�w nF�\��-4-�<ne����x�XI>�����+�4UeC[�^fh��t$�n��Ӓ��R�̫Ҋ�B*׫���QF����M�e� �6*��^F���
�K����T�4��&^/�z�	�ܤ��S�ٳP�V7�fpT�^)sf����� ��W�?�ٿ����57]�g�g����&�G�j4{�{��*�5�I(d��y���Mk���8`�P-�97/&��I��.�KUّ�Њ��6%�{�]l��(4������	�-���AxOyF�/�_a�#YU���W�^�}O{�_�n'�gmc��o��i+��i��óI�kx�m/�K���=�w$��C&�����ke�6<�+���IQ-����C�5��#��Q�]�Wi�M'�YZۊ��;-�L��bl�\��V��$`�H��/�)�ɫRG��U����\$�(�KH�����{FxQi�$S�+;�� ��E^�f.�:������K����˒��wyF|I�-�`�u�dg(�n*׵u}�+d]B�w�Y�W�w����K�.PgTRp���[ Q״���%{m��$)G�g�Lɟ�ϡ��,1��ǚ���+��u Ȱ���Đ�r�%w�|8��ل��ͥ	�n���e
�����	Q�C��a"@�_�1�5O�3Q��3fb�<RD
���b�ޠ'1���>ik.{�;3�*%}	�&�*՛��+�B�o�;�H����Xu��J���7JӞN����Brr��w5و�����u��� �2�|�ڙ.;cb#�M|i��X�����n%'�zB�`����h$�
t';u+��q���K4���>��3�����7����C$�jK��D���'o]��,(C
�׫;�Ԯ��XK�f�T%i��h�Ts�\�bJ�"Jޡ� ���fS�뛒��s�e��_�������"���Bk_��;�����!#��8'�[=�D�,�C9����I��!�����R���:�5e�t��r�zt?�U���-�98���!�r�\.z1c1��"�XL�S�rB��ۑ����'�P�S��i��-�HM��r.ꖣ;4e�dӬ�X�4�9P�^��&8P�����|�:�R������'�.3��k7p���my�o����n�=Ԗ3�H�ޥB���*�l�) ����d�:�Hf[�ġeŶ�3D�Yy���뉙��6�~%?X�������mv}�x1F�WP��l��Ȩ�y���y�W�5n@��H�A-G���
���h���UhvT
'��f7���1�]<�EJ�x�CNpɋ�p&��D�<�n������VČ�2~XdH�#�L7ˢ�3���E�F�k��j�ȨN?)�(��
$���_Y��x�:����Lns��z�.�o@v<t�b6K	*�5�6���h�?1���'�(��Zg�i����擼L$xâ����=��� q�NA���h�sGix�N�^t8�#T���	���J��l���Od�y�A��YE�Ŗ�B��ݏ.�{��P�dB+S�(w����e��b�=�d�ӊ+��:	�c�)�1�*�~��#�Gp�Zw4�03�^{s2�/�����r�F��`=;L�9�	�.��*�.�V�ܣs���Zŀ�u0��(�se���P��̥���
��.�W�|s�deGSBhF���� ��h��X�;�RSsA\F�:d����(:��>���=�,��,Lk��U�MϜ!N��i�)>X�R<�되�`(���VT����Z�oF�s��𷡙�Ev��P)���q�C�laަ�pne�=�7���G_9󱕠C����mov�~{�v\��4���fA_��.�g'��:��t2����a����&���;l)�Hz�2���_�{��V�£�W�_څa.{�C�� ���(�� M�+%�B@K���� :b��εW��;~T�/߫�h�Sd?��ղJ�g@)&[Y���I1Z�(0�s��}c�V��0����^/�c+�я�5���x�W��E��6]Z�8�l��LĭI�yAɗ!Cq������%�u᫮^����mV_7�W��j��u�B m��?�uP��J/C��&��3h���R Z�C�c i'��%d������Z���xl����H)��g[[���a�T���M�~���7!'�xˤS0"m��Fc�О�}�^9�g�o�'�N�(�m�a�Q�J9�w��*��J=�$�SM�{z���/Y:�r%�[�|���fw<��F>������:�r�Kwܔ�d���@�l�di�k#pp��N��i#���e.��b���2�}[���jF�{����Y3����(����W�c,2QMB ��r�w������>C�W?7Y5,�^�����	�?*ԑ��=t�R�}e��jIgi�#P�	-�"��0���`�y��_��ĕԘ�|x�c�+�G�\���A�/�,]vUY����J`����o���M�( )H����]y�p/��ؤ�N�;���U*`iq��ϬU�wzcO�����3���a�3��$RW���V���@&뤻�O!d� 5{���x�t�hi�Ʋ�-�SП|�}ma�Dĥ��:����P/;���n>������(���c��M�tt>�I=95���k��PC����5���5�FQ� m������dn�Pe�o�����`PԮZ(���!�*�m����~��io�KW�J}���$d!���0� Y�Kp�v�k��N�Mc/���SG!�L"�����K��J(���1{���
��=�(­��V�����><��э��ڗl��C-�v�AE�|Ϛ��\*�E=�����tt�W�w�0
��&=�īM�8e����N�������T�?J�����E�� ��?������s�(�|b5����LU���ZШ���og]PZ�{C���e6m[+�iU�$f���)�?�AW�J�?i���"����	�� * �o?�"m�*�ƦgKg&?m�tP�i~���=��X�����W�߶W`̀�򉛛��ym�k��*dn��+<$����(LDT�T�y���H���D:$��*/i�Jٞ��Hh\T�����&�E]p0�.�B�vd�̏�F�*�����Q�Ԣ��1�Q!���	y�p��U���"�֑r::�4L�|5x���60GԠ�0��zk|:室X���v�ƍNT��<��\���A�Q�����p��R�%�*�~����-U�/�(�^��č���ndB��勏�HI>c�͗�͛=���MKHr�6��z�,��.E�F���pO�j:榳���X����~��>��1�g�2���#B_�a���b_��5N�_�; �|h�91�v`TsY@�ԊN�ux/��{,�(!6��22V��4��<ը7�Fmt�JR3�^D��"~\����0m�0 �^�����yt@;�M6��(�+��i��\�U���g|������bu���W�!We�!��
+�st��r��iD��\��pO��}�����)�=�V�w3ޔSAҋ��~Nݵ��F�!J���nI�~� ʐ��6�[���rpv<5�v<�Bd��+-���/����reV�oˇ"kl� y���7`�A�vH�ɡP����\R"kh�Q3�J�����8��K�S�^5��<�N!N3]�mۯb<h)b�>�Ҙ��%���*2	�7v���*��/����v*��b�	�𢡡���Z1�F�9g���� �z�[9o0D?nJ�]_F�qN?%B�餣q����|�A~�t"͇~%{�ްj�I���d�)u���1��~۫����Yp5��M���Ŵ�.�I���@��Ă��L:�_�v�ȑ:m�Ĭ5��
H��O�
v���y<j��~{;��5�a�l,�� ������:x'SrF#��~�t�\�M�!����Z�` _(�y'�a��^�������t
gZW#Q�H?��:!��jE��HS���NC:�wWL����wF)������mVj4��*t���sb�X���/S�lq.�HT���}@��E�E�1��h�~_b���f(��[ܐ��Ρ���.��k�_lq"���dkɃE�R�(��+��j�n�`Xse
����!��i^F##":�\���rIy�����~'����U�+�s�C��&: &؎�;�`��v���txo��nl;+ ���@���/��I��F���E�G�{�1ժǦG���mHIr�ƈ���+f~�[��o�+���F�L��i�|kk�A_�2�Y���zk�g<��z�ý^{�]�	��b��h��\��~����2c��)\L �\i�8&ѴE�z���h�g?w�{�3>Q���-��g���o��p&��+�~��R�7��
?�B���d����K�����`���l��_��]�{t S�cu�$���B<�|ܔm��%��$�����V���v��r8U{!����m��z5 0X�뻈���;f�ݒ��;s�d����^��.�f�`�`���!(��ޒ59`�S�ڀ&-����.hM�+�%�KLe�-�%��ދ�΢s+Tbv9+w��"�����]��񷫉��l�����XUF>����,����F�cO3< L���p�l?��=~��C>1�n��K�U����,�a�b�9$l��v�� v��+���l�jj�g�~S�p��2��X~���y�ڍ�f ֓�o'i_�U��q�,VC2��K�Rdp�?"��b��\L1>� }fc:ȶڼm�m;&�D�C�9�'o_k)2�VV��,}d7���)��A`�����yl2��Q/��p�{�Q��K{�_�}aI�#�JS��l��>��!�F�U(�w��{PyT^��aͼ�	�#������jׄ�0t�>�&�c�3}�{#�{�AF�O�^�|���h"�������_��ǿ��$���#c�9���Ӯ��`�
P"��|n���(ۘ?I��Ǚ�7O�ԭE��e��7i��xۨ')�TW�<'��W�k%�̷���E�Z��?T�ثÊ�֥ �G�8�bǽy�h��ܴ�{D���P�I����� b�T�\���|{Yט꒾"<�9��mCz�J��� �3�б?�^;�?}S��ntD����y����._��uZX��ʝM���M�S��B���:9�O� ;l��o9��sow���qLf/+ϗts�s<!a����	�ہ������������׆���]u��
�F"��oV���Y�a��M����� �zy6�Ԣ�Y=[�t3aSF�/udϐ*cH�8�}�X伣�ߍ"�eid��IAn$"kT��{Ė�L�%�h�?�D�'-��c�Q�8J���w����-,Bh�ĚV�������}}E8mTs\��ሁ�L�I��~�@G�H}���>��ȹ�~�<uѵWXG�9�Q�z	XeZu��)؂� ���|IP|���ٝ�k���)a�O}A�r���� ����5
o��Ҽ36�U����dP2�V3^a�K�4�q|���0tYv<r�2g=Jcw�m5��ʷ4x�d;Xz	jǂnwnQX�g�j�d���������	̽1��:L��pI�z*�g�v~���eZ��Nqg��9c�X �;�W ��"K�}�Y����)O��N�␁*�Gii�ŧ��+��LC��߱��_����)1S��활�}�@;e���c��'2���J$�-��F��{�!X<f�'Y�p+1bؖ�qnY�Nǁ
�[���eN�+Gs �
bˎ��#��A��m��ac6�=�����P��G9&њ���*a+��2@�� �[�0�xۿd����#��z�l�]���g0���S��#�u��U�D��L;[�ZT�@�w����P�����=�;_&� ���4S�S����V���$��wAx����7���G��y��Q�ӹHůȢ��"���9�Q�y���WB�������pE�*�b���(��5Cqy�X�)Ct�p' X�G*N|�j< �$��E��|�-��)���W�J�(��Ȍ�$�\�eI�%"��/��Fu}�����O��V��L	W�6�O��~�m5ܖCz��~�RK)~[�y�s�6�BoGQQ,#�2}(D�p+����T?*�R?��:�rl���tbYL��1��2�>��ɕ�N��^ؔC��m N+Z���l����1b� t���H�-����}2Q�Ծj���h��,��;%W(�q�L���U�~G!'�k0���?�*x �ꘐ%�/�-0�E��
�CW �ł\a6�+�Ϭv�i�Q�('�@�u��lY�݆��[�R�w���m�P䚋�I�;�����U��zn�~Y�^��������-#����L��m�Fr��n_���9�X�%.�"�t>@������*d�mD��D����sM}�o���XF=���0j�@�T�h�͕�.7��
���/r��m�F���w�=�=ق�$�n=����uY}d,�X���0����nuh�3���Qe�&c5�z�o�%'��<����󙰊4�I����c�8�"q8���QK?��8�>�Ms$������qw�i���L`r�?����o���2����C��&\��S�_�8�A�U����t���坥uB}�J�J&��ԝ���I�|5���FJ�jQQ/'e&�<H�)��
4S V�dǃ?7c��馓�