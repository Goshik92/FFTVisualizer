��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5o�h?\bv������Zr]�M�wM��a!��6���R�}���h���ƺ{K5I�*�q�p~"^g�3��j���;�ul��:m>s_`�i��wi��2������hL��ۭu�+U�u�.R��_�o���%�t�|�H-�*��I��x���yiI��`�iJk��B���e����O6��k��;�q_�׆�Y+�M���´}��E7!��J�Ż���p��_U띕Pݻ@�݅'"`&�1�`t�z��yE�W�z�Ͱ�NBi�YJ���VM���T�y�f�rf̟	�-M{�>!:D�N�9��!ċ��A(�j8����n[	��W�u#kNn�.0��$�Gݿ?&i�h����0�g�kq1�;���;���D�,]*Z���3�>YɬK��w�c�hx�]�B�d��ۈ�b���Y�C�.�e[�芬%!-�~�Xa7��ؤ=��7X���q���z�(��Q�P
�!_m
��"y�%��z���^�PS��N�T;������o�C$��No�qP75a�yHp.=su]�B^��9�u�oP���Y�VƎg�嬧���^ʑW+�C�BW�52K�?$#j�PXƝ�LGG�c�B�V�s��l�$J����*���1����h� J'HUg�|��P�������M�{@.YT�Jb�#�Bѓ�refU!�7��A!P-�O�Yx,5�u���N�Cي$#���v�հ��.A|:��Ec�-an����!������^�,3�"��ӳMp�T�֜K�� �#��/~�� �gvWRl�L�c��l�\Y�Z�'��R�"�>�<^���?�/3���c�_�]�EP#YDc����5@'�/��r-L�������^e��pH��G ���3vO�)��Mx�ܞT�z̀�#`�Ye}�8���c%�{����0]��������'��Ӡ�sY��6��H���܁ʓ �6�p�,�L�/K׉�׿��&9�y�ޥ�U���n�0����x^�����4ͧ��$��c��׼� ��n@~�G���P ��BRT�9BPj^V>y�,k�����$�tY:���j���fbX� ½�]Fx<�"�p��(��)�g�w� G�����=�´������d�(��jD�i�D0�]�To��&++N]u��dE����^C�1jQv
�%1�&�08�[�9�8������C�"K�p%��7{ξRo����+�e=��V�j"i��������Fӭ�Y� ��Fi7� �b�!*}U.�̑�k��+͗IsD��~���(yd���IB�yq�' _�F��p�0\�x�@���~��H�Q� ����V ��#���a��-��<U-쪄ڏ��<�QRj%����K�\����H�q�6�P�������/uR�������*6N�0�Yl�E+J��]%��o|������᭶���[�-�<�(�(�Ѭ.�N�Vӡ�-�r��
�Y�7}$�#<������} KT<�z��P�1�r�\�/�t߰�8��~��CI�~xPRPV%�V��*��@ܔu���8�t�����{���P��bVxwޣ{��
/ϼI�
��M�Z	�cY>��v(������.��r}x)��B�7��y�?To0ߣ��9��4�b��2-)iS�iO�\��3Ԡ����A�:-FsV���`��q�;�����pA�%�V��:9�
�k����3�J��=���A�����"��ٔ*
� b|#��]
0o�u}Ɠ�tݕ��1w�a��GG{��}���zԣFb��&
�j)�0���a����힕�Ҙƭ�{:CU�Ox�H�эO�m��^ʊ�ه������qP�D ���'�����kQ���Z!7�����9;��X.���xa�zvqp֜��	�}����C[��8.	N"�unJ��`bO�yw@PR�Ҥ�Zz��C��B4B�~۴�
�y��ހ�>�z啚̊;.���hS�i�1��N���[-1��)�8�(�C�V�2��E�n�\��l��r4>��D�nh��^Z�5_dzJ�}���y��oA@��a4�p3<�D�+Uo\�+��O�YP��q�,�Yj��0��x*�)U���
��H]ҖaM���L�|�kX� -�7؅���]*J����$t�g�����!�*�G(������7-�C>�ћٲuB�	�RbN�hDau���ǩէ7��S��҃��h1��d_E�������isd}@�g9cSӕ�d@��ݷ`�_�����;�g�Eh��E�����93�D�s9�/gC�5�~�}@�H䄭��kLsy�Mܘ_u]���kv|�l�A+�S��\(Z�i&Y�@�6�Hzغ��
�'D1W���X�tb��4|�2[�Pk�!\+�i�Y��q�3���Vxl��݁���~�Ъ������qg��`�4��T�."o|�]�:85i�`����M�)��\8�4ȗ�g) � ������z7B��V"�QM�ӶƓ���n(�Z���f��G'�� ;Z
Ɯ0�~R��T��o�o�r|r��W���V������ �e����X����K�"��Gt�QVD����l�3�w����&}�;}�~.����Usc_e��\S�S1MX���S��}p�Qɨ )OQ�~�b�]ʳ85��Q�,n��<��(X���'KO=L}BY��~�Y$�4�e�G%n�N�~�"4H;{b��̂��>�CN���wf�Ǌ�
��\_[z-$� d�ek��4ɪ��(�e
` j�E�P4�?���hB��Lu����;�����OBo�MRmq�=5n$ռ�x���Dr�M���l4��{X�Y��|�5!J�O�y�O,�J��Mb|�(p�����2*DePu���e����WB�0��B\a��e�b>'@_����Mew������)���c���`w��S�E����&���ּ0u%b�Aiyh��n�GL�N�?��aJ���8�|Z���(��[e}6u�	sA�F`�m�@k��$^s�ߊ2�0�*�ؐ�ĉ��t�f��-x)�Z,�l,t2?��PB����V�Hͧn�����1 ��JMb�Hì�!�	�%� �v��� D�;�-ni���<Qd&r6��X|����.L��|>������9�
_��(�J�ARg��M��M'�w�D^�y��拓]h�[����:�U���r"�su��I����!k�a��6�M�Ĵ�ӉMy=$�AkNo�z6�{f�2�
���ht]?��oW0%ܲ�������X�Vg�B�ln{��q~vxs��7|�3iD��4��E�7�u�,o*6�ę:��>��჎�ٝ�lD�:m�����������L73��W����ckD�ݳC���X ba.
���F#�	���5�6���K�] ��`�r��`/���Â̚o�
!.Le����#�-1u�Ma,��C(8I�t#:�"k?y�g�e!�ӫ& >C{&����ce	7�wZP��и20�+��8O���7ͼF��(�p���+�r�T뵝xՓ~��_?aE�᧨���G�b���� ��\�ѩɳ0�D(��zQKsYGѽ�uo��W�<v���nӦ��t��I��;��t�u	΋�L%A�����_��ھqY�o5Z=ȶq�`�^v,aS��
?m���ԥ��Ϋ����'�pT�`Q����q��NA��r�!=q~���:Uv}�񥶩n�s��\�0��'�g8�V��p�r�n:K<r�� �������3}���D��c_���@����%�u+O�y�w��5��!�y&W���Ar/���<ׅ�f�(�����cTq��㛙�¥3��U�����N���v�t`����0vK���:�"��>����{�W�-��6�;��*�L��izb�>���َy��j�"�9���\ =o�9�xУp��ښGX�Y��i��� #v�$m럇b�,G�?o�����{GYp��_:�1�/?�p9f�������i&^����OR0���v�j	U��4z�3��8�w�#�w�-�腿F!+2(��n���-�1�dV�	������S|>��nN�����=����9����S��T�Q���n|ym�o
���Xf���ܴ�|�9�#��&���~�9�o>�茠�7��k����0�1�;��'H_s_kC�+�����eP����H>Z���)[�#�nj+VysT/禾d�K��6z;�+���l<bD	��V����v��|Oϸ���u�j� J(ic������(N����a���y5S���*6L���~����� �j��M��mxa|_��帜,!E��ǩ��&ůvH.��⻫$�$��z^����J�ܢ5�5RZ�YE2M�`���.��L��z�ؽm��M7����j��
j#�N��7�)��1(w�j�}g�5�<��
��
