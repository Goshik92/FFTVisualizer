��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjfm~���*�G�	3�`�{��G�W��;�
ֳC�?h��_���=�o��n�(�
b}?'Ǯjք�_Z�ϵu0f���Y�q[�m1�pp����&%�a��|:ꃸ���)�5�N��4k�, ���o�p��Z�c>���H��]At�$YX}�+��lj��^�E/����,I0���Xl>�_��_XLMUDIi#�����[���ZT�ˀ�K4�r��I:/��t]���"��p)��P.#�hp��/;=�@Fj����0�h!S�.���~�	��?mH�Ǭ��Mv�N�I2�y<�ck���*u��_+x��V..�����������`"�<f�{��ג���|��e�n���~����{��1��eWb�gsy���Fn���K|N�v:��Qt�ʉ�� ���c�0Yu%�m�Q�������/a�{����-G1��]��=Z*A�j �~���oRQ�-��eS��w(O��m�:�w'��/���-@Pb4t�& ��h�Z��9��������зs�J��\�����T5e����
�f�vݝ�e�c�9�yz�r~%џ.�Mzx���@��IJ?ļ�^+|�0𥓤���PԴ1���.�*�E�1JO��ʡڄ#�x\	`m�U�%��W+���[��GEaO�J?��+���֚���9Z��dQ��.Ei���4��^�p�E��Eq���d�k��[HE���.}/E����"d髣GE4�9#��s�*M�UU�	��G�^�ǚ*$s@���
������枢�eF�����wG/��]��ԩ����S�}ȹ��7���ŹF�L��6��C?���)L�g�U�[*��s[��!�j��X(?�#�9�����)!Ub��G�s��ZX!AV\�*e��d��=��M��E)|d��&��c�2,}d,*R��4��m��4�з13�BEͨ8�N���$t�΋O(w��}�^M�B��8P��?�w|�x���VƦ2ڰ��?:���p�(q�!�_t����B��$�f|�6H�DsX�����Ū�K�!�Ψ�_T�I	5Eqf��"��P-ʛҔ��H�A�dڞ��������^v�@B�^��s������]{���uʤ{��'b'�={��/��C�qy�ۼTM%Tp�|s�C�k�8:���!6�y�RËqH�V����v���Hd9���-�!�4��z��b8����obv�wѦ4A<ddQ�=Pi��N_�D���Z��RpTu}����Ϛ�2�E����e�e^i��;g��N�D*Q�z�B5B[����K�2�(�"�GY&+F�UA�����z���'�dQ_.�!9]�Y_����4';�����/D��������@S6�:� ����Zp޽2��5�D�KCU7�@ϩ�R�{DIg��q%z�6���x�&�~w�j�&!��o-ˈ�PM��tmKp9W(��B����$N2 ���F�B//�~	��ZVL$��R~(�,a�KU�^�gR�@�$S�)R^����r�,Bf��^j��
Pɜ9��G�E�G+w-t�9H�2+D'ƅ�V��-c�*�ݒt��ק��/�r�Ƙٷx�ۀ���W��p�=el/|
��J����RY�Ǘj� o�cH�Zê�HG��XѴ�4$;�姣���y[���`� ��=�-���1�B k\T �xL�����4���ʕ�*`f��Hz%H�Y*2�&�5���Y�+�@L5�Q�Fi�g��)��hQg#Pk�~1q�\*�Q�m�u�*T^���sF_k2`�����$� +����{~�末ОbǄ!}U{��	����.�[��\x��#_LP�YZ�Z��6�����11}��=�E];hc.�l-��(�aq�ئ%�L �\}ϗ�<�O\J��C;(��T)c8Q�˺^t����x�Խ7}�p���Cg�Xث��mn����8V�D�u{��^`�]:��݀�����9�[y����{?hDN�;7����FQ[ޮ�����ޕ��h���p|�2!�~+�	����e��u�ȆYF	��� r���)v��:���;t1�;��m C���SSY����Q�%���6��':r�6���<n��43��e{{ք{r�̴�3oU����ŲQ,����Z�e�h�Z"��6G�m ��1��LSDQ��ˑ��M���o��X��?���&ɫF�q�`�'��C�W��-�jKܡ�o켯�_)�}Z�T�Y�ծ�����e�����I�[�oGW*, �D?�4E��*Ǟ��'����'���E����ޣ�eA 1�#�F�[��qTڿ��	i��I
Uf7��m	��I� J�ئ�f)\������aMgV�����ym���k3��"l���j����0�����4���m%S�a}N-\KY<9�Jg[H�ϫ\��Ʃa�:6p  �,�0%_c@!�^B�V��/�U��X�_���C�_�S�t��}!�ȟ�
<��Lt��O���	�2���X�+��$ӵ�<M�
�+�)e��#�Md-��#�)xM��.~y-����c+Q3��!W$�Iw�P�����x���N�a��
�m/UP�y����ȷAQ0����	]����`�~B+�qIY�4#
s�8���%�A�L�t��J��kћDٳT+
&�Y�ܓ�l+Mn0i���?�;�}ǌ���)g��p�귊���+9��zt6��2f/�B.83���������7/
�b@����"����3���hU����o�����m7z����~�D���T{r�
��nk���O`5%=Ӛ�r3Xs�_Τ���i��p����]Ť,��h��C���_�i���?b�|~�.얾�\����fx�T���H
�a�̱Mr�A���D��h-_}f���V�G ��e&�<�/H'H��J��~3��a������$Qy2F��h�6�h�_[54D������~�S]���LBil�D\֒��U \<�`�z��q�x��(��\�<S��m?��7=��	�{���O���g�6V:�w��@a���A��#��1�*1�AĄ���%rٻ�m�f������;X&ڙ�$Q�*ϋ�֞(��U��I���}i�w�(5�Q��2$��h�*:>�n}��/�e��i~R�����S�u�,O7'2�+D�&_���D��ۭ�Vi���ps��r��IB�x':ϓ���HUKeu�G���E&�4�Ȯ� 𬧞��Dn�U��Y>8�
�BY'���B��6?a�n���{1��*�����4O�P��[�"#
�I��J��7^��\�	-��"��08�kP�J*����{�� i�<l�}$"�%����V�_%׽��$^s)��5����ZR��s�WR�A��f��S~��XU&�&�	��HqH�3����6ݕQd�~N}��3�\	#�A#�d$Bn!@��j�a���=�ne�����Yu#���0snv�+��]�6\�skah���.��0�x�FU��nӨe�������XJW�OX�]�n�ݱob7w~�qKN���it����Y��we%̴�<�Ԭ�Djk�}����<���\����Z�i�Z�E��<$V��x����ű¢�k��	e/�ѨVC,�*��a#Ei�;>B��y WE��<+�P|t�hܬ�Q�i��s�j,RJ����0{<K_Vn�F�h� '�����]�j�>�Ȥ^n��g��[�P�Y�p�����d�e�yf�ޓ���́e������!3.O�%��q�:}/M�#@��ĝ˃Or�j��7�^�JL��J��BȘ�L����`85������N��8~��H
�P�[�����R�����ąi,����؅�,&��4�
q��)uA����H�H��N��9yN�;���Nj�t]AI������Ď�C��؛u��qr��'O>/���>�N�<�%�32��
��(�H\6���1�u�6��:(��h�@�B��E��8��qj.ޡE]�oz�ʶ��ބ�����q�?A�d�n���ؐ"*�Q���$ìC�9�U��ɩOˌ���V�8&⇸٣��G:y-x���L��B�U`,���rMk��]K�@�q�\�{�tZI�VD��(@{��:p�ף�����0�XOhh`0*�_�,K�����Q�ݶ�S�����d�(,��a��BeD�ā|�w��s�����0b���mĸZ<�j�@�~Rchx]����L���>��h��ɹ��S��b�:�8����c����P \�lv򮑦yL�[i���W�9�~��w���&_���b�Q�}�t%�D����7�=*P~�1��U���3�����x��2���#Э/�=��X!�H�H��%�9Kx.��<�s��@#2���#�\:>*&$]��*͔�	D�z���M29>�$تp�)L�ة���	������7v�Ɂn
�Y�&�4��#�m�����1L1x���4~�n�@�T'�Y
��rC�^���jqz�:��-���}�I�u�gz�a��}h���e��� ې��!Rh�6�HL뿕�S�a�$��Cߧ%fO� x�eV�'�4إ��Y��ú��C;���+ݪ*^�� �;[0q{`�a�	����1���k9�(���tT�\��
��:����yYjR˅�'�ry��ճ���3p�gnmBz����4t��/4��&~��K���hS��-�t�(�
���b�4���V�в�{�^e�<n���U���n<��j|���B���h�^��D���@;=d��*�0��RMs�
a�W;8�� ��y��$z7s��BU�~2�y��:�:�_Î��Ԁ㿐2�HR�W�9q����9Wk�,�#���+��p$�Y� �)�ө���ֵM���Y�`�Yqm�)9���*٦zE']^���O6���)�hEB�-�s�T���q���*����K��4�Q�b�	`]�ҟ�U,�jC.���w�a ɰ9�	^	�{��AQa�5�`c�2x�
����e�\b�{,����I0�f���l�@ w�(���1A�uX�iEBR��6�O>��6C5��s͎��}��6 +��A!>{iCR����]�ɕ:���!)�z:u��%��uև,��J��fd��=Qk��,;(��G9�@O�D����'&V�dJ����A�.��hD͵Qn�+�|��/������ќ�PYSZ)M��֑��ϝ����(y�]��9��Ȯ:�Z��o�l�?�������1��d��Tɓ_��sV[К���,&�z�C��X�j�;Y*��C@K�·ew��G�D�?��4�#��t�;���<���+��0����0-}�g|/�&9X�9@�p.q3}	�Z��A�g���/��*�K�h7�������,S����ꇆ�Gv�_�qc�QJ�x�(���|�c�F(����s�e��J��YCS��K��<�vHr��z�SK>�-����
�!�s����d��Z��t�H� #���s����Td���m��������3�ۍƜ���҉�#��Ъy��mu� ���/���A��k����D�(7��E�^)l=i�UV��GQ9�1�<����!���9B^k��aV�����ă �FS���!����.�����ꉂT���|_�a���U?���KOv�ROA�.�U̬��[�@�%��0:m����S,�m��Yœq}�T.�V_����5�TUz*A	ÕJ����|��'zD�V=�i��A7es����:A�C	䌁�0�9�����5�����B^̐�.��O�~S�O���!jv �XKn�i[�bwŸk7�K<ۂ#�=�x��>��-��%4K��5�l�p�b�]��3sf��-g>��e�/�{�B�.�a&q0�瓹'笚��0�z�9���%��W?���{9G/�r���x��sk��bU��_���&��֮�J�y�8N��®/���ѱWi=jCy��Z߂�3�hR�~ڸ��������,�?2�d��̫�.S@yD�_���1l�"	=�G+y^@3ܸ���s1��t�q@�Rϥr��J���ëP�C��%�.����/���+�D��&0�Q����16�Wˢ��	Uֱ��
X��X�^ ��F�[Ƌ: �e�H٢���D?<�^[�EYi�����{Sc�P���U~�c�!ќ9�(�֓cF�L&��C���3R����f �}�kǡ6��95V��p�g)~��oǛ��l����V�!�[�}{����H�b��'_�I��۞��rH�w|7��ԗj���Es�@m��N�2�Tبbv&q�<S�R����W��߷Ql�k8�N���l��9�'�<?�w@���(bN�v��x�"XH{9Tϟ94Zgߊ�`́Wn�O$4�k�J{�i�L<&K=��f�M�h��z'��è7R�?D�nߤ��;b�F�h�6�����.Nw�P���$*� 
��G�MQ��Y���I0B����&zTո1�'	�baf��C��іxt6�=����X�j����~*���(��(�;X�?��&��n����q�F�?^V��gQ��:�L���1rXy���ḙ�ԦR���ך\]��4�Z��f���?	�0��>��ֆ'z�n�O�����\�����w��I��Y�������q�~qo<�9�<�M�D����'2-�ab����ko�XW3a$�!��
lyև�N��i�s�E�L\R��9	��B�YnN�����,����r���+��aN���0CVй8N2h��=�Y�B�ɪ]�oH�E �yn�\TW�x��`��L�3~�v^p6dx�n�����G������@c	q�A��/K��͊�v���W��IE�&��<��u:$���n�:/��۵��PA��un�O��pw\��P|I ���_$V�_D�����9�l�}�����s��b�Ѓ���Q��S`g�=<��6~�C�4�� |��]%���n�9�^]�fO�I��Y��pV5~^��.����OO3��n�ᦡ�!<�&��U�ǟ��qBB�F��Co�i
�����Ԩo������츬��X��7�[@�~E�N��E�J/�`��إ�������"�� c���y$�gZ�Kmi?ʑ�h$��6KX`�y��rPs�����o`6�%V�s��	,�p-W�$8�������!�w��͈����(w�"=�W}���(A���PL;(E (�0T�B�S^�9��
ME�e"�X����'��)�!�U�`�
�"�CO��x3,��0��'��7&�v��^�7���p@���	�__���G���^I�U��W�Tw���x&�<����N�*v�c�[@ۂ/#}:7����4��x�j���r��N��F�7	��4�Q������H�6)�& Rz�͞���~
�^k�wԀ�F�{rˤ���C��s�1��A=���~��������D�w)��!�}ɀ�5t�K�(�CCw��VK�t&;V��Y�Mb%���\i$��3Dؑ���}��y/�e��7�7e`@.���u7w��_�:��3�ȿ)�b���i�e��oh�"O%I�20k��=)#b�h��K3�&× �be��^<u�)E��Sz�Tӟ�>��ՙ�	�����5�!�Ap���t���p�~Mj<�L\B�Aہ��T@�-��A���]|�h�-�n�G���&֐]Y����,����gV�"�:��o���ݶ�mxN������%Y��sy߳�1�H�:��9�6؀:k�@	�Nb���[��1�/ZN9��'	uT�OQ�d�e	�5�Q���+��'C���]&#��Hd�D-����I�N��+��M-Bϸ5\�p�"R�až=�@�V&U�Jf
���\��E�8Ϫ(�r���Nt4G���aO�n� ۞�܈�я�]��6�i��g��m��,�8������&
a?�%s�&���5�`Nǃ�hƴ!�'S�`5��>S�w9�f�ϨB��h}s��"�ӳ4�6����C<���t����oEt�B3�F���_z�.a�
(�^���1ؾ~��"�S���,Vl-�"����eC]Uu-`�9���R�ٝ}�0jF�»'w��F����Q3�h R��{�0=��X���fNr��A"xG�'~KD���Cԡ���ҏ��b���ǧ4��N0���W�6%z�% �w ���}�X��	]�i�R�|l]el5{k��Z���	��p�ӥQp����e���Y������g,�4Z9K�y�	]*Kr�f�4J$șӘK^b���	�;�"f
T'�����!�.��p�1.��� �5���<�Oa�#�G+����������8��#��BvƂ�3G��Y�mX&k���p������N�*]?#-Ě^)nMw�%��/<&3*ɒ`g�\���$�@�n���vM%7/���k�[�Q���w@{Ε��2J�,�x�~z���`�S�M[�6؛�6?u���m�׾�e�W�kD��P��H��羊k��s 8���?�a]E�KI��ďF��,�Ѵ�P�7��@��$�ń��B�S9u�<)k���/|���o�+��0q�xO������@/�L��z�q�QyNT�p����v;���s�k�1��C� �)D��|ٴR��$��!r'G�S�7r�	�+r!$��+�B�<yJ5�м�����HN׮��/N�yvEm���l�[��Rp�a�ҥ���1g�S���ϋ��Z�--Myy�O�RVi/s��kE=W�Ud~���@sź~��T@���60V���Qgh`a��)'������a��P68��ķp�!ʃy�H�{q#��׷�X��jT;xRгm�;`Jr�Ec�]�E�,@!�X�Sϊe�C��,e�E�F�i[���ŜX��5Ha����
�VV}�݊� W��A͆��Z�
�Am�v�:Y���(�|���~夹(XD�	m��z���������aڢ��ox�MZp`eVe��U<��z�A�N�=]�$;}�..�%!di1hX�� n�}�e8���C�1��;��`TVj�gC�	)܄i5���9vx�(['�V~-ظ\���=2�x�v*ќ�B��b�ٷ0���qQc���.U��	M�xI�`��YV8��=��R0�bJ�9�
�+Γ���>x����t�(i��%nb���	�p�tz��f˚pf.���`��g����"�x�|�m����	;\�I>�$� ���Q�N�=RQ1j�F�gI�~��V���d�A#��%5��H	�Y��1	M�*��f6�u��%�x� ���;c�A6��e#���/[���e���L��u+Y����g	�aOR�D��H���ؼxM�e�H��#��Y_�=VC��I��6ga?�/{"l6�m"m��\��\�y�N}���C윘����!,UH�J��n8sI]��;�����Gj�,_��2z^a#y�h8��WZ/�S	,ůݮ,-o��|��U�"������	P-���m,V��m%ő�s��(��I�wO8D��9�؜���==8 ��7��]�b��O�k� W}ߞ���t3"�*��N$����U:f%��.��Hx �X���J�ɝ�!�+%���P��(��ɴ�Hj��cC�l��5:=��@x�8o� ��X���c&�*��� �;���H���ƶ"0�)C$�tɌf�.Z�"k��L��LF�!B��:�I��18ҶÝB_a;��A�s~���g���d�U���P�}���7!�W�� L�gX�@�-���ގ2�?�
�ܨ/�k�z���ݺ0f�����.��]g�	�D��R�l�\[�9�������wMR�_~��q�'**��uH�<~���^�����;�lf��E��ܰ�$��X7e9+跭���4��~=���Bxx��db� 0jA/��Zd�40�[7`^�Y4w�2C��n��������_TP꫅
@0<�(�[Hg� W���9�����P��[�k�~o�j[2����S76���=5ݿ�a8BI�����Q읱͝��O`�g��ӅAp����:Y���Ԧ�~��шM�PM\�!m.9���&�$��+Xl��j�K�m�wl��?ڃ7cL*�<	1b�����w�>P� �Qe�Fݗ���M3ت���[�����W'U�N�$�=UE�׫5�ې�q[:3��+T�Ц�օ}�Y�)�sy�*��P�F�ed�ǃ��:�+�fc1Ds�-�q\�8�W�ڵ奼���������(6*PG\�>�d����r̐:�7�t7��a������0�Q���Zr���z �U,^�";vp�e4{� P{rT�L�+aF�Z`���aJL�K8��&�;z�����r=�{m.�,���(��E��D�9��h���.�H\��M��K�T��6�td��e�����N�[�ۦ�z�	�"Q�K*-�+����A���ʒdj���?�h1�Yb���	�Ɨ�_�M�ʨ�7J7����&���k��Sߔ���v
D���~�����Zt�z���0�O~�tO�	�9�հ@#�:ǆ�S\g%�4�[Ƹw\-ZIwޔj#�U�vH��"��bq��{���9�<|�\�b���1�����H��������qh�v�z?��}��u� �V���ts���$�S�g�HV}d�L!5�=��6��߮n^M��ֳe��i�ht��CO�b�]�u%߅$��{M����/˝B���Z�CvX�?|����I�&q��9İ�W��	�Y��rATxҁ�?e(�Y����+s�������Q�s��ϠcW��!�߭A*��rބ��n'i�w~���[��;�i��}S��l�M'$��v(�Gl�����6Lj'�i[}ߚ�䞿lJ���f�\�;�#����"�&�"�ٿ�-mW��\� ���?J b-���,ط��N�M=	;���?2#�ygU��ș��W��_Rr�~ν���r�� +��b��4���b���+rQ��� �ؾ�b`
.Ǩɥ\��}�l��%�ZB�Uz-J�x��6��c�ND������$�^uWf�rA��,����<�ZdN��wĚ� �jP�*;��j���_��^̉�c�J��Y�d��B/�U��j��� ��E��uω�Q�-U�[)��Z��&1��T���ʔ��!�_�}T�7|K%��#��U��iܛT��_�KFt��Є!�â1_��vk�-#dO݈�����S�%dMϚ\����*:�Z���'W�x9�c�����hZ��](�.�39T~�����`�����o�t{���62W�W�����*f꡶Cy�#��t�9a���E�p<�DC����s*#��d�j@����G��N�.�-(T�u�pE��������J.yP8St�UF��"��-9 �G	��l�)+6,M���6��$?�;�ڐf.�8x��mi��(�����8l�����47���\�~��5k�˩ϵ�ڇ�D�� �~z��h�����D��xm ��S7���b��Z�PX��g�VuL���Y0Y���T`���{
ᤚ����u0��ur�{7��8�K��#��Y�qJ�p�(]^aS�I8�x]V��؟������� @8*��%����S3�����}^�97]3���_3hY+z�'�c,���ڲ���6�N�������/��l�z�Z �}��f�B�S��:�!RRЩӴ�D�1����{��~I�L�9:�9C�痑//����D���*|c ֤D�(�H�����|��q��y#z�&�A�1�K��WF����#ᥭ!ZYv��=����D�=�h�?Cm"ʹ���Ac��L�+TkUî�,�4���^�2��&ɓ2��Lc��`8���!���-��9ɉo�=h�E��¬�K�î�'	���-(sWoײ_@_7[Z�eǼ�+ez}������K���HT��԰8�1�q�ʖ��P� F��B��ڜ�b���`e�S�k��p�߱���s��qKU>z; ��N��Mݿ��t��̣�|�D���Ң:/8�
_!�w�!ٮX�(;�-NzHmsɯKV;�{s��V��8�+��z+ ��'R�p	 'Kfd�xͮ�e��K �{����ݼQ�h/aV��﹑��1�ƺ���xZ(�\vj>�Pm��ZELޜ�d�Qp����<:�V���e
:q��5��v��2��+�Y4��g1����՜�d��D1VF�<��E
���[o�C�e���������Ϻ����=�w��Lc�L-WEy��tC�)�k�d�K��[��9�V���㳁�M�o�0�ix����P�1e���s����
u�9�������ɠ�}��Z�sj����,����!6t�l��M/�����b��D��� �j�������$�(:�m�+7�_r=�I$���M��H�߄�!+7/'���<���H�Sꉈ�v���-�{m�k=Va�;��#���>�[�v��ҵ�u����� �8����!��2AE�j��������#��yx�	orw�����;$h��{����t/ڄ����+$̪ 
P�L6Zߐ�~Z���
�
�<}~��&��0�5����w@}��z~�W��a�d��J=�(Q���m�"�#uZU�r���1{�{`�ө���Ӽ}z����y2qW��R��<;�v�i��i����Q[�4��ړ���v_�:Bd>oxUʞ~��f���U)ڳ%K,��倫�Cϻ�JL�C!�/��O��,�	ݪ0mR��0veD;yk��P��G|TSwN$q��$���a��q2¨����C��;�$�!M!LI��C���Uf��͔��Dm�e��?qF�:�����B�"�Y����G{k�ҋ>�S֟}��XỊՏ��⊏I�Q�b��Š����Q��a����D��i����,>���֟e�0M'!p-��I�$J	��1bVJ�>��:X<L�X��ʹ�D����C�K*�'SjΡ�u�U��HQG.���?��Y�YȚ�o�Hym�9U�;yL9�o��I�Gi��b%��5/z:a��G�/v8���)mC:����--�Bpb�H9�%Ӕ����Y^cщX���%#�1ؕ�p��4GH���`̚�.���Ӑӵ�'j˺��,�rIfL�[	��G��iOR�{�fA뜴������wM��k"�47�$^�1qA��NA�^��O�W��>}�@�D�\����q7����C/ƨ�8w�d1�~��Uq��R������m�
�����a;9��U��llIC|�����_t�Qk�',��兒��E��9���N�K��:�&}o)�����;K����HCh�aYb��ݍA�d��aiŐ���O}�]�o=�"9Q�ko3��;�dr�̙�'b[�η�j�p���^�JVJɬ8W�@�8�KɈ7%|� /�.r���WR�$���%t
<����"m-q`����w�@9�~�2dLu�mw�:�Ѡ�!�X�2p|?pA����E�QH�Z������V�L�ɯ��Sm|�h�,��ـس�I�G4~���n�m��6}�+}�nTQL�5��fN��]���_Ј뒫&�����J_�w�'MK:%v��1�v.�}��Y�|�������CyĀ|D
�3�����BW��FN�+��H:z_Cz?���� ����ص.�O�~��q�N]z,M�#by�'t�wO��fW0�Pd��@�lw@�0g}�^��ڢUܿ���%V�Dk�΁�Èiz������Hï����V��R��`1+0�����1a+��@+з�ޡgkSZ�R�^�}��}��B(�T�%�l�K㹾9u ��;��d4���t�M7.u~��C�K�W~؎��^#�n�G�ɀ� /���4/�6xG��Swl/��(�G8UV���K#�2H�r��9�Q��`������A�^N1�7O"����or�s����e{$�������vU��<�_o�UI/�����xR�ٌĹ���Pp���<��i��V��[4�5`D$�%����R��n����:Vk_�)d�`���C�4�j��]�/)�bԢ�����<� I��@
].
�������ޅJ�2~V� 6����>��^�I�	�L��W�	mʁ�{�YhX~x�%����*.�L,�=n��R�k�ߠ^�<���^���@Due�����k��zN-�]�~{��m����)�l7p\��k���g��&=�d�!����^eĹ.����$C�PmlT�}�����2�x[�C>]_
���w�J�2�'S���W����ƈ��>.�x�Z�����VFT��k �� ��Ї��ju���q֤������@�D���4B�{���:g����=0���7_T�թ�~�&'M����0��GL���1h|�����P�f��Ւ �n�x�Z�E��9�]<��p� -EJAuq�Kc0V���(R��s���v���W��+b`Z������`�x,�����\�0��b���~�}I�ء��ub�\�T�wX4��|��Ov���F�8COɒXEV����4T5�_���&A�c+-�,][�����G�n�V��،�k)_�Uưyf�i�r�s>{\K{��q�ԡ����e�)�m�\��M�4S/���m^�wߏ;�+�p�2�.*f$�rjN]9��L����Tv^��H)��u���BZ�Q�m�*�g��*�v؇�{�'y��� �����h��eGc�P�!�WDH�qܘU�,~]�:�T�Up���fgf,����J�-;��9^���|,"�/3먙E������L�`�$�:����������?��i�G���ʟҥ+����|�m��QЇް�C��-i�����G̫&8g���R�z9�\�p�7��Z��E�~���i3�B�����\�D54�A��x�� ����4..�=����a�8Oh����(B< �e֩�vzpW.p��$���U�!"p�������%㵳Y�;>e���x�kh�hO���j�.��!P��H`Jбϫ����e��G�UY#䝑����vW7\�b��
H̳��F���A�Ts�Y��+Bzo,w��xEl	�?�v?8��Rg��f�o����<�%(�g�Z�@E@*:`��)�&�*�u�5���XS�C���&K|����1�l�E�S_�#�`�&t�ﶉ��/�5���T}"�ќ�ф�R���4Tdr��\Y	"�E�z^�9K�c�ZN$CV���Ρ�.ٴ[���/H����|wi�0� d���zj m���J��+����R�� &�:�{]�ҡH�$f�K�1ZAx��.�����Y/2��Y`�xo����#cB��el���F&���l��Ԁ`g�s�s�N��W�7��\c5�J;�Y@�´��=��Qt�6��EBi�%o�Q���l��f�l��;.�a~>����#Û������g�����퍜/K5;����K����m���X��Tb����-~X��ˁ]��v/h����8l�-/ ����`8w��Ϩ��0/ibʮ\[�`���k\����mN���K�D�R��`^z�\]���}w1*����. 6��3<��d����D3�r�{�G��j�OG�QNۙ��������pf��yY��4�\�U��m�Qmb�v��T��>���7U����Fhcj� �Vf!F]��߀{4s�/�' ��?�.�W�k�8����Drǃh��qy_����E���0K�XU�����S��R�LZ��ާ�u~	X�a�`|���N������=IR4����������~���Ƽ4xJvf�M�ٺ����uN�!
`��?��K8\�h�2v�	��|��ZG�܆�[���U~�Ǥ/�@�<�sI�%֠ ���͵Aq�f7~:؋�a=v2o"8�U�X8j��3sY���9���c���%�A�ţ�rDS/\qj��$d�Q�3}�����k���J���Ⱦ�|�~��E6�G�OE�)|,�nEO&/������ٞ�q��Q��X�[a�;��r�F%���>���*�[�X�3]�)�&�}fʹ��p�I��z�8� ���S�WqI"�-��2�%��[�81����7�+�tYP�oc�Y��tK�Vh�2N�������^�a֬q�D��º{R�d��r	�א�X�� �5�l^2Jf���a��¥;�א�f��p�0�R��j���&��rK&�
��`Zm��F1GN�$��6Z�e�v�zʛn��E pI6����"�>�2�����C3)B��n ';v�=�t�8sj�c�_��t�৵-�ןf�βK��#�&�/���3��&`��'$`��(��Rx{-�Ԑ�Q���$�@��?���u}L\�iS�+$�І����m�(�}i�&q�DI38��U�J7C1l�Vk�9�3�
��C�V1�6��}�?vF�J5���w�XC�s��-=�X��@d �"��Gc�L���%E򇔥b��y�����,��2#?(v��79�|h����� r�*��%?UI9���&U�)�:�`9&oϊ�P�����:[��āY���e�)��-Ol����As��0��2��c���e���Ux���R�?���A��3�e*��`���fW�.B�t�##�i���{�y��=Y��~*I)�?��䝕n��������?��x�"~{}�i�+��7s�B��9fHh��ZSI���?�zF��B�G�T07Q��F2yv��l�m&T6���ylÑ]�K<����co���с�m����Ѩ#��TZ��5�8�����~�/�\ǥɯ�[p�<�AM���Z�rK�f���Fd{�i�ES~���߹7���y0���;%���)#g�To�&���s�����S#0��M�DW��<�0��!���|K��z��|1F��|���VHT1�iT�B�u�{A7a���������^�mY�2��:�
Vj�-O_YsU��fw7I?�VX�!�^�?9�� 7�����&ދ�ja_A3��Ø�����|ʆҰ����s2�0t{V�Y֒�ʝ$]����qWD�ʣl�?�X�䳃��?ڻ@���T�F� �#�%�E�D.�s����E�|a^)A(eW��v� \d_���_��]ہ�}�J�A&�7(r�eF�0�`(��E�-�}�e�âJ��Y����P���}ٍ�s��ݿ�^�ZG�j�bf��h���V�YH�w��˽��x�y?"В�V�A�����Uq�	dr+鞽�?�ݍyK�}�Y��c�,�����z,�]�x�:�L�8�ب��W�D���T=$	Vx����h���.�'��W����{(����{9�����f|�|��x'?�1K�����5�_x[��8Q���y6���v��7w�>�v�`����r�����9�s�F��,-�}�"�%�'��O��ݗF�e��>�]��������:nD: �&��ۿ�� �s����_�m4_?��=P�8�Yg�ꓓ>ع����)��&���������H�r��la���Cᑰ59����(�Ɉ���Oj+?M�RO�-���;eP��J>r
�K�l��k�L�"&�!e:ϸƤY-�~��d����^�T�gyL5[�/�B������6���x[ ��Fs�ݰB��׏�@"��WNd�G��O���6`iؽ�}��xߡL>�a���'pop�A�#ŨQ����|J�����2�������2�V<��D�IY$-�P�(�^&0��}yfb�����7�a~"����[��+���"���s�KZ���ۓ�k=��Hة��;��ⰳ!%d��H�6{�P-�	�bWnY��/c+-������C��s� �?�vBPY��ޭ�/��ƴ!���\��C�i�N�{������.� 5�̢��{`v�T���^W�1���$�Q�4T
Y�bXQ���eFf/\���
���(��;��3y0�d:kȘ3��R	7K@��r��\��j���������Zk����d��J�0���"�p5Ø��rǺiH�ުK����sR�;�Һ�ťn�l�R�%��	E)�m!���]��t���?��'�GL]��ϧ��뀌K�n���i髪
cP���B/��Z"�3��P<)e���]i)Htm���^ڭ�Y�nH �����'d����O�G�"��w�����0��Q�h�U�AU�I�x�T�	��@�����񲒤����Ϫ�6g�j�۴�����w��)����p��xTf����d�4�}��0���tJ2�x�t�F����M���3�O;��'?�^BJ�h�I�j6N�-�W�Q=��!��q�H�4����H�%��m����op"�y�xu�y@f-�Fx4�m���,GK����?���]�R�,H���?��սV�����������$�9��Y�i�2d`[&rB�����{7A�=�*��9}���(���(M>(}�.^�;*ꦖ!T�)�D��-0Ht����X�s8���g&�r��W��Y
�`{u؞��|�؛�)�?��뻈��|-/�ht������@��[���f6�+��%�A���~��ߤ�N�	:�b����Wl۬�Xَ�fG8iPB���0�p���%�0���M��J�?�L20p���	F����3��Y��.�7v�F�ec-hW��#�Ǳ��fu��E�ݙ�K�>�`��)�t��w�E$��Bϒ�}�,";���8J\ζm�a[�ϤAַ#EP�G�}%���j�� ��}�Qv赨���-��d�×��#at}�+�9�%�#��.��*�
���Bao�3�E�#�B����)�袝]F4�uLK�c���gBKT�`*3�	��Gz���8+��ݶV`�R�6�Ll`݂~���%P��@�T�;~ì�7�5r����W���p�����g&�M �8I �H��r"�7���:�^��ʵ�yF\R#��}͋\u=���0�h?�O��O@{���ep�5�L��i4q�K;u[�}|��3_��/ ��y���ǝ�����x�`7R��B�O�cr+�2�u�@n�/(<�?��<	���T<�QϞ��O��v��
I�}GR�M�����q��(�!�E������E5����E������ᵵav���_��ބN��´%̿UʈW�Ɩ��*��1k�"l���r��������L�Dm�8	F���0'0�����ZQb�!d��?�vEl��U�� r6���74�F)v��a�@��48=WˀW���2Vwr���Q)���L��*Sp��M�Sw�dO7�N�2ؗYBq'��Z�5O�cU���_�i��#9�)�kbZ��Yr�Ac���w3N�4#h�����B�^3:�%5H�u�<ػ�b�v�eCB��4���W�o,H�L���Γr�x��w��U���KWdUD,x�/ \����|��h������3Kw�
x��l��3��TyTr�|Ȋ�����qt6��
g�q�K����~�Ki��)o���XY��\��T��+2c3��~�C�Umχ!s̕�������wf�k�c�,J����/9Q�'�Z��PR�Puz�EF��J�u 9��t@�:j4&����vV�L�/[�����c��|�1vQ."Յ�&�➶s�����h����:X=h��^�Rx��`�4��{��4�˯�AW��"�Q�ls�r� ��$}f�O�w'�
���!딐�l?���*x�S!e1~*�m_��j�jo��0���Z5}�F����KQǰ������[(���e'�'�L��TA���H߅�fw7�XQ�k��x�S�Ic�^�a_���Ҩ�8��B ��H/��y0ܘ9>ez^j1�^���~w���bNX���M�+�(��E�8�����ZðReO#	��s���i�8%�%�[a�v��>�t0���Q���C �x�U�䛆��%jki�堑�g��,�s:��HKO�,Z�|{ ��E+��N͘^�����n0��b�px��]�z��<67O��q�g`G�$<�G|��C#�#���ec:�&��E>��{�]�8����%�ܣVp׿���)�/,�ExZ���BӃl�&��������Y;��6����͜����\����2vd�̃CL��>�����.��s�g3����7���6 �A���SH4:��%���i`1��e���bN�VF��K��?�@zG�34?Cp�%�'��i�����	 �k�(]?�^��`�Z��=����y�b28${^�Bx��fo�8���5j�ٽ�%���Y2��Jh"Z��y	O���&o�dP�p�P��4��L5�11Bj�b�>�Tiğ��|F��Ǒc���&�Ҝ���]�C�%׶�*�X��ş�����Uܓ��å��P~�C�)��+���<>��&���08�r¯����r^w;��XO����p�w�J8��\!�L�rLظ����+F�*�z��is���Zr���r�?dj*p���xΖ+��C2��F#���۴��Xن+���:[TtE�M�LD�@P�]��E���6�O��J}Z����As.Ze�CVul��*���� ������0K;w�0�W��W�;c��+�z��I�Zs��*ڝ_I��^?sl�N�T\%�lhUXOj��#�?���N&8Í�t����Gy���ߝ>O8��2���^,�.C�g�X�I#�B����/֐~4�R�Tw��Z^��Pv�/m}��SF)���k�.��'���pDI�k;�:8���,�c�[��#��o�Qè^ee�H��1ԋ<�[��!%<�.�=����8Ҕ�ƍ���0���X�s§�)p<�v�O\��[[:��o�+�WS�O��'��`n
��p�,�5�,�֢t
��=����h�a$�M���8��0|�4=�yȲ�S؅���	JO�Fђ�=�1�d�^����,֧��[c�<Jw53?�&�.Q���h�۪ �����@���,�Iu���O|�θ���*������t���EI��}�y�7�5# eOW�s� F�EGi��l]�2�P�)�B�YD@t/y�Kd[��	�K��p��U�a�45_'���NKk������>/ޘS�����JÝ�@o A���u?��r���XX��I��!�
��h�R�����}TX�Gf�S�: "�SEUߙ�~~Ƌe�_����g�A� �8�B�-1ޗf��S.�u�N��-\>\>�4������F���`$���t�3����x?@�GUM��(��=�!�6[��=]%��j%�*L�Ά��yP��[��~'a�K��/���V�u��kJx=�dQ�5^�=�0Jd�c��*�T��:�����6���@a�J�L�L��of��F��*P����8�!�ğ��A4R(>�~G��h'���Ry�=Pb�D�����1�,>څ���1&���x ��E(Å}8[�'sR�SbX\�d$e�Hvp�}���T>ҵo#N���%~	ܧ����2{а��]ȩ�ֈ��b�I"*s����T�^n��&y_�{�-ĩ�JsΟ���L�.w��нF�=�\+6E�[�D~��S�Uq� �m�º[�ًq�vyJ�	�	b� ]**L.!O_.��؝�x���X�k`W����0/��H��\-���B����i�o��.��g���(���S�(FP,���>Q����98���� f�n��o!�����0�O*F��~�bɛ�� ��Bi��)�A�1�$��Sa��iI0����?��Jh��y��m�#�$��o����܃Ăf�j�[K�ρ�b��ʰ߿��91�݊�<�h���}�~wU���A%T��Ye%����0���β��b8�sN��W��p��'T �9���ԝ��`��9��ц̋WdQ�@w!W�3�{��$���r���^���&��'k��8\q� ~ֿ��s����3�?�΍�DՉ�d��kD(�7ģ�@2��@��v��W�1	��2be�߮/��4E�A.f�肀�v���x�j�~;����}l��+O"l�#�3"�K��>�z_����'�s'�B�,2����T�m���~�+�����
��2���V��6��U=:���I�S�B�:'�1q#yC� �e]��H�^�#w�cIT���
�_�p��`=�Jb>���)CKv<���ߔ*<f�8J#�9�K��hO�M/������	[8��V���7K*Y]6��cL��q�[��Q�xսa�r�~A�=�'i�vCsW�
p���W�Ǜ!/�cI�S3�N�֓2����E3���ygQ��}��zPq�!�J� �wd��9۬:Y��������|L����j���ĝ��o�tM��˩�J�gf�
66�Ո��ѩc�>��7֊�t��]ܭq����}���R��j���[��u� �x~#aE�"�i+_1|q��{�"	'�5�.���A�o���$��cͯ�A*�Mq��k]�r�� <�cta6+�u�;P�UZ}7ꪒgw����b;��.��op�h�uL]y0K�K���zK�WŠ���;Pf�an���Xs�Õ���4�ڮ. �-)��q�s���3�$�y��n?eõC/-�Xh�����_���p�e��w���'����T�["{�lb�9a欟��Z�[����(> d���\��n�Z)����{��"r�9�^~��z��h����a�Ѥo���[�?���v�7P@��oى��zbrU�ԑ D���c��YS��^�*h�|�Lm�]�ưCY3i��~�?W& �Q����63k<�*@�Գ��z��@i<�0�5��i�,{l��3�������=:?���U h�M̺��,_����ۆ�S\��ݯ;ߴோ��J�q��m�}�a�jgs��B�אY�s�MBy�>e���mM��%�n��o޻(Yo?�r�Ԝ��*�o��>����&���?!��>ZT���|�L"&�q��-s��Y��3r� ��v�!�������I@y�66+R���N���x���	�ۊ�k��Z�Y�|�`~*.9��(��6�չc����[v�
���K.�y|�x&k7���m
�$�����nh�����^�νN�ҽ\�ׂ�-��9ρ���!F���e�H����P��0D�(�[ۘ�a"4����7X��ߎhK| KQ5M�s���Ydl�ׄ�,�>�8L�.Փ�����	t�JHa�}�.#xْ?Yև9l� �2������x�*j=d�P�
?��@�����ob�)Ɠ
;�Q�Q5��7VnT�A�Z^���G;/ૢ��ޅ?'1����ʻ�0/�]�����+fѿ ���<V�po��eY�b�
�=�培$y�nΏ�C3�[#�C��ےo���0�J  ���^+�;P2���V]y�t�ח
��4<�cR��u��Fy��	�L,��a<�+���g4�,���	��F~89ف�hNE�#Y��@��(�M�8��+V�:�C�\x��7���G�t�N�C�73��:7����1�<<>��d�o�x�y�1 '!� /O�[O�D���OpG��s���Z{�5eR��<'����j�R��u���4��.J�Ҕ����OHc��G[�-�Z��Z|�|�D�2%��� �p�ǋ|��{�%���f+rAup�q$=��"�C���QY��!c�SV	��Msa�TT~JH�������T+e3N�E&�.��by�ubk�n�C�0Y?�R�]7��n�be�x�5j�:�d��r���"��y<eQ�6�E� `۔�2�m���ZŐ
�Nt�`q󖏉�K�W|.��}m~�4���A���P{Q20Fa7�U��s5����%W�e�\�rxJ�=���Cm���逺����э��9ɉ'c=׿��r:r�B8�*�l��?J^w{s�L��<�ĥ-_�NA�=���ȐYs$cPs.�����7�C�Y��j��U��\���Y�:��\��`׆�v;���>��y����<%�#��8�b�Yηp�a�D�Dw�}�e�`�n����TV��W�Z@%T�M���	�(��� +�� h���j�W,��mD�JjFp���G�ZS��������
�8��N�)E쵵��C�BkuTӾ�x�꣞��&������y����[ov/���5F����rm�wn���7b��?_�Nw8��qi�,81��d[��;��+�lG� o4۠S��'�6ph�˿��*6��`�u�������Ϩ���0�v��6�V�Ϲ�ڠ�?Tl��p�VV��.Os\Q� �)�=x�O��z�o��\�U2Ύv�K��yh�B��(�;g�l��Rܹ����=]Wb����V���Z�e�/�^���2s����X�ݠ��_O�Ax��v�����}��e�I2����]d��H�N�wHtυ!�F���Aq�B��Ӗ�\��{]w�N=��+�ɐ(�:c����u���}}�З�'�#���Bٚru����ȧ�S��Q`�
��SOZ�Ԭ7�^ը��F4�C����v�-��]V�	�k�%��^%� 02|�!S�" ݾ��K%���v��}4E��gC����Ӌ���)��ٵ �%Fc���G;�O䔙�T9M���g�}s4Q�0IB�Yܗ��W\tK�"K��R2�g�PC�~�~�$��yQ����O��3���r�t���c|����h�~�P�]�̳̒D���X�m^���۪0�� �5�oQկP'�G���#nk|wOT`E�k��dI���f+,On�]�J��=�W�
���°� �0צ�Ǔ�E�PV�����(r���e�C����b��rL5��H}F8h�D�Z&��mW���{<��r��m
��0�U�a}#S�=���$�O�A�S���Dd�Dގ�VӷZ=���JCo�8�r^��=]sɼ�����b]z�s�������81d��8R5 /�v�+��a�09�\�z���lSf7��О�(����jGld�'��L�5Է	�{)�T��hU�~��$L��S�}��H��k�y?�чJ�F�"LṬ��x�[8�3��v���,2���E���)^���O_ڐ�cV��11{ִ���M��=s��#6v�v��s��qxru�N�d\�<P{OQ���Ϟ�B��_��E��)�@qYJ��J��nP,�w��7�'��1�(�<3�aFF��R�r�����K1]لFJ��<�������<M���$h�s����q�.������V'�Z�z��M+O�1:u�^��2pJ�ă��?�9+�b�>���-���PW�E?�$���<��|�*���ÃrI����PwqmE�-;���������/!��Xg����~;O�c� �}�׉]�r#��5|iseZ�����i'Y��HVq��R�O4KY�L�!b���6W�|kb~�	� +��bЇ��߽�L$К��P���*���-
�.{Kg� �t��QS.�_ԃ��C8��m��$'7�iܸS.DMdR����ō��bF�%Gg�ī`�є�\�����{׍}b��Y�"�E��N��ְ}5�Y6�}Ҧ�d@D��[��R4���x�X�[�0
�vx�5�Y�C�T�l��,�$�&�������E$p��mqY���羪~�~����4��A�pn�i�2�&�h6,}�Q� �D������aT�@v�ކ���L~ =I���^D�N�~{,Jy�}wć�?�����ࠚ�i�oA1�4LM�[|KغB؄Z]���;1F�Fh*��*����	�('���̦�<-�U����V@��(���ra��K�.|�p씓��,n�ШVA���B!��8zg$3�g��8
A�(�Ί���:͖��L��a���+M�o����b�	G��z��!������S�5�Mx'̅�H)Eڙ/���٫���`�O�pLt�/�ɉ�Q\]M܃l!0H�cEQ�ܡ����칾��ݝ��s�ډ(�f�g�d+c�<,S�|�Y�5�,��)A��E�L�Yc���}}(��ҽs��'������<稥
��KW�K���*�w�e���TQ޳�F��I�\�4�Z�$1�:f��Վ��)��������˚7��;'�e���Tq4�fO�����	�΄�%X[� �@m�>�Cm[�ɾ��@��T��Lݏm[8��M���/!1$U:3ʲ��cV�]p��=�m����V��S�֮�_�S�;e��I�x� M������[�T���&�0+nwv����A�c��\ة�t�i�'z[ʷ=:�����,GIJ�`U��-�֚1�-���7%G~}����B��'�MD�wZ8����/�.�4�^K�}�
�E���َ�b ��T�Ho�8$OT{�q �ȹ/�#=��@�	:T#ŀ'���KjF�7�M������s(5L�S�E��-�G�ї�Y2�����o�%�����Z*�@D��2{XS���BnH�rU9�)��C��/PC�?�|�]�q�*jt?'��v�vk$EC	�NٜԐK"O�� ���@^��a�_�q�,e�	yEo��/��3�$)q��o�s��q�Y�"ė>����f���h�S�9�t�/����܆� �O���׻�W��t� "� `���Ti�����<L�HF �-�����߼�RByu->(�|�|�y�M3A�Ҽf�PtZ��rB����w/B���� �aXL��A~�-i��j�k�"F��n�a�ۻ����S?}0/��	�-&�������pw>���,�����`}A.؋�Ydoً|�cH��0o�/"p�T��G[��,EL�{��a�3�(�k�����������~r

��U�����	͝�M0ʾ��N���uS��vK�b^R�r�Q�3Pj�;zc��SZ?�p#4fm�`����&A�PC�<�=�ӫ�1������;G9k�/���l�H~f�-� ���5܋HoWn��a���r֍��p;M��X9��*�n��P�5��^��Dg��Z�9�~���N�@�)���Ti����B1���CIR�Ut�S����Ī�)�8�� �tRC������x^7'�o
{<�]�.��z�����=`>�N�H��B�^�:��\q �_c�p�0��1I� �,��
p�D5x$DHh[\w�r'����#�R_	`�	{s��ؘ3���_�\W)�x