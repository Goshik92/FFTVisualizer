��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn<����d���+!����-������F+)shxj�IHЊ��x�`�q+��"-�X��(�������*��4��l�`����1zyG<�Ao�&�I�ڋ3"s�Y���؉a�'3�s���Qm��B�" ��֖���R;l�L�W��Ȏ�EAG��2=@�ڷ��@�i[��oɚDj_\�fo��x@�5*��[���/&Co�g��ؔ���-�J`��Q3j�h����lIVt�& bѾ#s������g`��ͼ෹�C!���<5j�"c
��m�=�VZRepO_�ui��2g���3Ŭ��0m�ɵ����y���:���M��sV�U�!��������B�T^!G��9���/yVSۄ�u~%���O��H*D�=B'(>.4�TU~�z>4&���*f�)M��=�'%��+���w>b���M�ɋ�����"���'��o�^�tʸr6n��R�Jx�`�D��W�(�qVn���yC�k�4ƖaΏ��z��������k�~�^����fѻ��+ �2�҃i�P��&��n�������B��6A%��=���2a�kX�R�u���5�T�"zx��bM���4�����t�M7T1`�Df��L09�F}��Jm���@��.Ty��iz��m�
��-]R_I�B��� ��֯L���"�����܍cЫ�Obr�|�E��, �%�����X��6��'`v����7f�JsvzKI;9���v���WaAy��/ZB[���Pϝ���k�Cå�R�sd�P)(B��Q�����6s����oǍM��i]�zj�1�'�X|�l��Ѡ���z۷xBtϚ�o��_��=de�T���)�Ф�%�(<��R��0��ã���\��m�z��I8V�����B�{��>���I��	C��y�o�+�(�� @�~ǹ���N,�q�Ӗ��'�z���S'tt+ܻ���K��p���>ɲ�E�h�D��SB��6x�R��W2B<b��Bz~�1�1���k�̋|t�a����qIĝ��ջƠ��U�1|	<,�ܽ�Շ�C�7�����Q��b<�b�5��&X)ûӬ�얪���*���`�������\GAF������?�XӤ�,S�}��F��dOT�x��0t�F*��\�@��[ew	��%�[�õbq�����4� �h�6$�!4}��9�ܖ���!)�	�Ƣ�n���O��k�Q/h����V���Aئ(���}1�_�tX!���B�xMg�:_.'%�Ÿ+H� Z6D4c��Z�/ų"}6k)�x~�T�KI�e�����'{�N�
~�	_CG̙��C�r��@����~�+/6ܬ�j�i�E�!I�F3�7�(��� �%4��D2�=�� ��_��]^r���w�������rF7o'z����͝?�L����Ot�`9�
�!.n�cD7�����D��{xMT�"�C�N����	cM��>��A��M�P�����,���.��e���>�X�A���(����H��Deql�7�a����"u�᪎�a�H��Z��j��.�R+��}����ժl~w�=3͒����(�F(ҫ�6����eC�����W��I�ª%����Yү��c���k΂�|��ч���� 
���M��G����|���:����wv�Ѯ}e�3�5�b�Y~������
J&��;���L?%��e*²p��1{��&v�"Q�o�P����x���v�M��A���W��K���� �{F���c�,u�{?�G��?�kB�5j#����7QEU^w�a{10I��W_e�j�hQ1�ճ/ɏ�q>(�D|����q~�_ۜ����������9�ئ�x�2���a$�l���!�"Λ��O�glo�7ŉ��R�`��s�����p�ݓ�A����˛�fi^{��J�Z96IE\1�ê�e���� 8M�,����u]�b|�?�/tZV$c6�a��\�a6�����" u���!΂���v�7�VѢ�`}D e�+)���(��_�o��*��^�&�+��;�򰫪��2G�+��8\C�-��p�A��VYR�����w�d�0��~�76�P�#-�w�	���%������
�@ȭ��uݵ7��� v0����li�lU�XPp
Y��$p�dC87xH��M���M�����_�������ż�A��&v9�Q��^5��Gf�|*�Fs� �ә�����5��u�Wj�r��w�N��i<3���[&��ڮCm�Ү�0�-?��=���7���
+Yj���I���S�O"�}����9�x/�5W?��A�}G�������U�W�3İ�P:���1������3螻��O��(q"�ϳ� `���8Ǐ�c;Փ�P��3��gֲ��q��H3ٖ����2i.����Y�VhZ�ާSqC�_�����h ��w�^|xWs
�r;�!�`�թ��.3n�Q-��o�`�\o���p�V�pL	�{�<C�Q�N����s7����~��K,:x�w��5�![� �;�c�1�"2�Q���wK������R��TǓ`�\�w�ۥ�7A�>��
�3+&*8;����7gЗ�7�v$�"ă��}|�#zA��ު�p�)��{�k�� r�v��+�|���M^��p"I�Q��7�O�W-m�iՀM���,��K����|-���{`���{�ju��bu"*�Pc���Qz�;D���[�w�9�\֋�#<�u��p�F�N%ߎ���ܞ��9�pI3#�~k�- �$@�	��"��k	}�JJ��ޖ�B���y��"u(3�U̹�Lu�,d�Yٱl��*hV6��ߑ(`V�K>�_�ڢ��'�����&�����o8�*{�\��,p�!G枊���}u��u���tβ0}���wL�KW�35����)J�ئ�et3܀����u`�l>([��DS��xM�"RI
8z#�ॳ���kN��:<��^��B���ȫ%����(2�Q
����`�:�jY�������[�]3	b���^��֌�E���U�)q
��L�pL(�"�����GV��D�P�mA��Ȅ�{b��_b�\�iZkb̴;�Y��D����@����Q$�7/.h�߬�tY����G��Qk��eW���/��,~O���Am�����bm��l�[҄�Yp���ܭT��P����?D��B��!v8(Rtu2o�g�˜��;���0>�J.����2w��JD۴��i��0�$i��2~}Z1˿� ��kz���mQf���#���_��z�z�R�H��BG{[`��x�ePg��sr���"��ϑ鱲�Ҟ\�lw�j1*����/1h��p��c)���X)�A��W�ЌZj��(�����L v.���͊Fg�
[�2}�'Deԙ4�xX����P`���'gƫ�%l�����<".�p<�Sl'���,%Y�l���w|)><�,��L�X���j�#��P���Ԕ�;��j�����~�A��3��j_(ޕ�u��#-��ǲȵ�Y�k	��N�9������8�s~|�#�F+��>6�,y%ɺ���ɭU�£B���w�;j��P;�J6	�I&�������<'�u9/��v�jI�y�P���]*����Ղ���V`�OE�=F�	-(t�ٛY6�g7��b���m�Zr��Z6��N��I�f��u��H�8�m�7ǅ�:��4�|���/~�Ф�*v�D��j��?3����L��5��)N@K�n����j���P�H�_��Q�X��'��NL��z��Ğ����u�d��R7��<��;eY�uGs#�/N�Z�5b�)iR�L��:�ڃ~�N��o���%0P�lbY�_�b-e��x*B��5��A��O�Ö���|��o�p%��U���MgE�L����i>8�bx�RIᄦV���h��9؀���r贯\R���e ��-I��Ѵ�_ce4�:�o�	a����b����,y��\fk�5_�L�N�Q��q�����R ���͆��;{��5����хS�v,p\�� �T���A�Aq�_V����G�u�e��D�d�����H0(�~���m7�]WDG
v��F3�� Amj����
��7Ii	r�\g�����[�e�8r�-�m`�,��JBoj'�J�[��0e�"�ŚhCZ]�rN�H��-w��m`f,'��Ty9+��y�R�Y��Łj<(��ͯ�puT̛~ڃ�:Kɍ:���MzsrD
�ʨڟ#����ձa�fb���xI�B�4���������&�-S��S8�/�C�U8�l�Q��wB4A�/g�Ĥ���G���d��ޭ���6HU�>�1��/% �ALMJ�K�T;FC����`�%d��u���I'�7cz�YB"���p��g�0]�nà�z���>XF�
��6I� �P�ܞ%�
��p��	4K����A�����䘽�x��P�O��XJ��V��~���{�)P�d����V�S���� ����ًw�q������qk(��y�h�ϫP�ic�J܊�Y�=�C�W@�>u��2S ���Sx( ��a���Z�z;�����,p9��
3B�O�w%���{��?��=u`��e�D)������y�r�V� t>V�Q�!K;	)v�aO��G0� _�q<�S/�3|"�tŬoA9�3Ie�zR�{�v�<�8��_�� �G[��uo^�-��C��k���J��Iέ�ǌ��ÍUFi�=d�x�����ܡS��๑��.Y�4��pt�c-���a�n5��7+�''�Zt��зA_���I;�&RoH����MBx2���%�'-F����k=����X|0����I��o��ۮ��� ��_Œb���_5�q�t��V�-���K�?�ؐ/5x�(;p��E�A����y��W���Jl\^���J�I��Ll�U��g���1�x�vV)\��i�2]_z eN�WzM��+�S�
�J�W};����8��o��cA�_%8P0Nc	��8pг;ٲ���:_����ծ���c�J��	2S�=d�{[�Of�y�d����,6�]�B�cc��)��Sp)��"7u&�+�?��p�����T넗��!q�?]G1n�Bm�x�A�!t�ɮ��Q���^�hҲ�M�n��&�B���a�ʠ�v����\�b��C��O'�\�7���)��P��)Xs{�5���3�!�d�U�m�/LD��?+�
ߙ`Z�rxoe	T
����M͛���RΦ�ͩ8�]������-X� �I��I�J�b@��M'���:�m�g�,B��H�u^&� ;C,�����&�T��u��6VvP��%m�,��	���ʭ
J�jX�#[����u��yi��v.�|{��>���MFۨ�Rv3[Ia�9�\}`S]���߱k�u�d��[��^A%���>��O�`	�2"���b��Y,�\c��7��׹�<]9�bo�~*�j�����D�2�o�A,j�9��h�7P��B���Z"����➾�{����@Y��@�
�i�4t���I�[��6Kt�-���Jm�x��8�Vz⼰�&>84�B�j5\2��Dߚ�f
6U��"���ۧII|y���"�������q�9��+i�2���05K��HF����pz��Nϵ	*J�!��j�$d��߰{�	d�`D(<e�Q$]_;/��ɳwn��+���Eh�� (��X��<4���F~g�Rb�A�Ϝ�E,e�9/~ut��ы ���+Ĩ�����d{SSlKo(�i��_��7���Iq(a
��r�|����W�gtv��(ܒ��xb��c������⩃�Z1�'���%*k�Y���$(w�Ǵ��ٍq��&Bo����Ä�&*k�qq�e$��}��`�V\��<�����?:L�FG���/�ؔ�2Gj%�Q@��}�J�_��H=M��$���0��8�aK�#Y��Z� �b��L%��)ӥ�͸CaB�@b%?��x���(���f�x�� ���$� >ܸ:~@��d2ǦM)��̧TP���{͗�Bqΰ�Ҫ�O7��@��c��@D�!��� ��c�����;?���໹��[�<��շ8��r�#�R�YM�1P��Nr�Zy���&"�e�^GQW��7�t�����gvȅ �Ltr��7�lȀ�
4��	�G�`�EI��:{w��e,i�h>8��vwu���dY�J־����3D!]�l�qh_�����D4��}�u_p3(���ۈ��U��+���(�P�7�ⳋ���lJ"�C��8?��3����?��G��>�2m�i Ef�L��b�$h\@�����k3u#�#�m�r���? 9�aԑ��M�S������h_n�����TUQ�Ȅ�����ʈ��}�`8�a���.|Q]('�/���H��͒�%/���Nk��g�9j�!>+���h�T���/�˃-͹�����
�z�YǨE�TA���������@kMU�[�Ԫ}YBs u(�=5i�7ޅ#����64N��t����0���M%a�t�M�vG������د��pT�O�?�➾����_6��]�n�S�;a��I{bp�H���N_����"bPC}���|�Ȁmv2��]�6�L*�5���ۗ�T^I?��P�1��b+���@�7_a�pC��I�"�8�"�$*�"�$t�W��U`�Եr�4���m��4�V���ZCvHĸ�}�U�&�/���'3k07��}�f�:��?�1��ܓ>b��]?i��@�G����:����!;u�V@�~Wx��h�Xu7Y_aP���1��V��hn,�l)?�#�&��
w���vtix��x�1k�T�v0
���=+kԯ)����ģ8�E2���O�;���Tl���|�9'�WGB7�79L� ��M����J�D����e�� sA����?bNsx:�Ák� ĊW��!�8bh��p�s��-v9�_;2}Z�*�(�@�܆�M�x��?e�,A���e�gقwe�^���puw0�L� I��$��U�2~�('$�R_c��h_IT�W*0��x����>�w��C\�`�Ws50��ܣ��.�1跕�]R�lx�l	�!�������Y0a��O���b�}{P*�|N��@�UwaU����Q%Ɵػ��mOxiJ^�4�3ҴO��	�k����Y���,�	�M	���̯:�#���@�7�We�	�l�'m�I�X����J��z&���yQ��";Ed����Rz�831Cb`^���{�uS�OwWz�T����ԏ%4uB�G��)O-��>�8Vhf{�|�v�����(�6�o	��0"��|���;4F� ��KF�q��yXus~�zX��V�ē��O���7�?Ў�N�\�{�b#�ʨ���D��zk�3v�W�Y�@�ύ�?�u<`\u<�r��_�	´�"�P?��M���>�����#[�ؙ1�P_��f��C��a�jܢ�K�#�p��^�D���J�ܡh�pI]md��r\�u�<;I��-�?^阮j�#���Vc��B"|X�^�;���m������!(��L\�$*���I^t#-��Ҷ��D�B	1�k�l���<�C�'����z�M��;��d	�bO�V��h�Ԩ�"#�y*{�,i��D#{���F�>�ȿF�����F`|�� �Y���0�� �C��Pp�8NۜɄwU��Q:���� ����)�hc���I�)`\?E�Y�k���>�	��c�Y�ZHc »ضR������qf=�yՔ&�(�lYK�#N`O����kdJIq��}�@�+\�Qm���a�k���[$d�&����	�2]����3���z�,�AGĿk!�)�-�v�kB\��PE9}��T��4��*Y��w
|�ɢ���dP��#��[��2�|�;�0��;�^�9�?���== ��T+P��?��]3VU4c1�/uk,-)����( �ط ��,s�=�A屷 ��ќ�!9l�W
��F����)z������\Q�\�Ȇ�ܗ0�.)�b;Sws�*]�ڞ��8ߧ$�?.����Jgmm"a̛��(�C�u/́���:�Q/	�.w5щ!�͛i�-D(cn��Ӫ4Q���-4{���p{��D%\�yб=>�ke���v�$ܗ�2�D -SbݳMR��tӳ(~��'��*Y�}]�K�>�Fi`�,�^�{����k�T~��.���5�Ih��\*��374����ЪސY�[��d��%$$������c�j�:�%+§�71��7����x� ���ya�(=�K*�������^M�1��D���U���0�_s"L���H2�3PdW,��?���+�A��a㻷81��_rY��g�A�t2�V�A�b��!�G~&�C��JJe�,��������XYc�<�6�b+wT��T��9i+��j���5_ߘ�.}$��� |h����x2���f��t 2��_���4G
��,KP3��ʝ���g���~�ic�W����j!