��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��We����x�j��ӛ@�G�C{ �`�*��k�Y�u�oM_�#�,���ֵ(v���?���!��ˌlo��V��٧���7Slh�݀32�)X�"�#Ţ�� ��͢ڵ�z�Ґo���	d� ?�ШS`60�3���6�_�F�L׻���1���c��\/����_���w�6���,��?w�f5�N��Uk^Jt���'�[h�E�\��b�q�޼�>�����_L�P�6�B��#��܇E�K�v�%�����1��K�5 T�u�g!����ޕE, ��I���u�ՊAL��*BtĔ��{�3������nd��1
������� �<�%���rڝ �l�h��>^d}IO~/�/,��f���k/�';��iz5�
�=�~�茠X���/�����h�H��o�Km���{~U�r�
���U0����ި��Nh[Y����:��C۩�9�GNu�V���:]A���"w��㦻Ю�����0*��5qV�d��EH�LnK���}j�����3%�>�ɏ�<^-.����̖�zz����ib�s�ء���g��bƾ;8�r��I�M��!��~�Q�~G���Gr�����1�F�R�-�VP��C`y/�}&Ce�>+4ar,[2揉�o�d��r+�M2�jV|�l�1���얰W`³'z~a.i�fA��}��} M,Ϟ���8��\NW�Y�H]������(ڴAЉ:�P赌v�����4&�9f��H��(7w���úSf�A��s��1�46w��3�U�]�D��e�V���g�<r����}D Gь�C��膩O������+�sT�"x��:6 }���7�H�W%y�Ƹ�Y`���D@Oc�4�zq���k�r�e����K`9����;���}��R��,�l�8]yA��MV����$Cˠ6��ӭV�=�#ͳ�.2"c9G�a�tP���{���-��o
R��Ŭ�����Z���앫�����0f� ?�B^$��;b�?��ٲ�C\��zm����gH�_z��"*�("E�d��g_v*�;���dQZ��Y1�����;�֣]�dW��]z?��UsMso�9�>����൞ר�~��x6�KGęg�_~��$_�gu�l�|��$��{�I���H~��"X�����F�na�C���9��9���E��ԭS���D�*�8r~va
y7~[uP���2�W-�-�kc���ј���08U�2��搃!�%"d"K��Hp$���i�Ώ/�WÉ��z��� �y`����/�(C�v�D}��Ցs���lh�C�e�������V/��rG��zCl�y�;��t�K���f8X��&v��	
�m6��#�=�:���=�ב���7�k��h�e���"W�����t����U̦��zR��p�Zy�;W��
M��.�a����������V��Z7&\��Z�Eq�92zN���4-����$���6u�b�}T��\|2n��0@o���J�\����4أO�
���k�&U6� E[�f���z��'6��"����)��܍:�e]o�WZIѤ��.�;P5�|�V	66ƺ�d�3�)yv�`��fr92�k�X�f�v��!T�ɀ��:��&+�����u��Y�;rr��c�1u�C�/�7�T��?���1�"�YhO
�����i�Eo�����y�s�)����$#����;	[�ߕ"u�
XF�Ň���lx�9z���ֶq� �Hh�X�܈s�4tf��� E�eG�^B+��֊)�CB��	*�*�:����H��*�s���)���,��M��c�'�)��19��ᑆ���2i�\�I(�~�fc!g�[�	pE����S���Lcs2��sr��;��@��[CD��r!���:�pVK0AA�&K�J<yF�UWG��/���{o3:��(�6�����2����+��{
��VE�D:mg����\�~1�d�\sO |�@� x�S+H���n �F?�V,v��k�5!�t�A^��8u_2���E�%�� �d[�F]�tl.��s���{�J�Y!��?N��\��{�G	�����H�}DLD���'� ���)���?'��3�P��.�@å��J� �vK"J��r���Zo�[�~��
�;�����Y�{l�~�²�M�s^�&3q�.�!>�烿�%������$	���4��ff�[�R4�[�mC{ٲt+�C/w��`��UlQx��c�M|����-��}ۃk�S#�sJ��K��%��Kd�UO�O60V�z|��z��Ux��sC�e1�F.*A�Ju3���r+-�16K�b������e��W��
o�bߓ�aW����,�e ��+�m>�9�b�^�v�R?�
����.7I6 v��բ(���q��E6�na�[ ���ۗ�x[M���M����3?�Y4���0,�E�e����O�/A�M����_�4�&�|]Y|-�᪮M���r�c�.9%iȥ�_:))����}Z��~��~N�T�E�̚�ӂ������Fh�PZD��pآu��$��%$�h�~"�cc{`:�s66��>��tp�O[|�"�� 6?��,ɏkMq<�5�"�q|^oG�c~���VaC��V$�<����n�dh]�/hy�ŮEr�"e}V#��k�'���������/�9��^��9�-uz$���5a͸pɛ��	�-�ƹ�y��&�V��7R�ú�_�T��6�C��P�/�I�P�.��cW�#3��R�V�CIYlN�>}����L١�7O;��$ȼ�J�D�qV&�=u�tf��as�:Y��'dIS�j|��'����D��.�}�7�T�]FPA�[P�洵OkcP����ۈ>��mI�$�����A�X�jP\WO;fK2�;L�*��56�<�#<��5?h@	R�2꤅s�r'R�8����Dvd��k�h�Ŏ����x�$�e"-;%�)t����
��L���X���R1�iOԯo��6��{A��~XH�%'?�����$�&:zޝ�Yc�b>��aA�ED�d���l��֎���i�a�?-��30Y-Or�MK����aSgm0:��>��2_�İ$���Ak�!��S����'�b.<�AS�Ph`�U�n~�ˣ�T6D��{R-"�f�!Ժv�yl�z��Ѱ_ͧ%q�����bL��J�Pv�;�w&��t�v6��OA72p��Ƥ�[�f'8Fќ�Bi��-:U��ݲ���"���".����nQ4�(�{ɺ�~V�?���h��hF2�G3r�������2l�1� �5Rj�^�H�q?3��"x!��u�ܩ�7�=_L� ?�x(
O�b5�,wTN��U�Ot��2WO���e)����>�\��� }e[vNnxu��Y]U3�z%@~�N�!��v�"����LQ��
P�c�y�A�I��}���ƒ��o���Ăw�ss#��KU��S�����%z�E�\����ʆ�^��u)����	hm��1Ѱ��M��Df��ap���ᨼ�U<T֩��{)��B�3��������ʖK��6J?���8
�V�X��j ��o���F��HOd�0V��^�(e������ h�a�@��rd�f���i X����n�Ѕ�RThnFyۉ�v���i� (<�A�Ǌ��%s=3��)��:�����m?�w�w��%�����m~���-��	�*>�w=ZUGb�r��	�˄�Lc �XP��3Ԝj��B�󢄸C,Z��������c�ӨIW<q�k�u~�\���)���=�,��S�7y(��ɉK���3�NS�)y5ٽ����c^t�1��l�N�䊙��VX��]Ȼ��ѯ�$9L���@ʭ�~&6��W@ �]�Mq���C���cx��b|��V�gƷM�DXW�� �Hlh=4q[���h0�@;�v^K2�/F��z��꣇Ѝ��03�� :�vay,��Bo������V~>e����N�L��?q��U�����ս�h$J�|њh_hz����Ԡ���̑����=q�{F�,���W<9(/�_̶�>SJ�vxj3��h/�-Y=��	�۰��u�֦�&;��9	� �s�-d�u�N�-Ib��c��#��,Ν*!�SD^gR�rE�C �7��V��7?�����Ta:������TSus�;���
&""~���q��OT>����;����u6��㔊�j?(�8J+�U��(�0�a�H�w=��Vs�_u�2'ٰ�v����p�s�Z�6�yN��"�%�I���|�=wQq�Z�HL�Y�_R�:���6�P�sEC��j|
�� S�¨H���P\zQoL��P+5����6���y)�aͱ�z�TK��K��� Zt�$��Sa����<�2���g��Z�%����ghk^����]b�/G����Q����������X-�"�Ź4�M~�Ef�jxƕ�|e�t'5v�uuتJ�;\<:�p�7�yio넹";%�wd"��sơSi$����7(����6o���C���~$6B^D�l%"�B�~�u\���E�d`O$?y�����\�9����~���n	] N�g�ۜp�9��)4�@ne�_a��ҩ��y @����b�)�0�m _f��8�Е�RnbP!�n(��߼8���.ɲ�h�r:
�i���G���ع�g>72�T��m�������A��8#\\�m�� �ޒv��v�1�/�P(��l�� �b���v�)�ӝ�F����lDV�
��T
0R���9�۳�yy�?yQ�V�����IN�ߎ�Dy\��aǃ�6\�8�ѥJ󒧛����y�P���]�훒R(����Y�4;�P;>�T�)�U�B%�I��O:0�C�/^��Cv�N��_b?���km-�Su��|.�:���lI��>�Է�98+*#���@<i9%����a!�ƨI[�8ؙ#�&��7�m���J#k�u���"�سK�a�����@�!�R�@�E�Uz��]��!���H,�SAۖv�6�0��^���L��n�&�վ��9��BY�#��؈�X���i�}�dpJꏼ�X�[����5�r��PN�Q��'���M�����e<�O%���x�U�`O8lTcUN�NU�;�B�k{hQ٪/�����}{G�<?
ｼ�q6���^�_��Pj�+c����]� �OW'��ɬu����y5��@�d�rS�H��u¢҅~�j��*Fn���w���`9�/�M�L��iÅϛ̀�<��v�}`�p��|O���vd-����H�Dy�~���M�����������Mg��S���$d� �	�k������Ba����\,c �	���7���ș9qly�"	%�R4����
(�^!k�:�M� L>g���� ��s����#O<����8�
��DF<8{y��fرAM��B@W�fSx�����dI-G��JXr��~�)�Kl�$�]�w��G�}q�Xb�9A�U�j�7�|r�-�X�C�Z$ ��ۅ>��u��xy�w<�?�cuw#r����mG�9E��Z=��=Cb�s�N�+r���!^�������3�4c0UtLRҍ�==@}������V���*�~7�n���ԍ�l�#{�s�	���Wf�<�"$��*!Jj�df�4�z��`j���<���I��Y�1�i���s���H�����#. �K��x�{��(C-���T�Ǌ��6���L�������t]�*\��&�����M���rU��_W�,��q��Iz%���{�A�����[�O�P�m����ㆶo�/�t��c�JuR���&ŀ
~���wsc�oDg�ӯYW³|ad+���<H	`h��f"Uឪx7-� X�}W��]E���i�n+��ݠǨ�C��y�<f��y�>~��) լ�t@+//���2�`�G$��[:SEmi�gX�uQ��s���PC���z7c�UcaL�� �9��o܎f`Bo�Ԗ+��@���=n�� ���Ӧ�fƍq�� ������G����0�ǀ�����`x�lP���ў�Z����2p����[e����<�`�Y��0�o��?^afpTb?=~�G���4E�J�}6N�(ɢ+�L��$��-R�D�lX ���b�	UJe�x4#2Q�i���|��C���zڢ�ۏ
�-`�>��|3����D��c"��9�D$\����|܄�fi���xcB=�8�U۸��Bi�&jG�]���N��t��O���H��~J棯�2�4C�.j3�>����g�!�
]�&�'l�(�&- J��/x�YQ�Mza�d�Ey�����T?6]��<s����݌Y;z�Ɵ�^
��-�	����)�����֜��dV؍��hM"������y�-�ey��L����$9Ey<�
����z�(�gq�Wtj� �3E�Xj�_1.;4d'�:���)��n2F��O)�	�������DW\,�|j�� ��~���غ�%L����p�V��;$�I��{�DK��� .Q���dv*^tIi��F�MI�T�\�ZyNK�c���Y�ݸ�Kw}��7��7~�)}#�f��7Y�Zᤉ]��T�����H)a���S��^`	iκ�w����2�-��4�W��F�iհO@���TR�S���l�5~jVƑC:P�i[[�J�v$Ά�IɋV~��W��r��R{�7ǶTS`�{�v�HI�K����>)�N$� ��!"�W��Ԇ��ώ=r���X�ą���Z�_�%k�Y���F�u���"c�2wd��}ioЈ��k��0����v=�-M0�m�CK�
��⁽/펔;[#/�W� (��O6p%3G�V�~N"ܟ,,�4�gƱސ�M��PF����`[����,�]��7x�"��93.)��nkf��9����g�i����A�q���f$��(}�}�q\;�v�˶ᯩvQ�2DO̜/�m��f�Ǌ�ءB.�)^�7.����˴�i�O*l_�V�N�=mk�pgN����Z|�<FY&���Nk��4B}���2s0��=�����,��$���@Y�B�r���˂�׸`p���n)��C�ȓ[,,�4ᐦ,���zE�~���QUI���d��}��A�	 ]�eb��%���@1G-�=Y�ɀ��̬�v�J��E+K?F�#TY����uR־�_:J����{X2��1W�TP���� }v��P�˳�n	[[�-JN�)�r5nXv!�)�Q��ͽ�*�[�QE
v�Y/gW�ԧz�����h�u�sg�]��ظ��a�zi �&��w��O�H�����yG�Yu-�o������Ġk,*x�~�6���"��[�j�X`��˪_D�� B(}v[5�oiT�m}B�؃\}q��'��C��wz1g��=��v��Q#o�oYF������wq� l5��E_����d!����_���!^	���S�����P|̌�����r�(,�q�\7B�HŬ�X3�CN�Q4�YqG�Z�����L=cM*XPjd_psObD�Kկ�������	�OL�����
���w�i �G?���f�AEK5A���w ����'���}C�b��tX�����3^J�����@/@��42+�$h3ϼ�������8���qkyi,�]姤:���yP���ge�-����쓌zOo?$_�A/��=�~��폯��j�x}�`�s76��B��є�a��}E�+�?�h0e�l��Ha�赑����$x��G�Z��X�`mQ���'[�.��¢���U/v�f�c�>#�&h0>8&�~�h�Z�h�&�4B��`�y�E~��&t�PD��r[M'���o0���	��1�#��
	��Z�<��}G�J�[g7n�9y.�L��`vI��.���p���I��ⱞ�=5W�?��n�EOK��سY��_�gBP3�9�V�̙m?1�[eO��X�a��l�{��vvN�]��"b��|�>�O��v�����Oc����Qrƨ�����ş�rbY��k�����xYwJ�0�� E�"l|���X�M�����Y���`ͤ��+A}<�u������@dwG�l	�!gM�I�bx׸f66�U&( ;NdM�@I���� �E;�1
$AmL��M�^D����+�,�n|��c�������d�3�XV,CAòMu���M6vS'�g�a'Jl���}�$X����Gt���X�*�@T��	@���F�;r��@�/����)��Y[8!xy���ܑ�t�(�e�j�����(��p����8E۹�< 45�⧎�şN-��q�մ
��0.�?W�lT����a���<1���U?�ȴ����ʍ��ՐR��s��=*�l��4e㳐�M����>ğBz�����ƷV�Az{R�1��kd��j`��/֝��+��:-/	��'�6�R�k��?�h�7�Z�*�����)V|ꦪ1���'sZpҙy
��;����묻^w/x�uvD}�{�@8|xO����w83�*���K�l�gzμ�Ը���IiuC8H�09rc��RL���z��p�P��J�	?5��Ƞ�n������ȇ�����lg��W�9��Z��2�tf
�D�nl�]�w�/ZbX�B/�����������&�b��f��f��vb�`�����^��S��hU0cH����W������ss9��k��������Qoɳ%�LL��Y'��j@�d�3�}�8Fk
D��
��S��j3���$`w�b��̉A-�X��� ˲���>���a ���o2���v��C�ֻO�h�SG�t��\��_˱�a���H'�ƻIgU��
VG���C!u�Rm:Ο�A�5�(���ʘa�	@���u��o7�7�����ͧ���G�
��m�>� 
�&�c�:Gr\2�o!��ovk�-��W�Ye0��(�[���3`��'j�e���&�]����rx�������=v<�>4"ܡ'�!�1T�@GB"���Y�v�[�Γ�ڜ�3��.�.�!�]�φ �0J	�J����*�&J��@���]	���r�Uݤ��4S�(�j�C������5�
��:����'���T�&wM�W�C��D�����	�;���׹]I�@�+ �z�)C��;\�U�
v������@��[/���}ݾ}S�<(1���Ֆ���;�
?�S!��h���D��Cxo���N�5j�rJQ�X�,n��b�}4�������R��G-`��WJ7�1��9e�?�r�)'iT�{�P9�8.�Q����qo�+�7���P=���OPz}�f���	�鶨+��K���m �������u+�n(1eN��+��ۊ6>d���Z�O��'E1��CM�Q� ������z�c��uA��w���g����9pj �q�+x,\����Ml�/{���a(8y)��_��K.}�J�D=	75
_3�����5c��9���I���S��CO�h�^�9�����e!�����|	'l�l���"�{�1�r|�̙���8��;f��Y/3,���6]q�nj:�9�y��r��Ho�e +�+��%�OxkA��1L�����B�����"@Wb|���ud�`��>��BJ�ǿ[�?R�6($฼�X��|=6�O��(m@L�z7	�&�1���5���]t]�.�H��ޛ�*F��j�y`i�W
��R|��	\ȃ��5Oa�Y�`2^�����N����-�n�P�Ҩ�Aw3w�D��rݏ<?O�����X+��h|�f�W����N*.���[a�M�?�J���h^�3g���B�Y��bܣqH߯�Ӊ�q�w�����1�uz��W,�\��:G�I�8��Sm(ziH�qc	w�H�� X ���tf��Z��$DG&MR?l5XTmt��3�T��ݺ��@�׎�n�7Jv=��h�c�?�����"F�G�L(��O�V���`7���!y`+#d�gK�T���m�#ҕE��	��og�z$xNyq/L�J�x���TH^�{g��ҡp��@��4-Z�;��[gF��t�E`u�/�8�p��v�ꭾ�r��k@qogy%���ʀ_�p�`V<NT�_�dZ���~<�B�7�c[pF�3�[��M��a���7���D��jq�ٴ#�m������^k�z�i�^6���t2���U������Ս���+l���9�����_�x����\�	'0��n-."r��V-9���3�Y�"3+�ߍƶ��R�cٸ��܈V@KT��P�ƿ(YY:?m�Dv~��EN>���#Jֲ��u�"�zH��p�&��JF����ew�'�~�>'d=�t�,9M�f��0`�9��dDt�ez��M��O%�_�ȇ/�4]�N�9u�����5�*{�b R��R0>�s�/7��h���X���"�@�w�Hl`z��pc�	bL^��n��ଧ���?8e���(�%�o�A ��W�mT��F�?�R����~���t���x�$zDlyw�Ao�o�>�l��`n��H�g�R��
˄��
j���;�'��J鸁�.�&gy-�ϔC�<��0k\=���� \�A�s��Wν5�˥�Ϊ��A�+:���\P2����$�q��;A#���K^�&~��&Z�e����֑3��:���C�p�0D�!�������|�~!� �U�i(�ʄa�o��K�ϼ.u'�Zx������x��y�Go��$i�%�E����ct��S���Q�Ԡ-�lQ��<9�sU\�T�]��� ��9��Ha|,D��{߉E�0�&\ז�pڧ���n��Wr�K7���)VMkZKH��?�Bl�L�8b������=a�J�<묇"��*y#ǰ�g���L��E�e�ܣ�(�󔣶�ަ8>K��l�9�@���}��^�{B��lF�A-)�b��<$��g>��C�Yk��Ge
��4P
�nN�*j�wi@��2�ζ,���䛉i�\5Ӗ_�\�"F���㊶R��έX�u�Ⱥd��4�}��BPo͋�