��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn<����d�l8t��L'0��e����?�O%'ň�5Kə��80��1��Ø��@�>�h��EP�)��<�����h�a�;ԂcfO��c�v����p���u�ӹ�(�L|��<YƟ� �+ږv����a�yw�D:Z�o�RO˨B7�q�I�>8���d(�46�xEa�E�����
qn�9�w����,���f���A �6�߶��!�EݤJZ�|���҂�r��.�}�O�#��U��L���L�%h0��?�#�����r`�5�C�Q���_�<F�x�-��a(�/�NnݵXl �.�M""6�n�6}+H�i����Ep�M���~��=��?h�$�����!�ІH��X���{b��2����ۋ�� $�E1�9��^G\��q�����������SE`s�f�]�ο���G�ɉt��)��u� 4���	�������d���v���=JM�
��*�Tc1Uh��e�5#!�y*W�SX��Z%����^J�Ͳ!�[��;�L��$W1��1p������t==��'zघ"��A��Q���rd��Ƞ}��W���j��Ԁ=�'�	��%'L�i5c��퐉�[�g��"� �n?mZG8\�IV���yꚉ,�.�{qMT�]7~e���L]�{Q�P6� f;� s&+��]��\u�o\�g0E�#Ƙ�pp�K�D� |7W�����ƍ�iv,%�s�h�-T��1L-�o�\g��3J��m	��#���ݦ4*����N�M_͘��s�zX�ؽa��)wNY@��=�)ϴ 'b���W]l���=��H��s�����۰� 9mD���1����wa%m��Zj���ܷ�μM/��.)��z�hf�%_�V����ԗϐ��n��F�"H����)K�N1�����W���e���� ���Rw�����}�]�#{�m�P�l]VEI`�?U���$!���}n� ���jl!�':
�Fu�>n��$�|�l�)R�%���U��BV�l���5儻FETsT�&;����5P�C_�N�*�.d��ʊ����;j9cu��è�Se���*U��$��f�*7�Ͱ�$H�ė����Z���}di�Ri���1u��\���^��x�����B�XY�_�R�0���1n�=mO�'#ìg]];m����c!Z0�=$�J�^d�"�<�����5�j��ɲ5��w��@*����^(�x�x6��:&�k#OΣ�T��,��=*_��v�_P��w���K�Tx��ƾ���"�b�9�w�A�dw�K�r�eM7�
�e����5�5��/�Q-c�E��q�j4I�u�Z��œg�Ћ.m��.����r������5��ګ-�ﳻ�^|b��s��y�mB82� M�8�'�n�6�{5�nv��j��<���=���F�������Tp�W�������-u��+\��P��o�c\"��#��JT��!r�Ft�����ǂ�0px��5���gCu=����N���dS�R�v/.��2(5�Q�Z{�w�-U�y����s��J�'\Ɩ:Y��E9�f,�a���:ME��{�w]��<0m!h#G(�،���r����FC����BcJL�@9B�s��_q�c��{ ~({�K5ߝX0t��+�����0�4�m���׊2O0N�"3<�u���9��k��d1G�{�Q6ŉȺ�A�㫨UT-Ӧ|'�0I���9^G�����x��O`
Hd�E$��_��z1����/"6��6F�4�R�5@�}�����$�L���?�V%����
icf�eU)����d�R���C�1�w�lH��V�0b�D8Z/q�L��O�WǢ/�}�eW�l��r�o='�BOku����4s��Iod�+��oMK�T.��Ҩ9A�B��0Q��
�V���q�=��uZ�
�y� �UG�p���f:�.��ƢL�5�8r]��/�"��]�3�}�)�N��S��]�<S�ʢ]rt�w�~"���Yá�Q����"�0>Y�(�z��
�H�;�?*�bf"��/����Αۖ���<�Ȋ�Te�_��j�v�o�g��9LØ�n�}Wp�V����<���pM�ln+�9Ĵ�4<ɳM8�d`X��F���������s*�5x@�n��ܲ��'��=ݠ}�=�.�_�#�|ݯW~?��qC��E�L=����� V�Z
A$�H��5���Mp��3p3Ҝ�ׂ!y�����x�+b�q��Q�7��f��M����H�Ѻ��,�4�X�|����~��K��r���T��615:b�>�>ae����G@u���X$\�u�֊��K�s��P�<�_��[mX�<�Q�:��xP������yX�Ә$�I턵
VU)ro{�t��,t�)��`�'��}C��`'���;)}"�w\����:>�<H����֕M=�v��bw�C�@,�t��[�Vڇ��&-��wC7��kܑ5u����-�Aʮ�,F��)P�j�շC�Q��!�nVQ�p�8Mkv��Ga��3@,ݖF#���������?���Ȭ��o��&�����̪��R�+�M���	�R$��)�
3���k�
�q?�:`Yi-됉�XA)~�v���X!��}���.`�o���j�Y��X���ci�8�N�ga��>��+���7��E �N��^`�����
�W�0Y�Y�
[�J�q0�QK��Ga蠊R��mW��s�v���V�L�$b�u��i���F3��9��k7s ���K�����d�'>7�u�ʈk�?��B�p]6͹i1Z���$1k��a�%�=��W�|�L:<����	9�Y������>e�����YЮ�2h��@]�~ɮ��JiP&/x�K��v��J�g�_���:8RM��E���Ec�PKjs�A%���K�Ng�סL��(�{a��hV�1��+�up�~�-��&}^z9[�3�s�bzH77Dv
/C")���R��a�;�6r��hM6zM����W�����g�	d�cq�����>(:5<2�CZ�u�Qj"z�7�c����^'�s� ���2)v�HP⥡���T(w�ES��0�Pl�8��w8�ާ����Vٍh�E�}M�C�4Fw�O�2�t����;�l}{<I�&I�.wՐ�������/�xy�g�4Yqz{ߤ�Oa\�]yL��=�����~�QG0�����j��}8�S_��vO���s�@�4ڱ
PK�X CXA+���KZ����6ӌ; ��Y�M�Gm'vd9kH8�ZѺ���}`��	��e��J���mP�Tz�g�LD���ޯ�>��F���U����G�Αe����vy�@�}��P�̢b�9��(������@�?�D�	�K"���s%q��J_7P���.Ag�b.��y��˽�ۙU�
w��O�����y�VG��9��%���7N����k��<`M%�-K/�wZd
�����+в��`w8کVkn�����gC����Yl�|�	ly���)L_ٮ<�hd�d�k�V~f;���_�`���w�W��!�/ǎhM�P�4H���$;������@|���ϡSTg��t�}s� IJDM�]y�g1��g���� 3+��ЀǼ�̆�D�V\%g�ٹd�6�G��	5
��y��tm�Ȍ�
W3��]���o$;KI�Ҙ��;�|�j����x�)h�c7��1�&�Hln��l�}j��@Nȅ����Cp�D��X��MC=����Q�T+�zj\�=�`*��AC,���'^ٟ�!��`�:p��<��9sR�P?���&[���P{��o���t��}�4��]ńV�-�$��Ks5���l-�f��H{ώ�>���j_S�	�6z��7��`���W���"�٬�o/��k�I�n�� ˂o#�(X����C�0
x�)��t���{N"�8N%Ȩ���C��h���$�^�^�D�!�<�!�17���R��U��#��x�}���nu��}�ob��p��h���<���dU!OǑ��ag�|�Q���e^��`��>�`n�f�9�u��e�����_�)��
�)���V�&p�������f4��E��ۇ�?��$N,oU���ϛmڬ�p�M� !ß<W!�H1��>oZ$�%_ބ�X| �-!�ُ2�ngxQ]+-�R�����|8S�+06�4>��o�Ү���hm_�N'#+H��湹��df�m����͖ �e�tU��P��;[5[�^�Z��Z�H�Q�+;S.���=NrC�+O�2�Ԭkǋ����+��f�=�Ձ.h���u��1Q<+M�e���a1�"��ol0F��J�`�E���O�S���p��،l=��Ď�q��fRT�3@���X�����t�6�L�臠~:(Bܠ^��P�z����؂+�}�G6,�H��B�b�K�Zd�藻�%��q�~�_��s�Z9���9 ��3�?�'<V�,<�?#���M`��P��dB�ۓ�F|j��;&�6%f�%p����\)	֒�K�N^; �zH߉�����X�0�b�0m�¥R3)-Kjh���&�ٯ�m���4Q��{�R-���*�D>x�D�@��*��Ō��K�T�ұ,$���h�5�Pc�_�)b��Þc~Ty�!��u�* �
���0N�
�;U���j۱v��t��W쑿���V����r�K��Ҍ�w@��ӽ�%.�`N������y34�g="������pѠj����x��� �����Þ F���py�;"��X#��H��-2R�G�;�&���:�����A��Bosඊ&HULY�u%Z����;(�cN�OF�B�.)�i bC4~"��d�C��W��tw�B!8�W��ajE�������l������#�18��Og ���J��v�0���N5}�{��h��	�딙�N��lc���M�A$�x�%BH�M����<�챩�k;��V${��O�R']�o��5�+J�$k������-��=/�P���5�Aǀ�QAn�x5�w��1�޸��,�`�Q�"TϚ�!E�	��0gV�;�&��f�}���q��)�<��T.��� b��]�kQ{"L-�_PV�RK�B�4�3L�d����S���{��j[n)Z��/H{��̽�����42��p<b�3��"����ѐ��BHQ��Ԟ��9Wm�:�3��2�"�4�ķ����Q����f����:�<6T���8������+b��B���ANJ�}�<=ԫ��դX*�0G���=�YeU���'7U��g%jX;2�
A@z��CA��	|�X�O��ggW<�E(u%(|��=J1�.���W�A����wT v�´=x������z���D��=�����yzU�#���#�F_�2�9}V�WFR�3�v��8��5=��s�y2�y�Pg��xi��?� �^2=ō�ښ��d-9��)Ә���Z���(��m�W!x�vU�bMa$��  ��3X�!0(��Ĵ"�_ɠG�fLW��)��ሔ��?� �ow^�"���N�[���k|����a��of��+��9��X1��둖;�H��o|m9�f�Z�7N�V���Z�T ߮��"ǫ��ߑ6��{��wIy�ݑ�����2\6���s�[z�|7~>N^s�?c;S�'""ٱ0Cݷ����&�䓒����-�E��J�� �Q�����c�o��&��Z=vMx�c P�^[7��:�ի�w�R�ds:/<�_�KL+͜9˳F+7�ޖ�0�å������e�	�yt��G�mp7#F�� �=Yn	׏[#l��WFw�db�S�]���a���?	�y����S�j�Yv�l(�[G}��ޑ�%s��l�~.n�QO�t)g��m�N��Bi�f%��i Q�� ��B>st�H�n��0��J1���y�oa(��	v%_�o��&��}
�����Ahm5(u�ydל@#hsg-�
q��4)h�3��&f�s�8�.���嘬CJ����n�$�*ն)?��#�iI\�L�d*�� ��gp�׻�u�=DR\B���/����F�ǽ�DG���6T��oS*��M�#��8!c��?���D��D?�)�����San�6���_܂�<���5�E��R���ND|� ��k���0]՚#��	��q0�w��zs�|�.TS'��%�i�hX� �9��*��W�|����3^���XD���'�m ���z� Z�bHM�Oi�UR,����)��?�����>�X~+�^�),(�{���G�����M���*呌�u��A!^�w���$�u���"�,��YK	xB��Pe�#2��G��Z5��Cޫ�2Fu� �7ܣ���Ga���D�9�sGP�kuP�۾D�]�	��\��{�E��пr��N�ͨ�I���[m���?HN�����j����к��QcD�r���+0p�ԋ�Nhr�>6��Jυ�nRB	��~R'�Zo�L�/FPQ�S-=��Ѣ�b��2/�B�=2��^���ȓ�ǭA]�]S�I�P��LH�N$���-F����'O�#�8C`(ʒ�>>(�6�ég��I�ґf�������Q�2�.�|ê��*��T8P���a�;S��a�f1H���X�*r+��+_T�('zq���.־��SL�;�kL�!��$�#��fZ_�G(M�F�~GՀ�;D��$QsIz���䋔��������P�;����x�4����8Q�\^�D��>�R-�@* �-����$����k�]�����I}ʄ��04�JZ�z�����i}Ƭbqr�#@�شb�A�y�咄Q��{Tp�����z�{�'�h!�x�����1�	?��4�����uw站����s>��Km��F���-A_�Ѕ�N�P��տ�Q��Mr��g���y� �����!�T�zg��n�e)��o�L��޸WV2�t�@w&����j�-cg����8v�Ӥ����Jg7��[='�vo����B
t̷u��:Ew�-'p���R�� � N$�`���TnY��F�p2��,V5@�� C��?@�,���@�O���1y	��1<1+<	bD���P#Q�L��e{�-�g��q+���DOi6A�ӟA@$y�ډ�,r�����Ö́�5|���1�Kl�&����>M#�r
z�R�d٠���Pu�R�V��	Y1ğ�n&>��l��g�,�����!