��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn-o�s�X7��5�w�RB����F����{6k<A&����nW3jv��������b	'1���$e��0(�ǝ��Յ��c?�A��Y�����)�eD߭���Ƽ�j�p%%]��0���A��W���]%u�O"��#�1+�F�p�r�p\ �&��\KN���H�C/�;�[����`�W~��5�X�;�̊7��+TJ D���Ү��x� )�E��m�ַX���>{EdN(�zBx���j���́�(Sk
��& ��q'xG��0�*�S42��:>v~g_�o���;�|�H)^�єD�}��Թ�8��` �a�y+æ'!�_��3� &wyaC��
�d���Q ��[~�n)�F	T�R�b30�O7R$4(�W{&��?�esr�c{�H�&��U/�hT70<����, O�	�ٜ�zT��\�ғ��=�����r�:Ri�c�EY�W�	lH���r�|���}�Z�c16B�$�tc0<��C�Ӧj�2�׶W�! ��mz�س�� �9��G��P�No3��3`d��2��'Ԡ�I\'�O*�	������Ԫ״i��xĆ�f<�[U���5:�H�r)�H�q�u\����g�V،�]=��8�<�*mΜ.���_)����r��dl�}������
�0�[�@������zd����N�̧�^��ԥ�fr�*{���%c9��s9A��T�i��N����IX�"y�,�Z�z�ޑ�W`;d7qR�~Q�^~2��rG��y.�� '*>�!���p�zu-.��H���Y2�"���
י��S�?a~��'-��x�qk�eQi�W��:�#�Lh�,�V,kX�EHoS�7�Ou]o�����^�S��v_�p*�d�����8��
x6�.�5�����(�/����&}V��W�wl��p�.�
�U�r��q�^�u:��[�L-r�^��t"�t�ew�o����f�ф�l��J�&9�{ w��B�q�a������`,�9L+�3E��!5�o�C'�V6��Z���'�]Ԓ����ޭ3l��W�B
YH��'xA��i�M�m)�p<ي�?�}�%ŏ�lǆ�eK�rsu��넋o��/<��]<Ǽj���� �^�˾p�7}�<'���������Y�rL�H�D�m��3�|�>\l�@f�\:�X��ټt����`x3S��	�:�����ݨ� �./�ڸ�ͻת�����&���}�33{Ӏ+��3.
ONZ6.
���0.�b��t�����u(��fs?�_v$Ȩ�Z��@����6\L1���̙d$��!(��8`�v
�=�]}$fWg�q.��̰�0��:Je3��L�Ƕ�0�W5˻�í��}b���x�?GYǓ�d W���a.vR[���v�o�h�`=��c��jk#臁�e֌���,�6X�x���O���6w]7�����#�]}zik�^/&TZ4٣��M߆�wJ�^�<�s�OT	Z��e ��$�n|9�=^�>"�#��q����BΌ�ο�[g�g%��J\�?�In��+��6A?=�L��D��W�C��_Y �t��4׀��t���Rt����s�:ބ�	E19�0薌�g��M9	�ugv��hǬLOi�����f�2���$���7fqH��+����yO�\Rt޾����T����P)�r�X ��9�dH�
Z��jx�s�#�!r8�ch���%Îf$��P�x�OԽ>���\x������j9����R�|٤呷��27ɫ�\R���{���bb/�f�V�lx56���^D��HH�U԰~Z��E2�N�+*KxH�D�$��X6i�ٳf�k�lO�����#��� ��/�����"��'��`(
C)���`	b�yt�Xһ{�0B"�˔\�l �'$���v��ЊD������fb.�Y<�N�D�,e�q5$;T�/�6�x)���7v�y\��WFW��>�1��|N����fC���]���L�Ԣ��dA��L\- �*���v�ճA�e2��ff��
(Qe�gc�'�"J?�t*�D���:�+�.8��6��q�!� 3��wb����ő�M��ڄ��fa�f��+4y��v8>N��	�x1�ۚ����T�u���;t�d�p9� ՄRj�$y�1�{R�"�Rc�I� �ŊGv�t�v:�^.����H>)�2S��w'�Oc�^A�~&�
�&�� �/$3<���w}�q_�+g}�A��~�����(���5/���&;��I$i���lӯ��
��&����ƺ�'��T�l�?p����P�t�̕��y$���;��Ŵ���)%�/7�/���c�r�C��.�yl�Q4��D��WYf�rE퓷!��\�jIO��Taj���)�f3�@��h�`�Y ��w���g3�E������,�.���)��64TucY�3���en���"Fg#��]�#��u��;j�"�R���Ʀ��N%��51g���A�����z�7t��ʠ��QX�ߛc0�������cc6����U�'����dK;��<���0P�O�s�nc���4n����P]�JR�;p~4|\F����L�!�\\0WR06 �G3C�7�?FJ�I8�;�ս!k>>��b��u,�ZShu��]���Cnz���Y���V�t~]%p�yx�b�*Xv@�'�� rޖ��O6��ӟ>�_T�׫��)��_��u����aۀ���C�Պ��}�,�"�<��UL�"�'�}�bH˞����m)SR��Fþ�Iw����@M�|.�3�� �����X�)��`PO-&��=x�ɑ��:��K��s�fr��|Yv�[[Z�����ܵ|������|)��Z�WH�7�-5�<\�R�9��,� %ˤcd�n�J��J�m3���_�Ek.0���F��G��0�u�>�/;ӣ5�S2;�������}XB�P������=�ǅE�~���-���y����D�>h^��n"Ag�<O�3yR�>nb֠?)��5��1�x�[�F�$���W��)c=֑���$oGWyhu�p�@V��:2G��f�= ��]Y�J4/q�N�%boЏ˲�����O���)�_ ��U�h:�HH_�"�~�|X�(�����4䷃���9����k���)^1ځ	��9dkcsV� w~���=!�&�.=�'���muD�嵝���t<0.���q�H�7W�kXƣ�p�J�'��r�?��%N�Q8���9��e��z�����Vh���*o%��2p;ֳ��ٓ���Z��-�k{�M�BmAGW�dP�ު�)���K1�K�_�Ǔ���twJA]6C�E��h��Pl�պL���,����T�`g��Ұ��\����U�G-�paB���J>�s��{���@�<��5�0F~	����L��O�J�/���������)��J�*;D�nswm��}Bē�����	����]'�}�=�*���k�_uЏ��mm[`��YhU� L�M+b�
�����OOo3��8�%�y�^�)i�8�1��ن�k��0ɪX���M��a��,D���q3a����/O�yFr71��e�����M��� �ݬ	�Ȃ��D���d��b��~�X��OD�RBw����Wz$���n�D��Hſ�U3�N��"u���; =$^��y1T�(���XI�>2��Um�R�,����\�8�๾�
��:����@�L�1Gr|���C�gs��Ñ�M�c��H.�������� ,3�F>흹�J�K�H�G���#til��R�SB�'0q���@��#���>�L��B�#����HG���][�P?B)2~ј�}!)X�z�a�D=[q���fXi�_I�h�<=��d�n*��k���� ��"җ����{Q�$;J��#[e��]^���*��M�m�
��+��@rk3V��\��*N�<���l��(�Kj5�|;~����G��&������ܰH|�5\H�S]H��2t�?Vǈ���E�T�WV�%ޓޥPYW���/u[[�&��H�.F�����^��"���]5�;�U���V�+��`��$ٰ:mo�(_[�O^bL�QEuIZ�������Sn��̔��U���������8��`k�~�6�TLT�7#�0��	p��2�L�\7 ��s-�6|E^�﹈�qT)`��{
Eg��@'ONcL/W��X����&���Z{i��uΞ�_��3	aSr܍��v+�^�ğ�Q8&�֩���w���ҳ����(e����y��6�W�;����T�YM����ɼ&��̝�-/��Ɉ�� _�n������q�i�ZK���<�Jt{Q?�'����*�} X����1BWU	����PY�<�!MH��%�x���Վ3��h�½�0�0���ƙ�����6�	�G��7[����4]��h�������=��r���ϔf��r�C����X���|���z��-gʗ���>v���M�:��DA8ÙrY�3���0�`e0c���]�|>]���L�!�,��?�Q��C��]	�pԲ%<B�*�=�A����W(�	������Sɕ�^ݡx�G��8��a�
f�U���"f��֙�-�f�o���4�ɶ0�K�m8K=�;�S�s��/�H���@�0Ҳ/���>X ��T��Z낙�D�8ı�~���jC^�3M>�i�t�ƥ�[�V��`2�}o��"9X|`ළ������[�9��qr8E�6R��F�?zw�J�1T�֢�=��Z�e��r��˟
�����"�H�D�����i4�S4�������G�����:f�]:�����u��a(���˶!dhlñ��.^ ��#�V�遽�8�j7���1D�$m<(���9ZUg���BY�!�,t¨Ƅ����Q
��.n�J>�-]�)ɡ��X�ћ�]���}�;��m�w��B�$�N�dޯ���k)�pO{�N%�:�w�C��o�u�Qz5�U/����k#�HQ��-�%n��pb�wc�JΕ�ڈ�_xh^j�~�K<����x�<?x� /��7X;:1C{dp���Z�[��l�4@�pa�~Ϧ���R�g�G�����=�o+왮֊=[U����8�:�~��l��j��L�e�=Iפ������E/�y��DY��_�Dvi�����j���5ꁁVsy�G��#���Ο0� ��[��l9*N r����ޛ-��lc���x+��G�s���Z�T��(!h�?�Ue��]�����������1������a�$~�6�d.�<��ۤ�7��d����U��j���ʆ˧[�-z���Օ:$�����rA��[�S�6��T%��ΒUu��w�;��-
iD����JGł���%ߟC@Ki�N�p���˃����H-o�<4$�~hM�½�8����)��l�y��}]�Y3�f���yt��r؉cC���J����e��膱�K6䂅b1���/Z��J�LO:UGao��Y���;p�#M�����r-����*����)\r�����(�����.7��Ҭ)B��ab��k�ub�R�m�I`X(��[A���c��wz�����7�L�AMuT�<l��q�P��G,��� Q�x{�#j���	Pa�O��q0���y>���D�Q7�8YG��Yr�ɭ����\������M;[D����8�V�L�8���#����n"F��J��~4m�/��n�FA��pC�o'�Ѥ�q�S|�%
J�*cXV�;`�����chd&��?���T�e$'g�b`ڊ2��v�*�7O�X��v��މ5���,x�5*����֒�;2\M��'���L�غ:�c���͞V�sX�� N�G�d�	Z�6�������np��4�ˍl���!��#{c�ҒOu��p���Ŧ��,�p���>����ɯ�;���G�,Ӏ�,|
�v(#�w5�u� �)p�3։S���;f,!G�E82W�xe�㌝�W~��>�:�6ܑC��]���-�hĔ�1˰�ԡF��C���;��2٥�9����6)X������d��\97�,A(�N��r������卿�󃴆O���\��~eL�(�e��_<�)�'�{�╃�W%��_C�r���[�	ǧ�X����j����R�R�+��B����{�k��j�'*��rО�)%��?�u�bGq0W�:1���V�飬���p}��5��W�C�c��}v����1^b��l��Ό^Q������}-�u��Z�-���,��m��l�Z��45L����FRm�vR^�I�Dx�B-�`I����=�V���J�e�ޙ]u�ҥ�ZL�{���8^,\RPp�(������N��Y�K�����/A��KF
�pjʐ9��׾<���nyH�Zc�����Si�<�d��n�L��Co�ޣ�����Cz�;��Fu>�>(�B��f0?:�@s`œd��_�B�r�1�e�]� ��ڂ �{D\T<���b��P}�#%5;A�l�Z��m�o�nl�bO鹽1�d����z��������e`^��r����n�����C�Q��y TcȾ�Y��w��i��)kҢ�gÖd�V�
��6,��xX�N�9#�d����N�B�}�HF�A�4e��m�d�4�'�9�bDFq�� ��?]��R.�/7�?H���i���[06�����ma�X�^��y�#w�Ti���j���k=M���~t�I�C��J���q;�y7����.��U.t����8�Şi��9"�������-͝`���x ?�;y��vHHT>,���ǌ~����4������u*�f��+�:� �#\����#���ĝ��*����yr�������f�Ι4�M�++�󟒉\�~���d8���xo�൨��0�u9J%�G*�Y2YPLF�x��cx��4\8<'E%NB�W��0����MnA��}YL�S��=>qV���F����'%�ԝ�R�1_<��ʌ���
\��������gOOUeRjG� S�=a�A���<��R����g^�5������~2����/K�p���S��a8:�l��f�a3{po�������ʤ��/���N൤��_��y9f�,n���y�K����/�!�H�25��0{~_Y��Wc��a�!q�=�Z��D�,P{:��Wռ�Dg���f�����HR��1����U�\5!��f�ۧG��f,�.�r���r�^��Z$b�+�6��oQ^��k�P��_�TX��Q~�t����b�m�5����K��w���椦+�D�̈ds���f(�-��PK&��#�������x�䭝�e{j���I�1�S�4tX�p҅�� �(�Jt�s!W������xh%m� ��r���y԰�|�:�"��Ԉ��e4��荓��;x2���a	mxs
\M�(�	��r�ckU�=��x#��ݟ��Xb��NT��?KБr���x�y"�s�wf:!��cݤb]�m?0����<�x��G�I#�f�5s�L�X�E@�)@l 3`n����������ct}c�:��h9fd����)����1R~ߍ�]j���~=�@�SG�iE;L���+�c`7v#���EP3>�zj?q���xƠ�o�'c*�V��8�OA�`~�> (�~,�Do�]w�����6��F�/�Z��K��
	o���q����n��&F@�Ú&�*�*���L�Ѥ��e|��h�Y���$<A@:�x�$���Va��P%��j�ӛ܎E<����C�ԋ�V,�	��H�[d� ��6𾶱��\�U��0�a�@n蝿��C�3��W{o���ۜ��nS����U2F�x�=!�P\�?l�d�f�ٟe�j�Fo��ν�8��d�ZkjPL���H����g�
�J�}7�QE��^��$9kn9�xP+u#�#G�|�v
U���aPE^�?�1��w�:ܸܰ�˪��P���K��(oz�ϗiDU9He��(S*Ҳ�����Ύ�,��羀mR}f<����U���#_�v-G�D��i�����9����;h�0���)���ܒ��)��o�>Hy�(���m�Mdw���8�b+�ۉ����9ڍ�sXg9���X+�	�?M�N ��05�ȑ�.آz��Fl�bӘl���GTҕ�GZ&��X����1'��5İ�$��黸i�ue�.!�o�U�h6Y����c?Uw=�'�!Q-L~�M2k�R�]O��ِ�O>�q�V<�����^{��N�5?�W��/~��{� _��m���B�'t�7������O������a+�;���R0�h1�W.�0����l�@IøZa���X�����"��V$^b��ʬC&9u'0��(�ݝ?��.#�Z ��2S�����������<�����],4R����1��-j��sa���H�f~cT׉V6dto��8q������\X?���z���-�ۣ�}0t�͕��G����?*�x8�7xӽ����2>&R��u]^5`5�?$�]3�!�B~w�S���u�X�,w�,c|,��>�a�Ȋ1���}�Y�	�Rq�HD�"WM-�� }T�l|8ǫ~�å�$$+C��t9��rʂe��*��-�vD��r��<�&B/�?��uBȻ���!��_�fvB�� ����W+���kT�Z9�ƽ�>Q�)�Sp�f�~��~;,�9V$Ӡ:�@�8�a�	��rT{�q������h��FY=��x^w;�-� 3�# �p�zL��}zl�6�^֎�t���Ycf�%�/���D�1�wxМ�U�HY��%���o�4f�0<u�Q�e;�=�i;��MI*��/n~�[6�7�럱 ���j�>�q�M˧�����&���2ߋKW������q˟�~ҫ�c^��J�\�k�2�wȳ�I71�Ζkq��CƜf�-��!�7N�?�0}��w��Ɨ�O@�
��G����g�|T*�/�C����F�N�V�Ѷ�"�-|N~Ȯ�|�v���FXZ�%nX�:� E�)�H����J�*�[�phoi�_EB�!{�����b��˃�3�4Ƣ�|����g6��@x���uU (J&'}��n��ˍ�5�>��'B��8���<��;1��,�#;]�L%�{��6J�C3X���Nl4��X�й�;��Q$W���n�?�,o�{��(:�`��1����d<+Z.J?�"t(�g1eaɚ5�<��!���/ژ�"�i<������O��5��v��H�ޭVhBl����X�+��N�� k��ofY1i��a��C��/�� 2F
�BY�
"�?�>�9�E�Ĥ�b�!\�BC/ ����s�F=�g���+���;�����6�b>L;��
��*���i³~��X��������@��1)*��LE�T�Ř,��#�l�Ǚs��
v����79Q��-��K�uۆZ��f�m�A������]���lO%�v��
���[�.�� I��EoC5�X~�q������Q���ˁTd���U��E^n#7�r���we�yM&���B��	0F��O7\dd܈�U�Їc�
v=�^�'r{ ��i/��tB����bEy������ ����f�E��ű@E����l� �c9;�Zh4�6��5���r�N�FB����la�7T�u"��ra�^
���~YgM�V���C�:ZOr�8W��JJ퐘ȥV�����W^��.j}���y$@}�#��I'��i/1w�c�fE`r�f�Z��a̭��Ǜ�s4��~�&L"N��Sh�a9�X�����YᏥ�?^�;�+I�f��_=V�@S�(��f&nf/´3���P�����@G/�A?"�U���C'�����B�P�� �:�&RP�J. ���}���U�����D��CXLU҃��qBY?����8����DG����K�_ɑ�����N�b�*҉���������ǝ��(X~�QŹj-Ε^c�G�{|���i�|����M,,�k^�N�R!�F������F��P��6���r1_W0��3����o6���cÉ�l���}"1MPj&|��
G���R��EF�c./��C9�
�����U�/ ��F���ˍ���4n�	ڂ��֊���P�Z&};~������b!��.�aQ��}}҄�}��b��6�!��,Lԅf�!�g����TB;3l�-21����=��o��|t>;����l��y0������Bv��TG�8�&?�Rw�\v�����t�s��fq�M�m���V�	.dE[(����kr�������y(��Ê�x�w�p|����2˹��jbHɋ8D�z긆Čw���D����ו:D�Pw�[���*�]��J[t�|@K��������ա8���Q��.ZCq���ױ�E�bԑȢޘR��~e��g�j�A�(;1Vh�'��嘏}NWms�.�P�t�O�j�ܺS�9����Z]�B�PB����ClB��z��ŋD��ZL��j��tJ�c��̖��H�E/)���%�~����MD^6~�d���f5�_As�絜6ˉ�`\�8��?�˂�����%"����EF�cq����Ѣ�X�6���#_t=��Zf�'Ćq{���oY���jsվ+�������B�m0�o��|aQ����'׌���~'@�M���n�K���~~�H�Le��>Qo��C�l���=K=�>R�����h(P�=�3x�����]���3��h2vQ��Ns{�r3߉/��wi8|�ٳ�TS=^����]5q�p"�|+�X���xNR�5�$L������<����Gin�	[M�x;����e�	�����~�J�Nϻ`}H�Ԋrޏ�l�Ϙ��s��đ���S�"��0~J����"U���ܱ>�h�.�R�D���:o�?w~!�)���k�Ӣ�/^`�a��(��ϧ���*Y2�^Y/{��=I|�l����46!V0��s�S��dف�1#�L�rX��2�P'��F�t���)&�ޒ��ɜI���A,P�>6�G��v`;6Vi�W�VO���sq��:�$�G�k�w���E`�� J���S:� �:q4W_�@�}?u�����D�&&e��*K��6@����S���"3m���k4ְ8�Ȣ���z��Ӕ^��
���܂��73����8�����U�lUZ�*���ti�(Ddbcu��ץs�ݭ�E?z��C�l�z�<��� ��b�N�u~�y����%��ka����aMAW��%����(!猵�xh]�g=I� �ʏ�UZ�r?�;��&��v��������Ѫpx��)��8���7�%�Y�@�,���~�8��Qu�g��k�^=S^*&B�},GP��8W��V�A�g�P2wX�����S�1��ў��X�'�r��O)���IYj��,�# Zgzο��c6N$���qh�Iϻ��;9v��Y�C�`a`�������?�MeZ�:frC���s/�Չ��p�	�.��Ex��?.N=����r͑6�z��/^Z�V�b\�O��X��IQ��	�2��?��w<3G{��L��R�f�q��6\�sxƞ]+w��|�ֺђ�����wd�%9ṱ����y:9-6#�e���t��B���>�j�H����v'��������$�D%��=Fh-}:��gJ��J�d������[�;����R�I�Ӫ�^�m1��I�����rE�3C�)�g����A=�f�>чcK���=3�oˣt�j�F �b_��&C]��U�C���x�C����epٽ,��Υ��-����w��5ĩ���[�N�O� �����6�!ͮ��;z��Y�\�jUD�����L���
k�O�\�%���1�uFS�\ˉnK�)�cR�|k��~��VO)�g�eRp2G�&8�	p�t�'3�3����a�"�ｒ�@�o:'�.y�kX��o�d�����f U���>�/낝��o��3(�)+�p�W�,\����4�2 �j���@O$/��<��%m>��-�1Kj�`�T��g	�A>&̈�[���Ĭ��8�e�hO�rJ_Dkt�R?�I���,�d�N�;��~|u�-�'TB�/�!�t@n�	q��8?N1J�(��	`��:P��lG'Mar�N4�tL����u����%߈��~/L����j^��u�����H�*��|"�����\�A0�k�Kk8����Oΰ�' z�"إvʹ��Z�|���kIIO,�r�ܭS��S������D!�,��p_�3@�0�����ԛ�׬Hk���{l)6��Ra�N����������-��7���@b�����O4.�����FhmmQ~��!@�?K�>��6H��N��c�E̛y�o���j�5���;�����j�Pkn���͉�X[�c��=��-R_k�-���>dU|�+�QA_�~{C�9�Aߣ;2%�j,�R��dwި_Tf���Ȯ�7��Z|�e�Q�l�b�qi�|��W�"ݒi>��}^[�9J����7OŤ,�k��AUD�q�]
ݡ��c	�����7�/t���走k�g���_���K��l��Z�MW
x�����ț��ƃ���'�9�R�_���0{n*��2HZ�/�����≈Jd~~ y�ۦ��r���\�JGG-���Dy���(\�K_��o�AT��e��dk�u�m���6i7^��5�k\�dG�窗��|�",���Bz���C��~(��Oi����*��`7�D��no��Z-|(% i��c4�_6#b��'g��]u���Yؘ���GN2s5�[���yv����D���C2�U�c�s�\#��Śs҆+�M�G�Y?QjJ�M`KgY�+���c��S���0� F��Z S����K �Y.gh齢2��a�]�;M;��#�^�&�K�#��T5zXs&����2W-܋�p���� v�Kʶ�����
ZR��[�Y<�܀���L��@�ϩtJ�s�Ҳ�����r�����8�[YR�����>��4��==)���a���fp�"�<�K�a*����a����ҟ��Q�s�9QVM'���sڑtr��2�Y�kč�o�&h����z�)w��^��<�o�]�v#��"ü�q%`5�G&\v�Z�.���)�ڭtr�A���)�C>�wE�C� ��{4����Ј��Q���W�������D��)a>�Dy `�P��������VB��*�=�^l�㕝�9bX���C�Qu�8C���:�fM3Y<Q�s����v�O:!t:�χ���X��a�W�6g��ҩ��=8F;�P/��>���ph�?,��n$i�0㮧�$sЃ�$��� =:�r��4$*�)Gj������=�5ڢ�D����jvO��u��(�y�01�7иڪ�aqR��]K��>Fb8�5Gx�;�zD:��'l@���}ᐸ����|��Xm��g���������q�y �k��`�1�T@� ���#��R_u����~��b� cN�%#���3e�I,�Yo��t���he���M�*(pBw�;�v�D�Ts52jJC�y�>ҟߺ��5�):��7�<��*��tIN�nz<�����|����@�5��f��� \&����S���e����1�=��.S��h�B䔍z)�є�^�� ��xA�M���y�D 8�R�#�4`}�2�I;�gѬg6:���떶5V�d�_���,xM�he��,��L���IX��z�� tF�b���8�lp�߰�̅e�$團���KJ%C�s��� $R����]�*<��-�SpXF_@q�C���d]x��l�"��w2�8�Mԝ;�2��l�9i~gU�Zr�Xq�ec�A�}b%�+6�?W���_����ɳyG3�4��ď:���;�� ���Ctsmι�R�̌��i�Ր��a�+���I����e?s���eF�+"�Id��|�h}(=�� N;BG��6���B�4���!F\Ի5sxC_ITfk�Zх��	0��w"��<�F�$C���iuaoWg�)W�H�Q��\/����*��R�4_���h�[���j�;�˻9�b6�"+0;��Ƭ�p���g��22C�{�4���Po1�L}�S �-�9ֲܑV��
����_T#�u{�R8����I��O���V��_���Q��܅�,�l� ��36�#���ww_dÁ[3��!s�2;�����\�VC@w�o.n��|�F�6?�8.ׂD�&������4��V2�{щg ���� �X��+$:dנ6	{�y��'��8�D�䘉�^����!��X����bi�@��I������҅�g=6%��8L�Y>�+ֈū�"9�9�5Ƣ�mc��#;�:}�iFqt���M�tԯK��m|u&7 ���23�z���O!>��L�qrI>��M�B��b�m.�cۿ�Տ9Q��>���5��l;�Oz�MJm��񷨂���!}-�K�F��Y��1lA���"u�j2V�G	9L����>��H�i����_�)A`cI��x9!�ؐ{o�|/�!�2���U�~�C�{��`�\�t��u�+�'f�6��A���q1 ��-��Ş����|,����-���H*���V��%�cP�9��kzQ���Mvib����ˏ]yaK�|EA2I��s�%m܏�f✉�X��̝/�P_C�;�HĒ�����Iy�Rq��8������貜�f?��� .���s�_+��ĵ���{��.�lN_\R�ڨ����'�+�zeB�W�i(�������{�uR"�ALd�f�ϙ�m��s�6��e&u��l�@���z'����6'��C��3N#�ѕ�ᒖ]�U�(�$�`A)�/g���=�6YT��� fk���m�������N!kk5Q���'A�2�i����E��(+��N�_A���B�Rv̗*p���&`8 �LB?��@`��)3�˹��Y\��nY:�J����AO��m)s%p�2qd��(����Y��ymTo�v�N��<��p���Z s�|��	��5�E��U���=�l%o����r�v}�4��k$U�^#�+�&�T��~[�ʫ<�J_�u��DsK��\;�����ի�d�4muι�DV ��8�r�x8�AlY�m�HC��s}�kǝ�*��V=��i�+"O���8�
+[zc4W\�C�
BEr�l�Ja��C�#mao��^�?��$,}\Y�.B���N�=h$��\�ϑ ��4+�U7�y��b�|�-�mk�g��noz���o�AE��./zfX>R-�
���
�$�t�����\cwC�VHU��~o���?�p�u(z�	S��UA�w6��%�(\��y��>GLoѝV훽��|���3�x�����3�"]�F&�tj��k�x��T�bJ�y����A� �I�FFL��P�B&@r �e0�6B�X�&L[�d���7"��]�0��4�@�p��qE��-x3�+�is�ў颼���@���'��"T��U>�ڜ��8m�%-|�F���0U=��6|��J����D^�	h��~�n�� ٬u&��������_/�S(�z���M���U��`�$X�}2�z&�qz��喵]�#%}�����7���T�|�¸��В��@����tiK���ۯ�RZo_ۡ�`�}3�I�|��5Es����D�AȘ�4�u��K���i(X�������~z� �t)� M�uQ�&���1C�>f�Z���l%1zݔ$`6��]����PR&W��QPĺ�d��y]�EH���~Ͱ2	��v��1����,α���4�x:�b����!N�p��5p�Q���_�ꖡ�Zw0q�v�Oz"�l������@���Ƶ���RU]g�nD�N
����F�Zᷚ��7H+����:$!dD��ƀ�u|�p5��H�����԰M4�w�wV���,�;�x�_*�FXD��SH�$��`�����)*�������Sf��K�t��§vg�=	c��W��=P�2��%|,'�@�S�Y�\]��A�F���o�92#xQ��//�`��q_6��`�P����*#��D�U�;��}�
͂P��}Q����t�ůKѝK4ͱ&�m�*�x}�P�Rpe)�$)�Րţ{C�'���3�������y�?�᳾^�e%�).ls��ĺ-<%�K�������U��J�#���u�+��������Vs@�Jn}>EE��;Q�<,����jX�ůA"T�:�Ȳs�L���������8|	�]m�GVϊ����s?���,�x����D���R6�bz��^�*^�6(cNi�|>�8��v��P]�|���8;��p��&�S<����#�'����ܰJ�ʕ���f�V�Aj��S4�Y��W����a���Ӧ�8!�z��
�uT�Ê���o��}T�ף�#�I�ơ̴�����}� l�*3!mZv;$Z��^�/����Y�u��DÏA�bi��W$E��Xߪl-a����_TS�\R�(4�!��ݍ2����=�K`�&���Q%>� H'�����$�5�l.V��Ÿ#V�h!q{j���_6��ZU��xɬ�a�qo[Vhj�����Hn��\v�{2K`�� �?+��C�n��	ҽ��5��l����.�>� 	k�p����@������b
��$
J��6֡�[�v.�u������D�����	�m�rx\:yQq#+.������ֳT���a�7
������~1�?[�9s$=8�}M]bS7�q���ga��{m�,��1��aS.�^B�[k�-��A�`ið��<XX�Uk̕	7�}��e��R*�O�=h�ᕓp����wj����N;N�[3C��7�����(�R��1)E�������8�]���Q�9xD_�W��	�I|(�I����ai�����<��B4���v���3\n�^�� .�L���iU���z���%���VE"sj���i馘���|lCB�"�.�����W�ԁ-��ti�=��1�FE!L;[7w�c�JW�HL���?�?�BI.��;�S�G!�@=���Q�������l.W�Ȥ���`\m2n����״�/���?���@��r#;Ϲ3G�/��ɛ̧m��_���WWv7����Ը!f���N�:��7�D��݁J���+�^��~�"v�S�/���Q�i�M?Ǖ�&�
�sa��z����b��K�?�DU�W����4��� ��o�*����>�oeC�S@Ə��>��׃�1��K�����b��;"1*���&�!���4���8��$���90�$�&�p`��&8����*��x�vf���:���e���h,�?4N�5R�%s�c�<���T���67�"ϲ v�}.�}FX3���'�.gs�zk(0Ԡ���ݧ�L�8�Dq�q�́C�0iŭ$p�r�Nj���{8H��IE�!$�&t�G�Q�����w˹���kh����*V�=%�*=e��Z��w>O�}�f�S��A��cI4��W�#ŭ���q���W��Q�����t���3��CW�i��&�	_rrʆ7��#!�4|�u��ٹ6,��pU�H�fRm��
>�^(jr�cP�����p���{�Ag�E�(������OZsy�Nvy_m��' "����k�����H���ԻV��t�q��^VNk@�v���HYy�a�|l��Suu�A�h��- g���<�6��Zc�0�����wBrԼ���0q�ǰ	�U�sƂlx4^�h
�T�B����u�X�W1+�LE�Q�vyY	_9�'v��t���\X⌡�Q��9ј"�׭y4�3I�Ὼd(�?�kGe��d3|�-����n>}7�R>7r�o��o;���P��cu{�M�X�������CМ���|�t�j��c�S��|���c�������:�N�'#�~Lx���2��R�����05����Ӆm�C�=�+^�)'�~Β�ݧ�$F �����e� /y�'�]��L�}׉�?��Z!�mΎq�R�&K`��yG�i:�\^�d��rٺu����y^X!Z�Fn�!�Z�Nu�Z1�鱌8a��/���_c��{�f%[+�_0��gQ���U���^�p�ϙEXۉ����-Nh�֒�e4Pt��F�r���_!�f���"�/_"�5�4�1!�L0�����Mh�4�"�S���=�_���k��0�� s�A�f3��}�C���8C6|Rv�֓��#Ny�������2�!�r���v�t3n�m
��m 'aܴ�x�ٔj�5\W��궍�6[�zw�����h"�O�{z�sJ+[��\&�Q�^F���z,n�i�/�j�N��5��Q���f+�Ek������Zɭ�SX������?<�S?.�X {`��=��U���{TcC�
�(P%W�@�(}��R2��Z5�vv�A,iߪ����� �؃��J�D3�h5��;ghZS¯��hI���s:���ᥙ"�p	ϵ��r\8(��Y��n7'n�?FtK,�x�H�����Ȇ�[t�Se��݆�Z�#���*��H�%�)Ye]�κ`�.�x�0������`S;�B�qd[V�%'�nP���ɮ�N�	��+�V�(㙆������
B�����W[6	�2t�/%�dRMX�Q��j�]8����*�D��X�>
8�h��c}&S�Yi���;C�A:mAE�~Q0�'��4�~���j=���f��� �*�,@L��C
A�r���yKq��5��R3�(9�
�o6=��[(��]Z�s^�1���lC5���emkM[���+��u��b�]'J��ctʙ�.e;A&%Q"@�]˦H������#Pq&�̾Z�N�}��wǡh��@X�Wڪ�t�|*�ՂxfBYET��O����t����kȖ`#I;ԅ�$��x��3���r|���>I΂&S����z�][P�����;[��z���B�E�ht����1}�
?P�q-�N�(u�F��JY-(�	����Oƿ�ĕ��)��E�^�d�v���h�_��\B��u�O���*T���G�,�!sR�N<�E����#6��������*�Ȇ]��Z�#���hE��k�b8�|�u|���i�[{�xU�'�����!Z1�e������"sy�t�J��R젲o�qA�X|�(S�k��Q��i0��9�mBK�H�?����G���ӻ��d�"��~��-�M����\��,Mч�xE9=�M��.�P	�<�����A��6f&-��յ���)��VIx�1�&��ῖ-M���~m�W�mN�Lה�t�O u7Ic�.������k9D�8���U���l�l3a�W���-�O�Yh��Zq��9OS���
x{'�A�d�OSZS�����e������y�%N�o8PJ~o����v��#��J����8�(pH�Y�w!��~��k&y&�7�������g�N�f�{ ���Q<e��$�ZCy׹�Zƹ�`�]v�/P��-Օc�7m~�*K��گ5z�����<��}ոQ�QU��e]�)�������U'���`��56��ͳ	��J��Ǹ�'�ᢟ�!���l5�]���5�o8�&׃Pa\��i���Oխ3�[���U(�M��
�\]�=���_1������Wy0՞�z� ����7��Oj��ϛ�"���!y��ƕ�Ue��_n(��kM\lu,*>nkǣ0��C����D��_y5\$
��fĔ7ѰOE��5/�%N�*KZ�z�ii[�>f�}>|^T����{�$>wV�-\�S�;��q	K�4l<T@�a���Rױ�~H!�<���-O;<T��˩ � ��v)�{�:WE_��<�f�ެٞ	8|f�xp��a%�x�)v9���z�rH�4ӲXM�&Շ*#΋��`;���I����3�O�e󅢡P�pT�ޙ��!7��c�����!�Nhϛ(����#�ή�/�zE�t[	H@��6�u��Q�!y4��}\���9ͺ퀼�z
�qv�p�4�[��]Q9{X����iX������hdo��7A��y6�:][S���k#��O��*��^}9�1t���S:�{�\��������"sv˹�}&`�'R4p,�#"5l��g2]!���ܗ}I�?Ǽ���]����rh�U�k@6b�0�'��0Pl��r���Zi�T8y��c%ƫ+R�nd����Y{.��t�薭�M�E��# �]�3/�m���T�Y�K�sA�qh�����2����Ι�)�G1��RCԊA,�f@EU��,ŊU9@�<��CR��o=`B�����e�ˬ6��)�晗�駸bK�o h�đ��'cj=j�ճ�����oj��~ �Z�3C량��Ɣ���鏖�	�e{��%t�j��o]�
�" ���{�_�S�+��d��� 
��z5U��P0������R�j
�+hhP�c������[���EO��${�/�z���<��b � \�� �;q/w�{�2W��g�d��ml�N�k�m�?h<h���|����ăY�9g��\���[:�7l���o�		�[�@vZ����FIK0�o��_D��#38f��`;��䏵��(n���)+�p�u��ŧ^h�t���)��Pa�V���6�3M��Jܟq�o*'vNQ�/�{v�F/2/��Jb��,|7#�&�7��o�`(W�Z0��/��13�8�;�e��x��X�B�[�E.Т�?xh�Wl�VZH�\h���*p�L5St�����|��ј�E�݈O,79*�¶,Q�n��xH�Hmn��d\f�*�C�����l?�J3���/� ����F��5yȳ��3_��ͅ�����٧N%B�'w��� ���4�*ؽ/��K�N��>�IR�L|��_����tA�"�}����O$.P�BW4uTi������u7���
!I��]Q�L�_2���ʢ�����Z�~p͖�"=�����@x��J�u�Z�|�w�tG+����K��\�����K���E�!�L}��$���2H�3U&E���@y��P�}�%����l���4%�Cq �6�e����R@^�X���y /+�h���`� �¯L>�~��,D�<��S�.Ҥ}��T%;t�8,%b��+bm�5�\%�W�}������@���L��:}M�� ǻ�7����9L�������22���Ø#���uu��M;�R2t����	��l��h9Y�����o4f�nc<���o����2��(�������r\~�p���	�I�lZM'p�ֿ.݅Y�8$��5�'�X�Q{�h���O���/�c�ё�����60�|ޗEG}����P6S�)���O�0{��gK-wۻk��ǵ_��e��;M�T��� �����%�ѰFC�9�K��6�@�M�_B|~M2�s؛�t�|�,�6�^Y�?��h��\�p?U�h�|��9��9��@��"�P���Î�@�{Er���Q�P1�u��v�T6{���5���Q��΋EC��{ĆO�~E������ýo�D��t!P���V����u6�g�Q����{�n���H��]��N=�Hj��a�5|#���j���X
sƬ�E��AF�񔸠�|_X��GtZA��G���@�V��}r?��?yJhk���Vw�^���a\���
P!U���`X���"_����8Պ>d�fU�� \*	`�}G��~Ż�V��jt��p��z&:�h�hTnsq.�����G0%hF	�9f<b�Z$�i�7�G����Ji٢b7e3�l��iM��X�Ѿ�j#G4D���������]��˘�>�m5�5�`��#���$�=ʅ+����j�l�L�A�Ɯn��үߜ6�=4kf�c�S�"QS�����U�;�o�t����*��\�S�˟k��60V��kĜ�AF���"�s(i�c&��F>��+k�u���!>1�V��
�]̓�/?���GH���?gz4E���F���i9a�b�Q�:���s账�-yv^��o�%���n���Wq�P)��^K ��E܎�۷^uo&���|���H*�A(���x4���������T}H�<]O|�^FVNa���qFA�5��4���^�R���y]��L_�<9������~�'DM���<G��X:�2/Ce�v�E�$�������E޷N4qG�4O�Y3���<��]�Y�a�Oi]:U�+<z��:ig�W$����3Ei�(EXY�Hn�`'�.��U!��Z���o��@O3�<T��InH����^�E�ٽ�e_̰$\���E�]�=�a��o��^	��/N�H��`�ᨰ>��77�3Ӱ�_�G.f4���C��~^�,utӮ�s������ȡ�\^el(�2q@�b�H&�ձ�2,��ڵ�|΢�Ǫ�]6c�,���L��༑�� �k�^SGw'N{ �l�������̯w��f�P�T�V����_QO/#���Q �gV�*�,{GS;J�1�$v
,�Ap��Nm���a�QB]�Sv���v�Y����$i�� |Q�q<F_�L�_�[#c�ՠ���4�3Ub�gJQY�R��-J���堇�3Q��t��ܑ9����x"`��iZ�,1��bX,{�rI&w�5�c����t^���,c�!}���C��7/���{����[�v��v���]�1��hw�X6r#$��NY��_�,��v]ܭEfM����bo�y&-�s�L�o%������]#�V�l$͐=X?��A|txd��6��i|�:�[�a��W�\�z��ӳ���*���1X\��Uy�Ń+7H.����[�lt7��5��6��;-�"����[�O��"ȿ7�h�KK��>ɤ�TY~䜼��M?̸E�|���fΒ��	�ݟ�^���l�p'N���WNZ����6��X�j"�r.�����,P��f브X >D���SO�k��-�+G*�P���_�J4�Ro��`�����qIN���!,bї*
~77b�S��4~*>/mX'�V��1����q9N"�	��0sy��������@�:R�G�`�}������|�:����)0��R"Gg�=��4O˼	UN"��d,��|D�X��~��UtsلG�'1�r�ē�`��k>���=��ˋ��EZ�����]H'@x飆>�_"8(�HE�#��K!���7�~��|t�X�2�=�j�yS,iO�i0]�m�>�I*�$�.	K�z�B>��^-C�#P��uݹҘ�i{�QiX�6ùޔ�G�'�-B��|[�XF8�cm��cەO����Ii����#���a��t�/�Y�dpK��h�L�+@+c}�!�	g�ٴC�+�~�߰u���w_��.�Jp�1W���tM]�Gs��q�M�5oD?�'/���V���(4��v�y��^��[Ivk���i��0_�L�8���˹���,�=��<C!l���]ؑD�W���/��^�PQ*��k!�[�d�'d)t��Oo�^��[o�%XSA���Du����u��\*R*0���^AR�	�F��.r7�%Q*>3�+'^����I����[�|i \i�����t��v���F[	���#�K�Kv�� j�9�h���;���z*Fh�I�Y����m$�Z�b+��ӉO��,�e��:��C���VX^��'�N�p�/Ze���ف�c�37l�{Si��Qg\�!�ġ|J\��P|��5+�6~(���{��!O�x}�6�~�+�J�����{TM(��sVd�����5t��/��+^�8��xհ8�}�l�������9�]eu�5��{,lFu��aǧS�"�[\%L��ɞ��*��V�UKX�$��O)�2�u��*0bB��7M
�S'���+�Ct	¾�����[�5��s炦r� �pV��g������m��j�����]Y��K�M&A�ď�ƕ+�@�x�(�z��_z�#3(y9�1v�_�Ǖ��ʊ�KϓK�&��Ѿ��K������a�h�lQ�ao~�_mC�p����]N�*�_^>��(���<��xEs�V��X��2�*�@�4���f��δ��qʇ�H.�
yC�N��E&[�]�!?ʟn��Ǎq��E��o�s*u�y�W�]U!��;T�D�s���@)�s⃳8b#D����p��w��;#3��؄:�R��[�@M�A����R�Q�fD�b/�}��'B:�c���f<���^���s�A"r�^�z"��,��L������]���7X��#�.�[�P���� ��f��P�iR�C�R@j$ ��w��I�7��C�4�6��ɠ�9;M ��Q-��=t��/�y���o��`�^f����<?�� ��/�w	Vy�g��#�	�U��/�[�UK���!�u�HV����1}���c���]
6!��Ctl'�e����B/%ie��4l�M���5�b�����LBNXpՋ3	M��QΖn����#���-7�oR"
�(��8t��u����֟~�A��x�V��Yp�h���U$+c�j+]=/��aҥ���q����g�KP�&t��ʦ�
��%dA`��%�ES!��������FdL�`��N2CI�����r7M����MG�Ƃ@�O*U3��u�sܠ��� DoF�C���Z*� ��)�T\��E��z� ���+��	���������x[�[2:Ȍ�˧!	�+:P��{M���Y�8����E����V�p�s���L��u��63�Q@g�y���/�Zw��ܨn�:�B�ew��T+17�v;����j���0�� ��䔣ݿ��,K{��e�w�W{�5��BP�y�V+�Q
q���:5�˂��
�J��DQ˖Q`�Vm[*#Q}Rfr0���������KX`��z\g����ߘ^d�R/HD� 	L���K�ߜ�B����A6���R��5,q�a�P�i������d`�.�he�@յ֌�1��%�߿u^.�κxZu��Y{��A�1]�"�L.�YEa���KE�m.>��a�Y�U��n��5�9*���
�d-!ɛ�Dk���xRM��y��L�����U++�{3�q�9)8��0��E�����?�b���\��:�cc�L��9Ѷ��֑�3$������?��s?<T�/yPD6���B�V"z��M�Cc԰��R��c��`@�
��(��E�Cq�f��!���w�"
~�ؗ�J{�;쫒j�x�환;��X�,|�I�8�M��?7�.ޛ�{e�Ui#~�3,�H.c*;��[��3$�+ć2�h�f|�[Q���W"P��M7ր)^����Dt����\B��Ķq��'��9����ڌ��F����tv=�\���w��\�f��LJ?�]5ݯ�.F�	�5�23}�]�
�T륈��m�9�>&Ɨ.�P��7/����2�+���h�>(��2y,�髺�XF�e+�����������]��|Q�۩w �k\����5��"IiR<7.ՄɂP,��N�����8���3�f8�]�0��KH�Qh�&e�����v�(ݞ�k��{�$�2��+��xhQrE�,�Y�zd*7V�]�������}N]S��3�D�ܓ� �r!ީ_wj5����j�ď�0YF��3�.f!�}�����p���"��H���ee/�@�d��Z�n2�ט��"v|xg:��$�n{�o��d@c_L�{wņ=���R��J��9�����L����r�3e�%3��j�"��X4�|g~�9��-@n�����1���Q���q!/2"G��Kl�/�ya�=C=q��#���%� ����\��|mP;�d�8�:^�hC�*�3��E
�ga^W�wb�@��7��~!ou����m�}3_n�Ӓ�E�r��ӶGؠe�ú�cI�>F�$�X=9�(��U��^.y��;٦R�ʑoٰ҄$�w�k>��Qq���SN��C98�a���: ���v�'���q&r7N�u1���8��9X�ݵ�����L�W_�I��Gٞ�|�pܬ��$̙}:{�[GQ�@�fƉ��)��6X�h5
�th�]Z3��J�2���Y�'+E`"��D�u��eb�G'���PY9��7X�7u�.�y�Zi�8�|�e�S��lY�r;w���'�yS3�^T���l�ö�S���?l�xgH&A����`��[�]�9�����"Y��/8=�@�};m�Y�4�N
�ퟄ[(u�dCG!UEloF����}sŸ��f���ʑ�wV�x���$�BI�
�B����U�-�'8W:�y>Ə
��T=h�큡ے�m��7�v���Z�ôAa
4V�z.��5=J����RJь!�٩�)�����vW�*�����Nail�[#D�L��^�żC��y.���eN��BN&焈��$��rV�ԙ����DM�h�Hڞ�8�!�2��~�0?y����'2�4���=G�݀�Qm;)�&��&C��k�����	�+dq�Tm 9��r��	����7���|q�gwT���Zg|���:K����;��H�s�y���f�?�'�W]<Ƹ	�~H�\. 4��6�/�c���44��#��`�a)h�[V�*Z}n�����a�<�j�|�3s��m�f���I�c�')>��&$�[����W�S�x�Ri���a9V�:�r��Y%��41��XQM�(TS�n�=��Uk�IA;PҢ�ѥL$F6��0���B���q�� �߅Xn��7�%NѢ�[k�q
�n~mi*��˗��Ag�k_�N��2?�xh�~
rˠm
Y�{3��p��B7Vwҡ��Vm]��#�����z��(�]���o��G�����:Z%^I���&nvQ��H�0oH
��՗l^�Zj�Q^���i�^�*��C���h�c�r9�U��W^G�[q�p}H�q�v�"?��ރ�q�n=���O&3כ�A��ȹ�K)���>���:h�
����,���=�����js3�%%~���*�UJ�᭚_7��$�Q_�����d,���]�Չ�5s�A2���o���:�f��v����F����$-6�mxе$�eЮ̝����0�h�&�/i��<.`\�b#b��1K�9%��&����-P���p8&P�D�ߘ�������@b��=8�a�fdɣh�@���̈'R�Mm�<����8��?�P��m|)�=�'�|o�����U%v�v؊��]�eyWY�.���ɆZ=xLDܟ#�"uā�.�� ��GNtBt��rR{�B��f\aT�28�7:����p����n�V�Ֆ�./w��-�c�>b��@�SDG*��X�P�$V����X����] A��U���"uj��6Y㾳b�,)�t�D@&ӼE�0B{�p��/�6��b;R���򊃖߯�gHO���/��H���$�%Aşz\����vc*)}Dx]�5Z�0з;�]$���E�s{:,�dagX����ۄ�]n�!�a8g#A	��9�( A=��!0m�Ip��Y�n/�I=.�[�}S�fq?�J=Z䢫����+9��d㺹���i�0�?�ؽ|��}E͘��{-�I�l�xܚ{9��A�u����FV����+����3���4y.�vz��l�x'���,:LpSE5Irv=��ͅ��{�f��~`SmA�	�9j���Ά��B[.�gZ��Ñmܕ�q'~��+����~-{�IϘ3%��iZ��� �	�Rƫ��z���f�lK#�e)���J}j�ZN^�ZCQ3��R�xfP�5��~`{cHSIJ�N���Ӗ�Z�N�$ߧ����m/�~_�E�_��C�\�=8%j��+xŅF"����7Nb����kH9� ��N���&}ͧ�x�b�����q������h(�B�t0S*��� �OA�L��1�;7svO	\_;��T$�m̡Jk&3����(ɡx��-�9�{��ո��T/�d<xt��1��%�]��E�y��ic�t��I�|�Ҽ�-��8E�#h`�i�� S�����ͫLD���a�ro�)<O���H��?_��5��� G���U�B52vm�ƅ���}���8S�p9z�� �0g���УW���=iwY����#��cϴ!&�#�Ɣ݅���~�|c������(ICXe�?�Zl�(����H�����eV�\y��"͗�6Yx�j:Z\>��@�7�Y�e��ȂbS�܅��b7�]� � ꧳�����,�+E �Y��>�+4x�5�&$ꀚ����~�a���`ᖓ�OF�CGt�0���od�����Q�,�����p"��h^��yn��y5��@�x`��4� �P�,o8���P����56��{�X�'�v�iOB�.����2�Rp5�� �����Q`��,�����a6�b�Ū&�Uz�	ah�K�O�6b�6������1_��E�'{��JL۬�l�aj�0R�z[��b{>E�*t!w��%܇�8�=�!���ʌ	��봄��)���q�i�5��7��T^����E.fl��� 	��d���qD����u��{�� ��~9� 4�K��P�k�蛽�����a/eu��֦�G߄1#�J���݅�3h�C�k�x�׫C���I�5Ҋ6���\m��[x�Ӯk��g��	���hBfv�.�U��MI`�}ɴ�r˅�^1�q��-�0�;S������W8�_,\#Zu�T)|�.d�+��~�)hB���A`�2Kdf�㻉��Ӳ��?"�t@��+�}�������-���`�XTߐ�jl�XK��!� P iF�`	Yq�᚞jYF����d�u���!���u�xZ��]��l]�h��X����ѣ�M9�˫�d�R��T���g��܏�O�[���	������I�0�Y��u�����Efz�1��}b�%)8˗}�������S��le�Mׯd
0Їo��K��\��r4-5q;
<�A����~�>�f���ێ��dc��'�aO���Fdz���=^]\�X<�rmb��\6?�+٪ۈL����.U , ��H>4,��we��I��E�-�w˹O���e<0���d���ohՒ}1��|��;8V �dJ&K.F��n(\ˈ��<q��2��p�[���'�6-����n6�F9jR�njN�4PC<MՓ�I��#��K9��e6��訃j�s}��־Y
��_�����K�l�B���U�hY��'�v�()J�@١�GS�)#��6;�A�[.�vT��	-Rb�B,3ǋW��� ����o�?�m��c�������O�w c�=I��J�X��E��:�ͬ�b����>�(�!�r����ޜeb�dr�}L��?����j�UՆg:2� �l2C������E'綺����7��L�',��;�.�L�:v��N��^׳����un�h#T��:����5iq��@765£ �s���R(h��!��"^P�<3?�U�;f�r=2F�n,+\Emv�#pG2A�gw� O��$p�Y��f9�����+�^�/��:��HW�>�ȮM+�ٝ\b���1�w�=N��-wi��e41N�a�8���O 7�H��
0�C��0|R�&�R�q�D��m�Ӽi1l)����(�f݁TɤZӻEz���5ʬA��]�����M��)_}X�De�fؠ�f(9�qӗ��WO횤�(��Rg	�_�H{�
�x(�X�I�9`����]�`�yo�)2sb9f&IR�p���{$Z�0����o�����-���ʣ�"󢜏^Z���q���&�n�J{@`��[}G�v�@�ӹq<�7 ņmIʨ�3�)#C�	��9�ZxA�ӑuqS�z��ؿ����=�Ƶ-�Vf�����Y��҃/ܣ�9v6֐am	���{��+d�=�P䎂�*��Nt���p8&"��h$�?5�q�.�Kawݘ�|G�}ajr2g� �����υ�������[��*f��j�X�	��g��/�A7�����Z����Y{rCt�CvR��rU�ݎ��Ȇ�:]�j[�R�&ӕ��`�Q����V�x�XH$%�\��q������R�b/|��ܶ�q?�~,��\�̕
�ϫQ~|:�B>�񾹣����g�v/�&^�	��70�(�W�[���f|�dA��HR�;cg?07ܾ��_�����<���k��-j���k�Q4hq7z�<��z��J�QY���x"wRY��!Ű�mɯ��B7�E�T��>C˟B辣��}�������Ϭ(^ґ��Ϛ��Ck?헤X�v������N��^I:���uR�ȴi�;���Pܮ<��Q#Ӛ��%Ͳ��{�I��� y��O�e��!d�nU~}2���߬.����H{MBY�i�PhF>϶���{���bq�ϡI�%���*�M��h�58��쀞��J1�Oٺ�
BK�g�L|O4͚i�?	zX�g���
�5�a��+@�H����)����mIDv����-�H]�FE���X5(Ψ���'��M/����ᶻ��ә�Fes5|����)�jt������L[�N�{�#ł��+���qDz��Jz@d�o}�`�?��ʤ�<�D����G!�E)��K������j���椑����+	�J�p�����/GX�?m�$>i��O�ޑ�+�tUb�2�H(P�ѷ���.�̓�[����?`Ee��2��	S��h����������y�"�Ɨڮ��;��T�|�S$f�4EP���oC�$}sj���e��e+ky�{w�{K�244ǂ;��2�|��Y���;��!JA�1*�(@��xQ;]��h�P���1E�&1���t_>�J���
���'�UIQ�S�U�W��%�11����0� 7�u�?&�k\U�-�C�70W�$���>��HZ����3vG��������ֻ�R͎נ�p!8�C���a=i�$#���8���>������n��*7���)������=���b�K�Zz� ���T^Kw�� ��>�Q���(�σ��h��:�p�S?BB��Yc��3N��#^#f[���KORS�1����cf[<�|�:�t���&�?@7�ߕ=)���U��a��\�ێ]g|N^�	�Qg�id���>�I����?��VE�-Y����3�f���\.��	�s ����w�[tͺ=�O|vh���a��.��PT�z�Ϭ]/�`�i��f�LP�uj������4�li�Zs)�k������s�vQM��0�!a�,�h�*g�=����'Q$��>�9C��LT$�H��n�F�ˡ�2��B�#]�"���E5�]�|Q+���I�&1Ǭ�Bh�64���$8���p��3�c�3������Q�p� e��m�e�6��;V��V;���%�cG�l������lfJ[�K���C���W7�)4I��KNL8����uSg"_X�Y�b{t�������XP[�Ӝ�b� �2�|C`U#+������t@Fd�!)6���j�+Yn����}�۫=��5���5�r\Z��| ����a��+咓9d��6���#᜺n�ė��Gk��6֠��,As�A�©yLVJ;��������M)dQ���IG'�ڼv0�#]I����gn_K�~5R��E��:�i��Q���gAl�@F�vѾA%�R��
��?��ry�8�Pn{�����FwRT0;C{9�w���Jx�z�4�m�]�����jzn��þ�H��:��N~|���w=t�{�-3t��T$������I�"�B��9&�����A������pf�@LT��3��H�i�����!��WI�?!���E�,AD�$�fa��}Xp_Z�Xd㷖��W4no+B��7̀��Ӏ�c����$��ʺ���|ck��j^�
�������+կ�Z�wl��?'9�Lq�>&CGW�V��3���=BXY�{�.���ը04qh?�#�^�D��h�;�m~2R�B?�H[�mz�dR���F��5Љ*Y��mxvct�>1L΋7B6��J�s�>xw#:�������K�"?ik]�^�&GA�O@�;�jm�<@@�;j���
ȷ2�>Ue*-J6�����%A#�)�E��p+q�1���#b�ɠ@ǫfe[֯ $��%�*h��)�k�R�o��32��D��4�8m�� �Rօ�;�PM�Yf��^O�Y�EpR�&����&\ �j��3�w7i�>�|(���MS�P)ZT���֙ʗ��W!I�W4�����p��U,^�%���A�Z���X���{�W��܄s�:�DU-���3��<���#�4���Z��>+j!��u�9��b;�wX�Lg``J�q����< m�m�S�(��.#+���j�Թ�r	Zې:Q>��^}ro�4�_֝������8
X��_��5���A:4V]�Ԙ�@�y�PX�4]kD�P ���Z'��\"`g��g��F-���?�i^Kg�<���~<�9)�B��u�:Or�9<l�r"�eTؿ+�&-/D�;C.<�#�@��
��4W'|�^����6[@
�P�85L�%���v�:~��4��r����Q͜E?��R��k�{6�/3��S%4����7h�pU���Xz��X�0ّҶZ�0#�$^�"nօ�p�1u�ȘE^+_�p/8��^w����E������H����\?ȕY�{��I�NB��2-����&�XH|���`�_��R��9�x�Z��,��]~K7ADMh�gC�G+���v-*�{�A�I���D��I��g��蟦X��Et���g%�C� ����o9c�,"�7�+���2�Tv!�I_Wo�R�88%7�� f�89`�;�8�!j��P�izģ�yqVF#e�!OG�%&�1l��*��6�?��FDg/�4-�7��=�4��S�Q�.�j�x���[��p^=9�b��s������Y�%���d�<�8:%�^&�z�.�Nm�'/�0=�[�uj!��}Ƌ�}F��D��,��!Tg�q���3a<�Ŧa*���QM7eږ�}j����}�&F��������������+�1)'\��. +t��e�pa=�n�}>!}����2*�Q���e_J�@���)���^�ys�t��=�5�G������ ��>�i�w�"�[���W^{�:�Օ� +h�����Q	�JE���%V�mA ��ץ�m.wt�J�/� S|��������<�Y�����n�	^��G|�䰶3�&h��4�����i ��~�P�v�]a�B	����iO��E�Hc\�TU5-��m����|�o%[{�յ8��X��P���p����{�=�3{uO!�ՖRc��m�G�s����X}7 �.�D��6�r�<�4N�dx�ZZ*�2<-ĸ��]%�.LTHc��X7��*���h|9��yS�����؜&�z�el��YD��x~)��8���o�'r��a����E�%L�.^7~��fau�طa�-_:mKHu�u��]pO�3��o�]�CP��E�#St�/�� `w��p���o��),&z�`Pj�%~_���e�r���hl�~N"���O��e��6�}�s�O:�Iv-��]y���)�FdW3կ�/SfR{^tC:u�!g0`�>?�f�1��W��.�y3ͥi�'�S��+s��"4m����|^"{P�t� �X����_4�Y��oJ|]�&��N��D�zzg�O��.և�+��J�������m�F���6�4�9VB�'��'�T��8zz�^����	��M{d�x��y둙ꯟ����mC�i�,g�+0��,���bp0����{����KG�Oʤf��L���d�f��qe_��mT0"iZ��W VY<�_�q�^���P5�J�u�%؍6��P<�!�@\5Q�ڧd������B���kP�|�����.�O��)��k�;����Z!�$���I�c��f�(�7q���NL*���,w�	L�E��8���A�6������O;I��I�<+������|��oM-��\۹���
`�4��+}�}��3G@�7��}\dLp��im?�(�3j�]�T1]��u���gr�<����9N0`1&c$�e��@���Zr�((J�BTѨ��.GQQ���N./`U$�א������F�ʚT�|�l5뮻�4��UU+:���Q��+�����QgŁR7j��0�߈���Q�����~�{+|^%�{�N#���'!������^y�wH�5U����+����3>:�����D�J]+�Q��3r���@�=�pErǨ2�ÿb���!������L�:���ɱV�b�9`�;�������!R8r��j����ג<ս���Z:63ӗ������G�&I�v�A�:5<'�ߪ5��.�ݽ�<��T!����1ɶ���Nǈ[�	��g�4n�\7t��;Η�p׽=�#���4B��'�s�L��z�r3��L������\�HM���w��M��bRJp��TpNr&ࣥ-?������3z�m"	�Z-��%���fvC�a�o��)e'�ep?���>�:�� � ��K�Tُ�#�o�;��#��g���Εe��,��eŚ���6�L&%�Z�s��:��v���+m�I���J*i�F���8��3�+`;�W0c������>�& �]��lr0J*c������z��%Ç��w�
T�JQ�⢳�R��mKT!�4=�kî��lY�͕C��.���3jm9ku���;g�������-�����]� ��X�x��iu��MDh��U�U�2RP<����LT`��\�̘
���!���SV�5�>�3���h�@	.�>,�u8��V�ֈ5�l��V�������/Z��u`5�#KJ�~��|S� )e�`���]��,��7SqB��G��<�&T�� A�$%�+]h��c�L�V��x¯����,o>})>���{֣#vQ� 5�;h�@����g��l`2Ǔce ���Z2�F�:��8.�(���݉�z1@l�է8�㽺��� ?�,xa.��NU���{,��.����O'�L�5Ⱥ5�J�-��,W䛁��T+D�W,яPl/cvrC�=Y�4����G3tjn��^���D���c�<��BL���ݷֲ��]��1
�y�庛�YT��3���4 �T�	���d���)�C=`�$�2���aAUf��g����庫82�O�����A\p�BC�r�����h��d.�)�!�S�V��26�?4A
�٦E뫆���q�J���k	��D�P��e?,�ƫ�G�?�dB��Cs�؉���R������AqՑ��ǭ�}����߲�B6���cX=y�?	�w
f�b�k���[�@8���m���N�"�˳�LY�X��q�OG/�T��#Re2'����o�GzP5�-:�����=.�FW�=1y]Qi��.{���D����?����50�.Y ��gMJ�� �d'Á$F�� �3Ť	:��겱�)-���f)��Ot?�%:����B���\	6���S�����ӏ��i3(Ꙏ���/�O��-�<�qlf��βz�I�ػ�%+�ޱda5O���L���"/N�7bh`� <ɷ�����f�h(�Q���M ��\�t�KE�B s=��q�ق0�Ә�me�n����޸HS�>��[t������(1��+/ᦼ��N|��1,�?���q��&����Z;.��z
�t��z޻�b����7d��ߪ���Ha1'�]�}h��F���],��*��1Έ�~�M���:ש ���6t?��h�l��O���8;�Q�����o��?�wzg��EŒ��K�7S��bZ5��.�cso��K�(�Q`��������HS|���0�+Y�r��ԫDjx<�����0:m���9�
�
�@��a�h�M+��>���<&����"J�i�n :��sFXx�?���x8?I�E��z��u_�B�!i�jC���^�/�.����!����p� x�s��b���lE���5�&�b��hS��@�30J3y2@�$3��H��N�@z�W�z�&�[#�W_��U���j𩂲[oc����z{P/��4;s�r�R���|�{��#�|L_��)F��*݂E�ه�h;i��{���6�.
���nNc-+h"v4�9���LA�t��ԁQ�c)D��3?�\�[�M��=�ꌺ��m&cS�������ZP^�Gk���ggA�?�;�.���e��DY� zԷ״I�8�F-խ�;Bq�dK�"6)y�H�Y���h���+�̧� �F���W�������2�M�Y@Yu/��8��?q��RQ4@�F������⳴�}	���U<?<%P�i~5!D�x�2@j��P�8��*۞~�u�����@Q�v#`K��2��K�4�H8�OehC��{F��x[/�e>}ϐ�ղ��!.��faaswp�Hq�!����d��^V�)N+I�3M3	��6�)�J	Mh&���89�|��Ei����|DU�a�w��-
�����w?��3D��c��F��.3��p
髬���Vj��ǒpx��M���Iu�yK:����p<&�*�(r�P�ǴR�;��>7e�Yz���|��)|`;�01�6V.�Ft'��F��[��(b��t��IR�H���S�>�po�k���Q*�/ۀ�hcCEl���o�n��8�� niK�NÑSg1��)���pO���i^��-v��J�2�.G<,��|�K�gDu����X���7��ֵ��S4=��M�z��Ce���L�D n���f�iD��
�v�g�hMoTd�^�m"��^m��l�k������I��*�>	o�� q�C�Te�F�H������tj��:[�a����v�K����SP��A��q��#Y�؊Ł>�7_iiԫ�9��΅�0�����P5����;Ιt`����;%��������6Y��4��\�1Tw�sɌ�G˥�B��,��ˁ�0guf���,7]��c�ɛp�r��?�a�>�����"��R#���f*��ˍ�`<�G�}.�L&���{�=aP�/�4@�TЈ9(.U��QBm��@ �Z"��͍�]��r��"%{��%�J�cn�pLٌƢ�
����Jt&�g�x"6����#�6\vUt}���]8�����t�c/%���S�+��\ޟ�B1� ��;��N�!65#}���4F1E>�Sd�}�����'��i3P���L��K�טG}��s�O�藂D掃��b]t���(���%��"��ql�,Yq��/%3�QG J����{'�%Fh�AS�@��S ��,Lp$)4u�M%� erRa\�j�G-�Z�Nκ %���}I&���j �/J�O
v��h���+���b�O���(Vq3�#w�X���W��r�;��em����&��N�3TpAX����|N�x��I��3Ѷ��*�)f��p�1�O�d��*|��f1$�7Ʌ_��1������IPj�pKDMńPkh2(����u���!��_ڷ�� 'A@�+�`�'���n�.eKͺ�k1&'U��b��=b�l�C��
�Nb��c ���� ��䍙R���q>Q:�'oh*��*f^�bX�h���4�>��z��-)�~��'����R�����x�?�8ڤ�?aon����uO��ba�/�k$�c��G��:��}�⫾�����>��a���*;[�	7�NM�h��l���B�J{fwu��E�U���7+��9����!cZ��vn�N�_�"*b��k��P�Kl�3��!�f5�}���J{1� ��`c��#��G�Ή����8r�q�����Y���(>0��W ��旵��E���mT��7yv<\U]*#��2@q�C��q�ŌF��EXa> ��.�PG��������8%�s�2V�>����G��HJ̅�<�l��Y������%-�̭ ��_g��B�.,#�KAu���jb�኱
V�]M�y�?��p�u,KLS��|,���r��9��bl&�\Z�H�i�at�
���C���Sx9.���Ü�>����L�����[�>]��F'	�5�G����5����]�B��[o�ߡ��`!�{Oh�36�����_B�Fj'�7e���-|�\8���0��f�Q(�keB_�����j� ��͜P_%�I5��"�֭�9؉5�A��$�tiw��)_�{�mgLբ`k#E����#>M}3Ǌ����H����:�����[l���}r�JG����B
b�P���p� Z�	C��1>����U����|���:��k����$� ��h��	����n	��e\��2� �+�t�u{t( �ǜ�-ɔ�q~)h��[���+�_�57���9	�tV�7���k`��'��O�P&���<��d���ҭ�|��h?K����ax�M��C���`�G���j���,�TQ��e�O�E�m�����Rr8��A�Hq�>ԕ��-���E,��d G�0�K�ul��Rm|�Ӡ��9��z}��XՌ!��*>�O�C�r�)|��U\��7�CAȜg��S��9Gi�e�X��J��8/�t����5r��-��b��b¤�{�T�j��&�]�,bL�&���~a7_��oDڄ^!�F�����j���{�.2G5&�J��䴜>�w�J�8Dx�����ͻ&s��p�Y᥀�7�/~e�����p�ɼ�.�cln��-@�zȋF��>�D���i�Ը w~��0 W9��>'yKxq�����D�ԅ�Ք$�|آ�+�(������0;���w�w���8������_q��1����w�C�&��T�*?ҋL�D�bԔ���g��Q�j6��.a�FDTƈ]W��˅��]����lʎ�*!1)@]'f*����G'�4��=^zg�/D�Q�I�kc홋� S!POg�U�� �}���->>X�Qvo�jOk)�t�P���s ��>_M@���R��ժ����J�)k�;�E	�P��)w���F&�ʵ�q�P�{h|%6�����'�mCmM��@]5m���]@]�I��5ӀA�ȘIb�(�)��뿜gn�ѷ�B�!�:/˙BJ�X�,��|�&���P�.�2�0ȡ����(�z�Q<&�j�9V�U*��W@�G	TO�ǲʿ���@J��U�۫1Y60��rۓ	�ܜ6��U;K�$�;�ne�$7:@4�ǘTxx���N'�8�1^Ƴ4^����?5�m���R���>�&,.�ʪ�#�ZxGK�|3��x���]�c�XS�'[������B��o�_ψY�S����@�|����Z���p���5�2w��ˉ����h�z����Rr��+O�F��e	��}��҇�z�)纮���%:U�n���:C(��˔Iu�����p�TjP��ɀPiw�� "�<���$������$�/�&l)��U#YC��Ot��ϐ'�n��@v;����z8�+��-�~5�^������ܲ�p��J���O���s
Ǒ#l��g4��:Kk���+s
n:��!�=�4C�>Џjcx�&1����7Թ���2z�����ɿ̃Sؑ�|5DE5����6�6V���Q����7?���L�E�n�<�vњ�������e���������L뗂��xU��C��t1�y��;1+נ��QO���6�8	�+ߠ�HYN\Z�ǹ�ɬ�.?�%����qF�L��!�y���nq%��=o��e�L����֗�6�(�:�Q�o�UM��`��p��@�u���#ۘJz�o��J��NB�1�J�Ǭ�-�W��X�0k�l�Ku�%�Y���ʆ�~9������l�@@z�8�q7��c�X��m�����q4RգVk�+g�&�>�x�ѥ��|�u����这��"���	U�h{^����%ʆa.x��jU�SG"12S
c�n�=@F�R��ŉph��3�ѡI:�H434�i(��g�����U�VUE]O䷂��8�s�%^.F�_��,�.�o�m��'4�ϝP�L�b�30G}��17�{m�ӄ�Zg���-\�Ȣc�PB�{�}D�t�w�+bsG _�0t'��}0�-�]C������[�z�z&�|��H��c������3	iU�������bM�w�޶L�쳻��Ա��Gm&YC�;�ՖW�_�.���!=��e�{ʜ���[��n�yr�BFAw�p��*��ِ��O+�3�W\[�w��WV8��c&��y�H�Ҍ��7U?�Ku#�����b?Z��9��e��'�]#=�`���w�2T��2O��{,��q�
��T|�e\���Ίu��|b}��{�Q[k$ۭ��a2Q>�G"R�;d�3t�7��\[�����*9C�;���6���[�f����1���~��oՌ`�\]v�f4(��V.V.���2uŇy������}Z��"#1\���e���הD#	�5އ��۩ٶ�u�A��M��[��mhӅ(���Ks=[�mJ���VZ��[K�rK#̥�0��$�丌)�E0�^��!��O�݉Zt6�����گlV�=G��Sw����	ŋZ�9ֻ;j3��|���G�0�����mڲdߢ���w<iα	�O��H���*�?��M-ǴVFh���ʻVM΅B�QK�U�S�3�fW/m�֘�����'si,�f-��t�ůJ\*|4�"fG���O��)C�(�M�X�*�$�Q`~����8�n�L���Er������n܏O����/��g����s���bR��)�C��vh�&�y�aD�g�@s�j��q:�Ϗ�����)!�؋�\��k��]��}��JNF�D�[�^e�R��?�S�� �{��o#�&���osѡnk���ՓH2��rC�& Q	��6����sc#�x@�۶�Zm���D7,+�*1�otCiIL�#~;��͕�SNS]hN�!������B���D e�R �IH�����ѷp�g�i`��E�e�|ɰ-�>�1���u�?��m0��y$d9Eu�*\�a�z�Ծ٪|T�Q��ՠ$�W�p�=�0�w�פJV<�b����Y��D���qlt��ir����]K#���14A����m�'i�K�UUĺ��?�ڐ�����II�b��xq�b��g��NR>ڏ��g����>��: w0x#�_Wn�~����J��l�yl�f����'���3~G�)�$��F�*�<���Gć�ͼ6�8���h�j�U�4�PV�5�����%)����l��JI�v�N�V"���<�6�y"����������>?W�z���~=<'��P�a���Ǟw�����S�4%�eS�AnJ�$�.��<RE,Fl��&"|�N�<$�F��+ߥV��˅�B�Q:Q{D�(��}�E�zd�L���w�\�g����>J$�F]���tǍ����V��=C����ty�&#��]��qi�[8 Y��sM���LU�!�*����?����j�ū�%��bO�,��ף���F�i�=h���TDi%�.4;�ی����s�{*A�r};X+�])q�P�D���^�)?o������ݰ��Y6ՌD},��LV:i8F)Cz4��I���7zG(Gz�Fmp���nt~ߗ��}��[�$~�%\Bp��[�C(3�W}�	֊��V����5��������}�����H�^+��G���v�3I[R?nD�7�Y~l����&%����'��p�mC�4,� U���^��\��E�m^�|���_'������gRF���]9G�^�5Z�y�}�P{���IRĬ��x 7>O������'O���AF��ݪ;�²)
0.D����m���᧙y�8���Cۥ��x��Á�ir�c����E�X��v'��PA��/��"!S���U#,��C�n+X#f9�@����<�vP�Q�N��
Mm3*�[6�Y��)��w��[�&�J�uz�H>�+�m�WY��z����5c�0�*U}����x�W]㜅=�{����u�Bia:����4�!���/�e��q�ܨ䪚�OR���S7�'��7�+�-88s�o 4N�B�:���
�@�k I���J���E��c[���E��w@M��٠���m+��&� �b:;
�u�ޱ��TPW�'���՟Tn{Zm�!$]"s�NOc� �3�tW���3��bMm ~�{y§6��qa˳��9"oԁl�&�A���~-JMⱳ0�����`6�#{�0-n����~U�$E�˄�!ʱ`�r��^�*\&��!ˇ���M���e�ZĘ�{��t��S�Fb���7��A�����^���u
���-�!ץ<��8�����j�@I�0��D���d�\P��!Ca�8�x��S<������m:i]\s1I��O�4�%�`Nb�3���l�<L���2ҳ;y���%U"�9��
7׷:���)q�e�W/����'*:Z�^��	w{l��b�p�n�][� �iM5��8n��w��D`�b����徛0��MMbx�ħ���ְ��6F�G�8�o��yF .q\h��U��-M���lY���S�U���ڀ.���j��6*�g��P�\g���Z���5%z�M�"A�m��F��@�X�D�x9�����x�!��x�زT#�^�6�i�]��}`N����j�k�=��)� \�qGr��g�������+��s�
�cG�Эθ�B$�T��N�M�c���@�̄/�����������4�Dnpj�3�q�Y9��Np Ԫ.2y3����6�W�"܇$�z������  ����$�e @�M'�iN7�[�-a�z������tL�wq���ˎ6��"��c}��)��R�M+�nN�r>�3f�����U���P�76��0f�	�Q��V��'w�s���cA�|	:��UW�]D.]����T�%��lMX(�Hq�m(���35�bخz�P�����^[ߊ<f��r�b@G�2�8}cb��$��4�I3;�y�KɚΛ�>��/��K���R�/���x�+�	8�nf�$y����}�slZ^�e��3l�!�rfzFV	�D��?�f�*��]��,_o��pIK�bۯ���v�N}����C|�v��p��v=ޑάF�X��2�9	[`�$�g�I�GƤw�aK3v�z�ӛ�9VC��w(ʷvi��<��B��ۤ��a�J0A7��׉�
��W�(��K��M�����6ݚM+a@�x�Fy��(p}���/�Y���\[/Ϥ1np4lϓҒ�^�i�T�>�Exg������zX9��.d�/.̆��n��o��00VY�c��p��J�����!#��W#���a��/�GNg	����}�9��of����U���-�՚hφf#6	:�G�n����������|�f0^�>�~e6.}�WW.�]�К�?Fk�D,}��g8���W��Bw��h$FrR�|0�D��$�r<�;��U��Zو�Һ��N�{�����Ϣf��0t�u�\�F	�ұ���(���e}续�<UWEȡ�^��LQϠ������CTW�'��F�u��r�N'���x3^)�b<�PJ�*���QU�RA*
����AF��!���5�x6}���3�6+�����&ư����1����K���_�[�����d�Q:R�����I����=�-��C�.�u}�6I�-:g�!�򋷃��ެj
1�c-å,D=.�r`�*��Q�s���l"�>`eY�S߿��ʛ���Ӟ{:Y]����Yx���{M�ŵݬD%��\egDP����aq��c�~�d���F�@l�9�ӌ)KU�HLǾ�w��n�1X[U��^N	0��t�0�P���������i���|��6F�i75����}��<�|1���<5z"�I�rÅ������]ĕp~$d׆��G��b�7ar�z�6���V匐�d��$�O��lP��-C.B�'0�`�[��U��nFހ���H�Q�w��n
�bY𥶖��#����/�Jo=1��[�p�ͣztܦj�����yg8��cR���I�6#QJZI5I��8�b<G+*�R�~�#�ޱ�%�ة��oy�*ch��3���\�{�8M�u!y��E��z�F<�4�ڞ*nUw+E���O5YE� AL���p��P�ux˜�v�����J4!+!p@$7B�8���-�V���c3~I��p'+.�'?h����b�)�>�ns.��k&́z�# �w�p��R	�o��B�������Ӄ�Rɽ��%������_����{��g�����#�P�k �ꊪW��jSS�:�y�Ǝ�m�!��}���1S-���Fawnp�K�7�h�����, E��ҳmO��_������ �B��J��{̟�|Z^�2��]M+���Gz���#&�W��[���A/ݏ��>�j�W���Φ�r����[;M�L��ۜ�F������Ն3�`��S���+���G6$B�k�h�ZU���{�PpIZ��j�`�(*�&E6�]&�K����m��`�!�5�����ғ�c��/oz�N7��~����f_m��y����`��ã"�FL�Η*:OS<W�zH�Z:|u�˹�]��ʧ���X�����G�ue ��/QX���+;�N�x��>`�P1�3��wn��l}��&L�<{�hr�X�X�A����L��V��Ϳࢅ����!"��+��6O�g�¸�m��O���*ZL�����rzi�Qh<����|�WnV�?�튰ϑrToiI�2/W�
����}#���b���iQMC�
�q�w �gv��}�
��,olD
�٢���Hh�+k��<�>�� �C����®��£���+H��%y�-)	ֵ�S�i|e� �y�u��yv~׷��Z�x�2�����k;;oT�5{�7oQ��_5E�f���ۯ�����w� �a�R�8ԢU.�'Q����J�6g�x����3��̓s#��m��C����.{Λ��*������m��V+<�[n�e݆� �I��F�r-]�(9�$>���B�2%������Q�m5�^∦�"�2��VM��L�y�-r�4��o�N/��JXy���/@m5�P:�ajB��l���D��B�Nd{�ן�..��X|���B{�䭶�>��]E.��F!g��$8
�] �;Y=��2 ��CebL���y��<˵���ː��̝̹	kؓc�z-6>���kZ����+<�RRP��R�?�Xj�����um���j�Ĉ��r�Դ��j��)c� �)5�|����xU0�`�3%BTQ�h7�kuz�:�0�Z~k9��7�Hv���.���k0����J��Z^�r�S<+�j���'`�t�-�|x����ӷ��W�їY�y"���v����.֚ϓ��Z�r?G��Q�8�]r|�yx�0$�Bѿ7���h���5�,�"R}�ݾ7X�t�W<X�?�]2��[�Fw8I�Hx��uI��o�c�*�V/��zB#�@s�nm+�<w<���D�շ����T��$g4^��}.�S2S�����0}�XE�H-{���j�H����'���kX�|QuXJ�/m�]c�~e�n�"V_�`k�/��[�����q�io}�sMs(��j����cCV�s0���l0�j��;�,��oRmXn�y+��)֫>��
E�Du�ju�?8�{�"�����C�	�q��Y4r�NL�>�:�]7���d��xe��&t�N�� d��Qd`�;���$�H8�D/z3n��}K_���#��eȓ�}��M�#I������ގ,��K��]�N�xCW�ӷ���Gk��!4*�#�����j�|��$�Z�#�QC�T�1l*LY�šՠ�oPo�����CJ"	X�
S�?�.��S�pm5't�7GPv�6D�a�K��ޱ�Q0\�̛ᆎ��H���KO�V\}r�?�취�����>Xr���o�au��2��A۩��	�{٘➪@݄*���nVMbD*�O62���v�hikF�aXДÜ�F��5���z蛞���z����u��}�3�����e1�i�8�h��_�f+W�8U"\H߉dJ�]j��D�X���e3��H�b/�S�xz�[i��Es�6Tc�>3��:
G);X��J�ەK�ʾO�,��Q��c�H��b�}Ĵ�U_�zx�Ԑ[�Fv$�l�u�=�&������W�n�B�/������Ꞗ�-at��!;�w���Ø�Q]2�emzS�o�v!uчH8s�*k�����g�gB�0�&�q�������&��.)��$f�Ź�o�T8�m��ˮ�?��\�֢:K��|
޽P�b���׮UTY���G��U�m:Xx����)ۃ��DoC.<�#{&K@�/�9A�Y���VD*K7�w(Ϩ �6b��Gu �OR ��B��37�fKWo�ؕo����}�$¡���/ב�J�<�	2�� yZ�I ����`p�k�x�~���2N�I���)��b^�/�
o��y�_�4��)�� �A�W�@�E��f@CU��]���ݺ�,�W�J�^d���Bh�\���?8��p�՗�f#?���\����IH���B�	e|Q��)+c'7P_���E"�NG�Ϳ�Մ9��F^�v��$U9�,�W�����Ї6j�%�C��԰�o������6?�^��R��_{�*8g��R��I��Ta�.<�f�&���l|X����n��ڼ���<L?
������ӆ7�}��?��a`!eY�nw�]�9��k�r �üˣ1���� a�#kPfly����8���<Q�w"�>�e2'�<̛e��l�7��ȁ��IF\�(4����x+��ˎϽ���<u��,��WV>�fǲ"h1yɻ�}�A>�,�0;Y��L.���CS���$��P�v$byK�3� �\Q���>���k]��'oRL��Х����~����6�ˣՅ��m<��� �>�P ���17��R��� ѻ�xe` i��w�K���/��ϲmo�F�yRk�8�S�j��z$����vW5� |2tn��ڂ�A<�x�եؘ�JiO��h^���ڜ%��q}���ozlI��eOC0n�U���D�\���֨�����|wz�\},��{{�s�O�����q��!�����W��(���Q��-�;2�Ӎ[�>2��b�$.�on6��f�':�0vv�Z�������'��E~/ j(���S��z;V)��V1���3h����͌>�w�����!��Pf�&ִ�b�30�Q�������pؖ�_�4.��E�O��HuE�n����Sl)�Z$��XƌXȰ�G�;&Ϟ����NB�nc����5�3�����KۛJ�m��]v`źZ m�G���RJ	�c�sӆG��<�]V�.�����)�8�$�nߴ~�=�)�Tf���,��T�{�Н`"_���R��_!�q��{);|x�ɍ?�Ù�RON?״�=�X�y`�[�e��Y�(̮w9�ubCװL@I�<K��UňZZSs�T��50�JE�s�}Zo��X�n�6pȈk�gY�-���&�}��/�}��+5��0���pf�^&�����.�X�N�a���:4�b���q��2��8�°���h�˭�����ʁ���)�[įq���"$�?YTg-v��JHj���� 'P<u���4�%�j�kW]�el�L�ӢoLQ���	hX�.}�x�o#�����$>���ɀ����w"S���vwd[M�i	�Dlr��F�;I�{p�E������*ƌ�b'��n7�+~9��`��;~����gL�.R"���&`|L�$�k�����{CT<߾��8�M�c>V�&����H����|TBCaAj� ��8\{P��o4^A��� �DU2�;\�c�S���TO���1���6����V���d�zI�g�G�`��D7_�]�QE�<�X[E�iU ����o~�i�!���ʡ�DG;�w���R>�ζL�fB�(u�W]�$�� rP��q7T���+D�C��ޱ�<-Tq�T��9��Q�j��muX�R�)�k;��sa�1�Dd���C��?O�� ��;�Ǫ��3R=��Y� D�B�;�vj��N3��+sζ����V�.)��HN�����lj�Z�o��ny��?$A�$�Փ@�����������Y�g��W��#E��|��ǳ�Y����~�n(�DO�3;�E�֘ô0A��Ux߫^r�:�����!�f�����AҦ+��s-��[���by۷� �w`�6�_,(r!�hk���0%�B��Gy�Q�B����j
�z��	q�f11�|ٯxj�Y��"Ő�簆qG|yB�_�v|�>oN���5;�;�����B���Sz�p\��c�W�&�/�u��4���A�+򟾥�ɧ	��
��A@���`�r�U'K��}��Ny������>Pv|bQf���ˬE�#s���_���m��
���r�lFf�ς �M��b���?Oǣ��l����O�G"J_��Ml8Y,�8�hA�iU9�Պ���:��o��--��s�IN�x6@a}�^b����� ��s/�p�멖:��/<�v�M�T��1{kk~w<_��aYi���ە�u���8b�ڸ��z����E��gyi��P&(!m�br�p�1�]�1�(��?�W����uq��%b鉂�&8�`5��;{��W���z\�Y�n��UI��P��k�)%N��H�2������~i�'ٶ����4�edn����'�y�FyE�u�Bo�JG��@����I�Բ�YD`J/���AkA|Z_p�Q��O��~��_�M4`�%��_x4_����O���ާ-)�o�^�?���3�l81��F)��j[���)e���n�ƕ�X���{z����u�yn��;w�����d�{º�����Q@�o�U���R>�"�J  ܴ1y��t�1�݂ΟJs/]���#:Z��*ScI@��k��U�S(��:�+�R����C j�������,�M�tڭ��x"����?8Ƌ�yk���K�������M�b6��+mߑ	p(��8�H1w�r�bgr9�Oo�_H�c�'�Z���<.�s_��X�p%{��I��Ɠ�`O����5tIKQ�ſ�]HL�X����k� EfȨ�O��k�H�|fo����b��2Ӡ��9R,��_a���	x�rh��dA���PS���F3Y"��0���
��䚳���T*UA�*��5�A+��X��O������kq+�y�[��?�,簎CS�8�MĪ�E�ܺ�2�L�^IEJ�֓Н��5(��e9�p.�p�o\O����P �峋��N;u��é����1�A4�λ�b-�������l�c8*Pq?2��p�E�N)G�x��R���A��إ�7a��~AJȈ��uC�L�V������"[�v����Qi����K���}��R�]o�oS�ܾ�7���`w���bؗH6zG��xi�6Vzm]g��DJ�b�����OH��D76��Q1f�����,ާubBK+0�S���Ė<{rH�1i�H��f$���/9��.|*l&�_���RR�9t>��/�E��^i��Z�]��-eƍ���G�1�l���(�L�'��t]B.YG��s���m�M�,8�ȥ
�ւ�#�!L�nR�&#��@O,`����J@���$kSM��1·Фn����Ʈ��gru��;����%��/NU*Z�_�C_���Q�D2d=_X�ӝ��C�2űūQb����>-�z1t�!Ĭ�@�7e���n*>4�"k}�c	�"�q<O���������ks;����o	�AQ�曦Ԭ}q�+�����Ж�\I�FxG7� v�G�E���bC�G����Y �Z���+�O}
�Ma�8N�3����^:�2�:K�w��-Nԛ����_3��oD���Os�ꕑ��l�G�`�yQT��륰V���yJ߹��p���4&�P��{�b*�6�f��w� �>d°SK�Q��;1�3���Y���5�1V\g'����(������ /ʬ3C	�����?0���v��!�,îxH?n���>��ۙ��/�G�>�|�3��0t��Te�&Sy{�����!�t���1�����������#�G4@;�c1�$��T~|O��5�?9���gh����WJ�q� \��6^�]���ߥ�/�D�dQ5�+]�)�;;�������2_���-�L��,����!$"����Q����pg�z�}�FbN,�Fg�8����(";�q�su'��(W%<$17c�����q/��Ͻ��}1zQLwu��ͤ�!K<Z��j��׷>� #��
p֢QS�w[1��ԢQ2�\.�D�O�¿��u>���=�X��!^\ґP��X�r���N~ �U�B�I�8�aoP]ӓ��Tx���0�&�\�z�K�+�����?�����╊��y+ �)�G��A�����vT����K�Rp�f�̘�.��84ʣ�?{�C�[�S�y�.�hߖZI����In8AzW�>�L|�h{`'j=}.p6A��.�A� '*\�\u[��4L�O~K���?�/��I�;3���z��G<9�\M=�����Hz!)���u���.B��gGJz�1����� ����CH�٠hX�S�D�rTy�EY!`A���˧9�U���Ht���8�,O`�C
ޘih���$�5�I߽T?��/?7��@��Eq/j{}Y�u?��y�鑢�[����c��Y©�U3�q&_E�.Ϗ4��48��o���y>/E��e�4<��d$�?��­�?\�rV\FP�X[\i8��Oz��_�[��F��:�Ђ��'o9�Q�S�MJW�z;�ɖӎ�kU���Q(�@=c1ۯ�����!�G!m�m���Ztl��,�?ྈ+{+�c?��_��>^@�����ߨ�`�ʿ�Kը0�gN���*�u�6
���Y	o��6�D(8�rI=]���k�P�����hXw�N>�a��P��D���?�z`����416:|��mw���+���l��l����b2��UJu����j��v�`N�Sk�����fe�#�1��Ý���&��v���lLZ�E��^p^6W/�\B���w^�j�\�aJ���2]�����i��n�|�������P]�2Ø0(�#k��}���(�\yI܉$���x逴8���ƹZ��R]�g�Լ��D��V+�"�B��[,Υ������}�-�;:��q̣�s���4wV��#*H::�KP6v�{?-O�C��>��8��
n�^�� ���đ�XX1F��g��FI2t��=atk��`GNnX^�X!����g�8�̀-��^Ә�\x{9�]g�i�-��}�jz������r-�(kv���L�����tr�Q�0�x�xunm��@Z3��iw��Z%һ�C:��׵{K���G�(qd$m��s�a鍌��9`�K� �جߧg\L����F���3�c�xv�X~���ɢp��xѩ��ϸ�CE�� ��zB��K���4DS��-�	r���z�̶@Ŝ�4�����K�!K�8�<�;o늞x����,���&N��=�e�z�1�� ��9���L|K�GDo��F�:[;�������e�j�;� �k��2r�P�R���ߕw*B��O ����xA����@���w���"
Nl�v�ɩ�n<Yб�辠�ؗ�fW��3,s���DL���sn��t$�$�Ա��;��C�N.Q1/I~'�t�T\�I#ɔ�����QZ��N�@�N0��!�,��}�@���Ͽ�PT��Q�b����0��+��~*��:�8�Nn�iO�z
��I���z��>�?���}��!J?W���Z:���j�w?�;ld��"[u:�~U�/���H!X��ź�x���k�nX
�����0����n;�����X�5���o�Hdd�,j��fdc��j�V�<�Z��.�;�711���D&-�c�ڨ�;���$|/�A<W |(H#Zm��#����ld�R�4��p�*�{�`��Ʉ��6V�''��M���QҐE�[3�|����b�2���;�}��k4���dٖn��졧���(��[�8����E �I��V�Xn����A�p�<�L��fW�u]��!������{¥3�	!���æ��y��f?n6�Q[Q���"6��|_�3L��є�n�Pxw�ӓW�&}2G	,�m�^h�����+�M(�˯mS�aF���o�	��-󩕼=��9�*�A�;zc��+@��E�$c@ةCU��_=Kq�j2Y7��P�b
߄�3��@���h�:�-&��(��$���N��GRG�^ON��x(�K�(����%r�ȍt�!�������l>F��h��3�yS�0����!QR�ݓ�ɏ���H}-R�.3�N��I4�a\ӹ?��ѓ�*����c8��ᰒW�h�QV������m>��q����/��qLs5���C���IÞՂ勐E�%��!$�
*��u�~�����l�]HG���]�,���B"`�)$�����u���~2�@����2�d$���) �+��/��z�:Y��6�|�ZV���m��M��/�(����>I�����_Z�t��V7�S'�/����f=&@z�ս?L���Y�s�9V
]J~N��ͥ���YRZ�BD(�w�>��e��"�,�G��V�����S�p�I4^�b��e���[�ׂ��K��5I����"�KП�aGcb��N{*�����Ը7G�S�k���#�ڸ��4�R;a���z�Av��!Sx�V ʑ|]h6{\�V���h{����4����U�U�>kN��[Q���^�M���U��Q�L��&��cj�4�i`a��]�#N$s��������W�]�	a���^�N[T�hи��m֪�(u7�{�p�dǓ�J����cz9K�>�&2�V.�'\λɰδ��Q�� �H����3[C�tȚ��<Jf�Q��}��VU��ڹ��ʐ(1P�wف}.1-��u��]����QS��n7�[ 0=���.ڦ�h�a�D�D0��K�Xh�����p2y�۟���+���k�5-4
QZdrˏ7�H_�|�Հ�]�ɡ��RQE�gޤWt!� ��5Jicr���=����j�`Ư!�fO�;6��R��%gH0����}�sF~�\@���������-`�Q���*�pt68?��{�˧0����f������p���lm���LO`�st�]�&�]��D�Dx�*�4��W9��9��W+�p)�MFK���;bd5>�A}3&��T^�E(�<�k#�󆈆��ͩ�� �[!Pb@tW���Y�Z����.4V9���"V욑fe<|M��Sr,	2/�2�G|lju�{�,:�=X�3Z���xI*B�F5H�%�X�����[�Y��:	��j���u��'��������TD��E���1����=g�TB�#�9!��Q4L5�8�!��󲠗�X�א	8�'�%�����,��E��	��&1��Ǖ��̮��x���:��PGh����@_}���ê5Տ��~�i�7�z��V�T����ڦnI��b�Pz��(�V��8�}��"��C= 8�ߚ�����ǉ����%x��u��k�|n�0Y�L��ڴ?Ag�#��էw�@���^+��*>�QD�e;^�h]��f�p��%x,�DQTt�S%��P�jSaR���o#~F�%��-�ZU>��`�"�0���-2��ZDds���#˛qS��J��'�G��4�<��(�>�b ���<fh�ym�����W���rB��-4�q�}e|��l��A{� S�׫���	�αa$�ډְ6�9]R�y��96ݪ�4|�eF�82�V��q����X�z&�|�S�Q�..c����M��{M���<ȴ`�T<�i�#���E�:hG[2��z%s���Se�qU����a�^&�w�Gd��+�E��F�fVA���-��<m�����bN=��'�ƶ��=Ru\*��f�u��
�v��hw�B(�A�vb��d���\䆨�J�ׄ��P�S����=��B��i	�l���T @�����rH��� u
��4*�\ZS$��D\�3�m@e.��D��*3ǛNA���x����Yx�i�!A��,+�������ŕ�~	�'8��j��8Լ��YNuKFpkg(O	U����X%����Nx���S�C4W�|���m�s���n�ř<�Fn�/l�{|��ȃ����CpVo��O��!���@B��S� L@hX�Jl������=�劥�_v'���B-�p�P�"�:��'+~�S��q���� GJ�c��h.�?2����/��]^E���o���y���$���3�^Ov��1%[�qMh���#}������dAԑMؓ~-7��PzOS�3#�m�B�EU{H\uh�Cu���B�ʔ�۳ͣ���4~����J+��S�",)bg2����حX�ދ�3�c�u�#��8>�bT���)F�|��Ex|���A���3>�~P���˺kï:�_�#PQ�?ʂ5Tx@4��q4�o�7�픡�zU)=C�&�a�*h�pA~�L� �#
�����;�l8nQ�s������]��4���T��M�(	�
W|���q(H<!Rw�P��j�ۘ��Q�x��w�!6L z�ua"ł�j�3�B&>��h��p +�f�εP���^+Z~$�!�n_H7p1�	:qDwN
��	�c�ă
�F�c�?��R��iw�Ԯվ�K7��y�"LCI����G�>j�Hn�vf��u�AGj�KFC=�5�R���r���)�E��u�,ʁbbT�猃����y�8�T����y�i��nj�$��Wbh(�I��t���|�A�W^���a�� Et� 6J�E��1Ȕr� �g�R��f-.����,y����1Z�[jٖzs�����J_�O�uF��ir�����D���)�L9���K���y���)��.}$�@ec�rB�k�@��x��{U`���|�NKl�[y����=F6�^N�?(3�b��e�|�Z�6�V��:�>�G�$��b��<<l�W�z��m����\���O�F��ѳ9�,X�C��	1���)E�M�1 ��W�5���O�^Q�����tv��[�(�Yݾ	�F��yEEC�u��<���A���cH,�;!=*�5aI5���v3�[:�L�G��۞ǌK��\v�
Τ����9���#����a��jFe�aMʬb��� �7&�2��`�s��K��_���r=V��F���)+�/��Ot����j����hD̂���#`�د�t�#ӴuE0�L/G>��c�4^7q_�B�F��H�"cJjv�=X՗��x	��L��>\z>Us���Pj�T͛������;8� �;�k�Ѣ�4�u�$�~s����H���E���1@�t}���%��ar�ŉ^J�a�n�l�|u�$x
Ϡч�z��>k7�������I��}%C͠ub���O�ȼ���iP���}Nw�4wj�)+�1��.�E�8��;����d0Ѱ����5@�:w��ü�o����l�b���-MO|� �ƥ,hw�Ycԙ6K����jT�8�Qf�w=)�O�hf'��A����iU�Aݹ��6ܧ��47�e���!�s�+��^R�|jy�
	�]�})��X�s��)"��Ir��k��xɹ#��Ȑ�Hd��,q#�Zr4�Ŝ|r(��̟?_d�|u�1F��t���f\ǋyP�Z����d"@��SV}P�)㜡��Ȋn?�Eҳ5����nf�P^&'ކrn�*��bo�)l
��ع��u7�E[Z'ߏv��D���$�����D���{�D>�� ,��	��z��d�9
��M<��h�k���B��TH������ÀT�E3�B'�m� *�ҠZ87���)���F���۶�_�{���&��9rd�Qk8a��ڐ�-�!�X����IKR����[�W:m$�6U��@�Y�a���҉�Q���G~�_�U�m ��ػ��{ҡp}`�T�i݈��۷�߬�'�"����gNɭ�8q�#Jdt�z��b�yuFD�{+�p��ddm�K�Ն���3�!P���E|�6���0�`�R�5���!
���쮙�@RE8��[Z�.���*s��G`F�aռ�tx1��d]B�G�\�fb�R�Xƈ�t� �񯊚�/�xsŋ	:��:ڀ�^>�4��z��S��"��m���Ɯ�:D�՟Y���Z)�٤i��_���Zy >��k`p�<-�~���$�st-���T���+�ڀ�����<�,��E.>�-�8n�w�aQ��.�ZH\���/��TҬ5�jI��L4c��P[��p���P�pˬ!����z��Y,�����JV��w�)_.��8��/���1ޥ7�f��(<+;��x�v�`�E"���(��!���f.����EJޭBϏֆb�8W��� �,�G�Θ1n)֯q"�j�y��/#K2����2$]%p��dQ���GVq�f�!��B����9<�.����'�E���ќU4` �Y�{��߁7��1��}�?`��^A$K�(�b�z:���CTa����J�B�e,�(�ҏ2�>Nɓr� _p����Ŗ�ND^XUQ'�m�g�R�^�^v��3z4Fç��}��Ћ�(^ru����a?>�i�"�T�3ب�D�fA)yp��հ����y���Qll׊��W;���XJ�j��X�QWMS���82��65
�}}v2d2q�~͚��$�ͩ�SO}�a4�9���\�1���G
��z���a	��_�Z��qO D�0�Hm뻄�����YP}����S)��/�� �
Vy�%HF���TCa�TH�|ݲ߈��)��	�B�
!(ǡ$�'x%F�r�]��*Z�_�َJ"<�:3&�9؎�x I��cܧ�q��?XRv<�衋���Q{Px���=�^������ٝŭ��^�D��p��#�Q*��?��Ǳ�É`=:�q��캱����(���������fwL�!��"�H�n��;�N��H��f���2*��H6�S����AeĚp@�O'��v��`�A��֭����Rc�<l�3�N���.k�g2���D�F�H�XS�,f%FA��˅��{��i��|̅��-����q��4.��)"n����o�9J��ѝȫ�C{��b�ahDsGˉ����.�^�!�7^�,j�2'���N�k��>�"Ŋ��Q� ��d�t��������5��y�x�i�8Bه���>v�2H�*�f�� s��\� ��<�V��:te��8�"�ƃ-�izzV|�ɶ�.0c;�<q�+�~js�t��i>E*�Z������	l���8*�؇�sWh̒ila�H�5S�N�w�H��A9=f�h��5#���#��jhX���&%i)��7½oM�/<��;<�>o����N�k��#�-�'�jN���J[R�A�T�2]_�]S�#���;>2�ӫ靨�<�C��e�rĉ��A"G|�3�/���N8+�KvѠaLK{0{��;,��,3n�g�|X�T���F�h����,E6#��j^���	���d7K^r��X�#wv��Jy������XL����!.��i���X n�X�{�u!3����2�yj�R��9Tߦ�����{�P���C;篟���ҹ�u��ʹ���s����GN,-At�I�mt2ӧ�~�ٛ�k�FFo��K�z�Β8���4�~���Kt��+�H"��-��ߌ0�5XD<��(�e|髰��l���O�PjfD�u�9��[��x����¢�,Er��T߾c�(myP<��s���7�z���`H?����t� ��\����9!O�K���M���cN�	q� h���~P����J�ૹ]k9[2�#W]N�!��O%9��iq�)�M
�4/��!�y��u/-c>Գ���hOb��S�ñ�Q�z?���N<c~4��p���z�o���F�:S}���u��=9zq'��}5;���0�����I�ۤO/���R���v�#�y�z�R�� vA���q��m�͔w<�'�v��.Z���ĔU�d��ǀg�q��P �2�~���LS1�x��Y�'m�k;l�R0�	��^T�I*s�����.��)��k�?,w1��,o~Ɂլ��"����CɆ�Kp䝜�"O>JŽ3�v6�������"h�@x�5�QX1�w�O��Ѵ�+���)&��է��/?
��錚���pG�K��U-�V4�z�Ј��U�.`�쩽��"-ի�Sx�k̔U�}���,�;Y� R���k#��q��ou@��?��uY�Zb�C��H�FM��[�P�1��=w�8�Z5`n�l�T���N��f����F�c����,��ü�{���o�e���'���S�L:��qc��E���yk�X����Bs�r��[S T�鏞�(�:��3R;�W�Z�Qs=0���rG�D��O�ԙ0���2�5�������S��v�-���.�z+�:d�L>K8��:��A���M�ٻ��4�x|������iS�
 o�'����df�5ْ�8�)���O��$��@@�Iuc��SuB�n�\�ƅ+�8�O�A���UW��ͧͳ%ľT+F�K��S�d��S����f��N�H~�g/Vkh����&�/h����z��P����(���0�>pzҁM�2�aRq�&��t^�z���nhj4<ΑpP ��ʦJN��Z��h��p����85��)^/��4�VR"-�.po0Iq��,��S9$�
Vk��F?��7�����j����qT>LT���@}�������.U��<����������`���O� r"�"�	v�r��'@����R��T[�/9�UKRȠ�-%�0��{�[��a�td_a8D�C&��Oig����qzD�y�SnDC�ї�+򝺵6��W�2�{�YG']��7��<��<1|>�5{��q�!��qS��Lwxu}Q�ש*` �n�G��4\�]�CEm��S.lǈ������ξ{yKͯ#>H]�Vz��^\���-�Jb��ŧO�!.1��v*�7�������n��6�+P4��;��)S@.�<8ن� BU'�&���^�� �H\��t�N�բ��HG�Ƃ�8p�Qh}S�d�,�[���.�� ���g9ŕ���t'�O�/�m�\J�m���{4r��&#���(^�5#o"��xE�H�&W���1���}�������fDC�
Ibq���N�����1��n{�ϔɆ]���fb_R�J�rUz��VҪ�j����&�hBK������Hl
�A�x��$�#�[�R8�+0f��>]�t��8 ���Nt���"8v(x������]/�QH�W�Z�߃y�:��TUc��(��$!���e��"�  �����co� ����H�����[�v���9u��[���f��Zن:%�m���₎I9�f�r�ƒ�6���<o�e�YXBݼ�����X1|ԥߕǐ6*��$]��v,���5�İ���وM�z���c�Zi�ZτtI� ������������~7����T�SN�}誗IP��R��
���"T@����3nV@�G�;�<f����is�ٱ�6x�[P="P�iҞi}&=Cs�*�q�l���e�S����)�≬�2I4��/M�s	
3��C���%Z���i�Ǿ�O�����A��+ �&��F~�j{D����G�3&�-��s�� D���[�B���[[�j@��������O�7_�-K�8wY�;��-��#�!�GO���B�=5zr���/���8���o���\� ��2���%Ԓğ۾x����鋦��-Ԣ�f3���[7��"��<T��z��.�>����`6�1�j�ף�0>c񅮚5V�& *�?��!�w%��M]�z�q�\�Q6��"��PR+����#�M�*�Ɯ_���n1�����µ������o��>�H�� ��	M
w����T1^�+sSm-�hl]x��#�s��o3�C�;=��l���I�"q�8�P��?x����yX�"<6ܷ�����K�(AI���T_}Gv�N��l�,Ь�JS����截2�ʢ)~V��z3�.5�(J6��=P��"���Z#������P��!��� �J������[�Ǚ�n.�-f�<��]]�bu"vqM}�Bi�
�GV'V*�:Wz�(�����.�B��g��GT����=��ʺ�s)�C8�3D䟵�����|.j����9��D���0�`Ώ�;v ]�B���þ D�7�^�_}.�0����:)�[g��X�3K�5D���>��hB�πSl(��F�����G��� ��3j�����Φ3��|�!�J���ɕ���3��y:��'3U�\n�p�CI�f�Fhu��[�֯(Y�8�c	^�(���4G�n���I���pa��)��R���^*y�ri��Dzc��ոe;��mH_�/��6�`�m7O����7��+J���+�I?�%�Ԇ�"�i�}ʙ5!B"�R�����.�i��P
豽������Ž�x��U>�*����NT�j�U�_�d$rj2�YPh0�V�St=$��d-�ͨ�y�l�KR�?}�˜Z�*�##�o�q��tQ;��"J�⾈�K�k�Թ�#�!'V�ڹ�������t��mB3�6��U��:�;8��D"��8-��M��Ihg3C>��O\��,�eɿ�U(���{��}�GШ],�<�PB_���a7�!4+��j���G�>VƼ(��Us��I����`aSٞ8+��=h]O���r��[��W�m��	B���H��~�^��0��D�~��=Ј�ȼ@=��px��Te�;�LsҰ��ݖ	��ݕ���S}���@� [�!V�q)�man�|tC����jfx��ӹ1]�~7��1?j���)�b�s��L�3;ڍ^�]��-��S��c����⷟Ţ,�ml!z��X�0
W� ���Xp�i]����f��Tsm�|Ӏ0M�I>M��Ś�H�
eL:��dy�k~��#Vo�\=+�T5�[T�F��y�Jvwn"Sr�\@)z�%�ҡ�"H��t=�R/a��{�փ��$�����L֠޼h�=~��V.iI{�8	�|�+��;_�hc�[��,װ�� �{F@�f��ZQE�K������QMqy=APs�Mܘ;?� �6Ɏ���x���S���$	r���j[L	s�fIȄ��t�H:|l�� �@��T%�/�+�4�n���)�JB�>���Y���R�yls(3dU-$�m���]�O� I�|'k�Wr�b���z ��`c��f(��M/V���)��ga�۽m��8�4�g�=�|�����{]��g����ы���6�G/aAV��C�\��g��\��X7S�>Jf����S8�k�*�_7-�LF̫��"���s
����G��G�Y�4Y�~�#{Cm9�cƖy��eq��k��L�����Y-��#Af����
��#\94`7�^���*���>��'�^8����IxZ���y��gktt�f7�z"�>ԓ�u8���)I�#��A��IW[�ؙ$tw�����d5��H�U;�W�H�>�펏tI��l#:��Uo붸�!8���	��]�]����.��H���T�%����%B� ����>��]�F%V�[�e�c�]LթϿ����cl*V0I�u��'t@[ͤ��L������{{6I�҄���jd����k�Ȑ'�,��8:7��6�U>O�a�Nn��bJ���m��E`D��O"	"d�v�|��D�?��Y�F��*AJ�-������)��>ŧ�o�����񫓂���ҭZ�@�Jc�=}�L�c���Ǻ�G{by؇�/�/�$���I����x��;���hap�B�����oA9f��M�Q������p��Z3�T��%�!�$b�������~݃��7s�!�jO�Jzu��e������Y����Is�7��At�[MZ�ۙ�%�%D�3�W�W	�H�x�u�Q��0=�x�j��+�gtb)�
�Ya�[���S��0���G:�=e@d�A����03A{G1��/j�5d��/�}f��G��ôEN��괞�aT��dHk�K��?�w�.����)�AS��ݣ$ʈ������YMx�	Z����s���kZ��1��,�SS�Y�GA���{ISM�󾘷�nܠ��%6>�I1'�w6�V��R� i��ɑf,ʚ��C$x�6��фF^�
��B���A�� �@�TL�����a�D&�S�;����qV�pt 8�2k!�rO�b���B�J���f�������*&T���V0P���w���i����T��Y0PmK�)a�"e�E~y�I:�q�c�䠬t���<z��iK)T{���E,/=��Ň��(fr18��E��4s���+)4co��u��aLί����iV��]i �B&�������z�O�
z:�無E	v�_?���?�"�������� ,)��"�)#��A��Y��Np�slo�	�-�*/�Aq�j�U��w��f"w�eb��n�,����F�����sZ��/�ҿ�	�Y�m��d�����4$c��>����D�t7Ζ��yY�aA���cȂի�x��z�P�;����a�t�Fy_�+�muX�`U_��#����Ocq��Z"C��d�Z����è����[�ܡ�G�ɍ�d�g��*}���!�`I��Bj_�^HC�3�7H�D���M��PC���]^ޞ�g��'���8��_��(r��.���vb�+�J��h-O�E9�����sW+N@�W�N�ƅ����tF=��	���o3$�a�>�%�#ez�Ԕ�6�P=L�S��[�!�l�?c�H0���_��+�=U�A�Q���f�^.b7�J{�q���|:�"����A^w'h��Hs_��+W7"�ky�S�\$io[2�WC�� ݔg��k����E)����e������g{���в���@�ֳ�dX��0[fj�K�)�E�
V���Т��'�x��]��{��#\�q�>����Xv�?�GG�(��lT�ivR
�&�@h k�m�u�����gR.dU��<=_%����������U��:J=1�o�t|4�!�QIU�����@ڹ��k�����@t������:F��ȹ��c��O�BÍ%l� �&��y���:	����òl#ބEP5GH�
��� �IȖ���,d��.9.�ϣ���(4�l��F<̻���i��q�&�HWg%2���V�Xj{�(�k��o�Yk��5Q�/%�*$J�� �"�zkb9�:���'i��؎�W"d�d��/��Mg�1U ΍,bT-��|����Z�� ާ��@����lcIvȁ �a��}���/ix?ظ_i�<a�W�]	�ʮ)w�h#��eQʠ�.^�D7��D�w��p6�o�ģULM����(�m��o�A/=�5@{DO&7MKm��
}A�Z.��!ǻG�|�h�V����3�N��{ah.�����s�)�wf�T�S����:*����b���ÏސVs�쩬U�%Z��������`M7_��&�3㝩X,N��Sׯ�"\�>�F�iFk�u�V���hI<]wRz;Ƴ���
_<�
d�O]����?���`-~.�b��$�0�c�����S�#���=�sډ4�է`�	^7o��#��gA�Vq���h؅0�x�&Z4gc��F�A/�S����*z�~�P4�
�{��=2!��s�I����Rߘ�}����v�L������X.|<% ��;�F��M��W{A�"2N Mwď��CS��[sOK��*>��T,����屮e��Z���-��$��K�%�R'������d9�J�u�+�(�(�������6����y쮊ob��Q(]<��nI$�AT�vB�3��i�p������*^���ā�I������y�ʻD�b�ϗ*=%��׵>;]�Sj���o㙪h�.�<�U�c�"|W ���ԬX;�Y�os��܇���)dOԶ(	��U8|k��m�6��|�i�%ړ5=�	%��(�'�._����&O��n#��!��8�8dak�7�m�!���n*Y��C��a����v�����w��w��y�;Lȝ5A"�slL\�԰-g��Uq'�X=`"T�MG�e^n�>Z)�'���a����TO�]�d��"��UCLG���̟���c\��jLQ��G�vL� ��<$��W�����\D����6�򞒯����j"�i���1��r�!���<9"2����Z�)����>W5�b]���� d��4�^�4�W c:e�{�iZ�י�������V��δ�ћ��3�W'5O��,��=�¹t%����Wt@z�9���u���͢(��+���5Bb��Oާ�挞ߩ!�a�L����;Z�ORK���_Oh�̂-�D�߾��R����mB�����f�f��`��9��N�v�g~�4���R!G}O�7�x��{��K�t�S�yCr{,�� �(��!Gp�v�M�����l�DX�P��3�(a����$CN��d$���u��66:}}`G�7���/���8]R�(�.�O�mw�:ݹ=ffN�ijbY�S<!���~?����ę̩ͨlL�_T�kl����؞VR��j��'i�E�F؛�HgP5{��Ul�zY)�Q��HQ�����ߏ>�$n�nt�!?X+E��"'��f��00��p��M����w�O2aIc�<J�8��pS텥�
�첨�`�yu�
�0����{&�e��F�kH���|#��8-U}���A���woQ���˝��F������*U���S6\�z|Cɲ�Zv;��͔o�E���b�c�����r$�����. p�؀�}��K���U4�sV�����]Q�2������u�|qzp,l�̣���zJ�6�  ]����B��ct/��t����9��HL&�g����:�jέ�\03�</���؜ty���� ~9��jz~�{�"�O�4�D�c8H��"���&9���U���,�n��ȻghX9�-���y���4+xT@{gF?�����= ��SJ�)�r�bu�zvy҆[4��7d�r��h_@]�h�����`1�8ݸ^�gR�5:,L�g���pA��$q���i��|ק��uz�d����`�V
��󬢛��(��Jj���A��;jD���)�9��A��zQ�P����b���vW=������bfXC�43�.F�e�o~1֔�5���om���F#FI��C�o0VN�;�l��(��ހ s��ՙ#�a@@=n��v�Y�Y���x]=��.��qL�����S.�4��g��gR����[$J/�8 ➱�k�)�׶�/�Yu��+���<��)���7�C/8��TV=�dc��l���9�b(��U�"�,���-����˺r\h�5Xk���B����-�y1�"���_���i��L6)���0�o^�+Z�Sє3>�GzRD��4.��*�a�(��*�uϖ�t��t��AJ$�f�UD�OAX��5[)]�ͭ��~��u[���W<�]j�<�n��X�##	�#oo�ܜ*�{8�������33�K��$#|$��<Z�z�3T�,��V���������Te�hWz�H0N�k�sD�E���9�5�&�t�{\��4�Ĭ@�H�T���%�H�C��(w� :�mӊ���=�����+��\h%�i�L���x5����	ƮW�77��_�?u1CE��񆚨z���0>W�a���;�����-�q.��LH=)l&��Y��&�1�m����{ |��߳�Y/'P��Y��F�-�kM�2�l�kX�{/5�ɒDlΝ��C��c��:���g�����$�H�7���f�@�-�V����/7�MްI�����7���W_NU�~�iY�boy� �ˑLf|� � v���ť��}X|��y��<��'���w�Am{�#����F����"�~����iő��|��ɋ�_;�b�V2(7���$��Z�d���Nec��H�G��NC�Jdױ�T\*�ēsx��H���(򣾀�Z_g�u� }L���yR@�'��I:�ix��i%���(>��1/�S��~"vyn��*-ܯ.T@�9�S��0!�9{3��e��bP���{M�"���|�=7;�zt��B}rXD6��
0��z���`O���\_�T7g��o�n���N��	���� ��m���<NL\��$ͼ��h��2�a9���e�i��O�L�7�c�yp2����ɿ�C�]�U�o{�C�� ���|��h�W�חD��Iۆ�6�y��6*�'�\գ:gs0�z��Σ�||�SOd3/�O#���ő�zw?�Q!��4��H�i�E��=��'���\c�v����{���][}����od&˟��
����g>=�A{b�����ˉ���v��Jpz�ZNnv!5fb����׈���u���Q4�Sn�vI���Ja�?Q�.���Wd�^(����k�Ec�c	�R���Ca	DK�r��oI�:;~�jZ��-�8�w���efiC�W�R�><N���D��Sv�u����c����$�o$�2��wh��I��*>��mR�^�b���Jsh�ג��y�+:���W�b_�O������N��S�����_v��&w�/�!�:C�jv�k~ �*�V�9s����x���\�0��}M�rR�K�B�n���H��^�[^J�
�3�B"�Nӭ����:~9�)x����6�
ѹM��kY����l�]18Ywu�l�?�/A�r�_���72�k
`F(2ܙRDI�NQ1r��=L�@�O�+��7S�.g5߰>l�o��3��0�q5{����H�D�g����P��eH��ێ�K���YQ����<�^61���X<8���=`
Y|n"T����WC$r Qsf������G)����E��VG�	O'ӕ�Ij�-�g��,¥��rB�
a
=ԋ����j���n����; �V��0	L�pcQ�7��;zцb��F狋�x�?|F�:h���Ԟ���a}��FX���N����.'��>�r�=	�Cs���?��>iΎ�H$*�G�Iu18.�Ğl�\����;�^PAQ"-�*������ ��mH)�/oM�/��h�g����t������3�L;���
޷��"i��0T�Y���co��������8�<��W�5�{͡mV��iw��ױ�LK����H���*h^�~"5]|)�0�6%�+����5*=�H�B��kEs`;��i���k�4��u�}��ˊ���s�:�M)�I{u���W�w",Za�἗3��A�ɬ ���'�f��Z���]�����`�l�����c)������V�|�?��A cs�� �^[KZ'��� �9��5f\�	\x$�C>k�[��o3�GA"z\~�<�]�7{�}k��T��MBM����e_�
J�+v�o}�,&H�`7�3܃��;ˑ��e�R�S��3U/�gS�؝��H�5�t��P�ϙ8�D�d��}�_'rp�e�CShF���ez>H��	��x���VI��RK����.K�SH��BH�g\y:�et���_B�Ȝ\�L�f��ؽ�f,��\�;���;v	��F��(����*�O2m� ��@h�����)���*5�
��ԓsfZh�'Ɋ����#�!$�w������%dXϹg�SW=�F|�����;�Zw�RK�˰5����r���غ�Qy4ċ���f�ɳ��9U͍��]��ɎXc�k�^�+�)g�T��c��E�	K3������7�+Be��v4���O�ky�V�WkQ�ҳf+C�Po�:1_-������!����{} sJYJ���u9Jۊ��j�u�O&0�F/�*.�A?;n� w�jKQy�0��*����x� �>��8q0A�,u�=�Z��_M}��L!�'�f4��b�M��M�Y~��0��x�@Q|�c�=뛀\��;R����4�k@i�e�4���`�Q]^��JW.g"V������Jrуt[5(�G�P3n�;�-җ�wk����9)H@Sn�x]tČ4AeYe��T4L�H��f�<����7~��>�E�'顳v�e��o{𱽾��)>M��+Q.��wB�)1ͳ�R���^ho��ޔS�I9W�X��D+W��4];gN��Z!T�,[�xP(����L����ڑxCOa�ɧ���'ޚ���9�kŢ��\7t"Cw�1��H��ջQP��-���+����z�G��N%�ì>=}2�kȼ�2�8k��V�at�=��E㊙���,�����6~���Շ��3�vj�H�A'��"k�Z|l�����P���������$���:����X]�W3pm~�i-��%��kU&\�W�P�!�i����h�@�]�3�1L��$�j�N�!VEW.{�($t!"<��y���oU,�ʑffKr�d��tE��R�]�n����u�%�!8�B_
T��+��~&�*d%m��=�t-/��<ט[*�܉g����j����ֿ��D���c�%˿z�
#�s5z#!�v `=�A���<g��"!ڳs<X�kw��V����݅��0�מ�9)�hwQZ�e�x�}����"����~�]�/U�Ps����s <[�db�#,*�+�-����+Vă��%}�|�����d��Da4�S!��U�q�W�aY6k6��D���x�F�}tj���jùI�T� 岚"����T� �Ꭵ���o������Q���6u����a�n�̒�j��;j�k�E����V'�I+�C?rZ�ȼ�pF0J��}�1�%m�;��#�&-��7�_Q�����ijrX��$�����&��ҷ�|�_)���x!K+���#i��G�F�YK��M��Bd��j}�����<���M��NJ�[e���-ϸ�E�L0��*�����2ڹf��T��/p�� ,�����~�J�&��sm������ W���P"�dӚ�3����c��R9T�JoAL%�Yu�VBo�&��<(&�u�Ӗ��'p���_�_^�	d2������?6��|�4>�=�T�!�d��z��p�Q28|�<�7�z'��D���[�X�1�RY��N�+�˱;DW� )�����\�ˤP��������JE�(V�:���φОi��K'ȬVS��ٻ$]�i���u*KA��)V�Q:�ÒOxø}��@i&���x������������찔=�+�_��Č�ݬ��Ǳ�ht@U'�
NB�Y8�A�1�N:(v� f����!�	�{ބd/<ӧ,���nM?�o���DdAڷ�f�'���n=h���ֶ�=i�C�Jx���/�����vD*�@E���!g�Y2H�M���ԇ�-/w�@�bud��(���ک��b�Oӯ#�6���Qk`�������	�����ܙ��5�������D���NF����˓�=�� 8�0�+�� Wn��/�nlA7��	U�7>��A���k�H����g��g��0������!9��.!��B|�9�뽜Iz���T��-�p��������
�e����6�����۟&�P\�hm��l��+�q�Z]b���%�H�NJ�ٿ$�L��t�m��v}ۦ��s~�dE��w��v+�wĂ�o���eƻ�A&�~�C���n��}X<26g���.��N>�M�F������/����08&��0-���W]+�&:u��VUf��<i���s���B,�m��:�)Ʌ�[��p��?�.:���p�ѓwg;�D�����fE�z��#bԔGW �O�����z�D-Tt��}��I�\�y�����\�����`���ȑ����/�2Ei�C|�+�A�����.��vY*��lW��#i�?�@�����=����#X�cɦ,+��(�`�U ;h���ʉצ�R���O(��V��`EM��]D���ISN��U4*a+XѠa<Ϋ^��0B���S�\��I+�VλH
��q�lk�^ґ��Z�~	�7��m^.K�v�y�B�D)lk��������9���-��@�|!v,i�S�*A�k�F �7�vF��84v�	����C��ڢ�3�N�_�ӳ'.��j;L�6�K�$��0��(�BԷӴ���r9��>(8b;��QsC������%Ώ�)5�×J�N'�e�$9]����S�ɷDw������CUM���?#���.qœ��.*�������}=Ý�E��y������W�aN����Y�h'�~��8M"�E��9�/�-O)`;s����0/� ތ�xc��=���b������
��&�b��Pvz̻)����Nu��##����8w�������x{�����;@d&Z5Ԝg������7[
��uI�<F۔�c�p?^�tA,�3c!R�
�3U<'�P�k8���X&�P`�	䗛@H�\������ I>�V�X�O\�L3�[��D�∓������>,u2�p�ي�I$�%[�+P�"U��^��.���Y�1m'�� �o5����)��"�'&��݋#X�-ӷ� �C�=�G�9����S�)�ĭ߷�"D� q���$�]�e���Av�.ih�U����x35AW����A�x�ec�bH+:*��Y�?���v� ﰅ�-K�3�6��Ž�1��J��$�����_�N���(D��A�.r;.'lf�a4�0����g\���z�g|?N7U{Y��C���Xcw���޽�k���<;���}�m2Bx_G���H55�8S�b$&ѯO���D����Onc%��f�.P���9�|��	
�P����*�]|W��h#�O��S ��O��=-��(Ez#�d0#_�'~�I�,?o��
��\^R~G��y�M��q�ީ�ۻ�]�&�:����b����f���-)��>� ͩ �[T�������F�@8�����c�"�\������G��чw�7A���~�)���px���b'4G�fA��]?�	L�`>�J�g�3����H��k�d=g�
��?���$G�sƃ���Qk��K�������I�c%�����^^A���-��ȡ0=�\�)2y�YӇ���m�0�;H��Kպ�k��^v"�R�9�3d�e��a��"?l�"\F����j�r�S�(����Q�J�m�����I����T]pK\]�G���Z�W�/h���t0�O@����o� ���HS����X��&���z/�'P�M���åT��6��-r�_IM�j�pGuA��x��)�t�������=���:+v��|a$Ϯ���4��f9yX#�x 
T�����c�z�<���isZX]�G���<�e$G��|U��X'�� }��;��;&���Фٸ�?�]��m����v�\9�:]�w���OL6FІ20�@q�I��~"1�4g.�Mm���ɤ�'I�'���2V-3�8��1���e��p�32����^�>(^�ѹ�[鿎iֻv=xTv���N�F:�5��L���;�fP�<���j	�D�d	�F���ά��Pi;Wn�AYF6(�c7�$�\)m+&�hl��B�'l�8ߚ��U���E�cM|A��f�a�`u:��=����ÐF"����.���Ϥo���s�;���Cw.R��^,)�l�7��[� 7���C��� .J{�G�ܤ4��{�&X"��Q8�w���.d/�c{�l|���)��l�6]��ه{��8n��*�qs��!��Ɉ�YCF��~F�b�'���M�+Qo]N�˩�V�<�զ�	��ڢ�2�~sd���M�-�Ǉ�4FZѮZ�4�����|����͂J�j���zGI;Y ��#���N ��*�%�Z��m@cw�-�;���t���?|7hJ���M,�
�Y�,�_;q���1�^3��4��	�0��+w�|��#_�,�e��B+_-��~k�W˄sL6���$RзԳ�����OF��Y(O���Q[h�CX�&�,���)�E+3��e�oVH��CB�80'�Z�R*�����_N.��6]�.�2��(�5�S�PW'�I@NM���O�`�)+��U����M�~�j7���Q�nq�J\�8e�ǿ����!6_:U�0�k��yP�Sh��O�X/��<Լ�d�cKc�O�2p��gj7��M�|\%�a��t}�[���n�_�����j,K�'�\��VAP]��J�vX�45孴s�5�O�W�od'�..s(�ZAQi�����}y��`�40#<i������Icby���S!+A�I0:��! :��A,��+pIgV�x^���o�<O�_���	]B�~d�cL�5�Qlc��]O��>  ����y�ł�G�,,(�X_���Mi��t�׎���Ĺ����=32��lv�#g��*�:X-[�.�/���VH���;��WZ�V�9�&�H�Õ���:��r�p�Ǫ�@�d0礈�=Н�tS��]��$\{��-��uFkͧ�p����߭�z�.T�j-1�կ�]WO��n?��{���W2ZAؕ�W��ɼR�z�1Rc�sV�4��<K�.�8��7sE�K�s��j��W&�����t�=K���g�D�~�����fe2\��_�x��J8���0	�FfK���Bv$=���0��qe����= "wc&K�e�֢��p�r�}Y/ z�h*G��H�Ω�=5eM4n%���'ϕ[�f{�o�Wi>c>d?6�ݳ�A��]fcRu�դd���heK.ϡ^�+44���|P����a`5��Ӓ��sl&�C���CW?<J�'�M�/ڎ�}2�G	��$�K��O�0L���zd?��j$�J��L����L������]�y��K��������*��a��33��1�2�����*�Q�5�f[׸�0[d�ǹ˚b��-��T����BD����� ��1�԰e�;4�D�bt�N�3�!�6�A��q38r����[�4z�W�����<��s_���M�觭���(��UM�%��O_#L��w�A��'Ϙ��$����⻔�q�~�ɑ��2�ń�?\�vJ�c��_������hx��D�]��S58JL�3��w�ׄmJ6$�L�&Da���h�p�� �(��S����x'}�Y�Y�'��5�@���ˢ��) e�jܷ����-�$��DPS�Q��F�F�R��̾�Z�V��KY��4v�D�br����o؅fN�r꣙��D\n$�%n�N���h�����L�!I`�=U/���Q�";�v��q�B�p�)�m��7]�ׁ#��G���������z�!U��+����r�Kw�[~����o۰�ɉ���œ8��������C�J�V@z��,��¡ЊU�Y�apͧa��3�M��=m�~�k��&��=4R��~��.��
 :�|8�a�$��mE�vXId����R��fP1�]�=g(k�kK�q��5v������n�J�����f�cgXU�!����V��QC�Է�ѳ�HM6'�0����!�) s�ʭ���=P������f�Yz�Z(�HYg��:�?)�5����]o���ܶ��ֶV��
f�s��xs�w��k?��O+K�k"�[_����H��z�l:z�f�X�45P1�Ϊ�ʑe�g����д�n�&d�t��u>�UV�Z�ܙp9�~au�*튄w�K3��G��B�������-�h�S���J�	\)������ڷ���t�.�JŇpq�<%�Y�Lļ��S��9��Y0�V!��\h�rP�'�Sf��?��4�@��w��K>���ؿ�m����^B3�0��d,K|�W�;�RU-0ŋ������n�2\��EAM����S(Ԝ��z_�
���!�?_�bR|�-�	��de�T���	H��4�V��$ZZ<I�ֱ��k�}���QG0�3T��?P�L�n��z;�x.9{ \C�zB�Bo�|�&]�@~���x�'͆ ��3�~P�w���TDf��Y��8P��ؙ[{�q�2+�CD�ϲ������(*�� 3������8hTl�Q��u�#�9�J�nVZ"��J��~[4H�r �c׈�
U��D,|ǜ�ﹱ}�.}&n�e�!�S�����>.fӓܓ��l���d���b8ǭ��)o���q�MӰ`�4��?��]О��|�}�\tEޡ^� h�)#�vv����V��|�w��� �m���p� C��=2j����,�&�%E�v���0&c>Ol�mu����c�5���)r���h�nkVĭ���I�@��6�vT;�Ot��,yˢ��\��E�]O
ϰ�ain#Q�n?�(bWe������ �U���qA U�"1�1nx
��E>�,�.e_[�ԁD_&l,�u���o�M+��V�5��R�C?~|h��pk�o�oV;��E� 8���̓Ƽ����ha��Q�Lq���`��<�-�PCփ2�T#�d��ٙ��8ʵ�������׏^�+�4S�5^��+-<Z4�<�!i��	3���D����5	_��bz#!��v�2�)��e.�����vB)pҐ�B�~T��<��*{����5�^̺Z&��m�C
C:�$��
��C�|>H\�k���dڧ�&`k�����Z�0x�~8V������cП� LN�{B6��ìd��C��^��ͦ�~x���c
t�9���� �^ݚ${��1F��s~q��79�O%�Y\uY�{R�8��\����~����n�iT>���_��I_O�3����=°�Ԋ�}|qj�[k�a5N5�hqt5\FV��V-�������mLt1��%�;�����` ��[Z�$��	�������!e�F̢2��i��Kx�f��aa�	1��@���:�vB�/ư����v	���߹�v\�%X �f�r���4D��c꤃3���`kW�s��%c��9�S�������aQzX'x��"#�|��V�Mx� ۿ��/�.٪4�<�����(M���f�ق���j$�q��^�7�*FG����m��	����w����{Y*�<����U�MC�sS��:�9͂)�Ra1Sm�mՕPcs"Q�]��|�K��1T"�(��G:��H�H6�hHz��)���%[4.�ö��f��|.�Iλk�z���/> ���J�-��?H,���8p��V��+�)��=�j~LN�3����r�x+�(i3�%{SaK�zY!A�����c8�'�q&�ȉy��U���}y����e�0��ғ`��/g0��H�V���D�+�	��U���]~�-,6K`�ց�+���L9���ƣ���09����:���-,�d��F �6ӳ�8!�},2�5N�b��(e�/����HI���<U�\�5�`��@�ݤZ���vR�W}��A3U�g"��R���������)h
|\b�~��A+H7��xN�����-Y�6@��B��)������El�zM2HA��=P�P����1:�w��:UJ97��&M�����>;V��cp���ë�1J�+VPI��r�s�|4��ᤕ�j��|롿�����e�� �#� �4CB扎V�X���BHI/����X3����(��_��'��7�<!��}����d��N�f��
�KjM>OX�~��E64�͖�B����kp�)$�_�Z���b�����Smc23���^e�_R�Bq���J�e�c�?� m��\l��]"��=��6U/������^�2&��8@�s���Xe���q���o��-�	S�J[�e׊�[���šp�/�^�rP t�5�F,�4�/��;��Fps&�[���A<n�_����%!����&u՝-��� 	�l�HE����J��!G�؅dm��L�Rq��$�(\㍳1��0��&����w>��\���;�=��N^ȳ�.$ Y�|�9j\���ϡ�
}"������-+\pB��o�Q��m�j��$����oiHJ줄�슣D���m�P�I�U��/c���O��Mɼ+��lC�G*� ���s�gu5K�*$�02���_žZ\��[3�Y��x�},/��ѕXW����׵���F3��5WQ���Զ��%��Yz���'�q��:"#�E�¯� ��ĝ
X�����3���t�:������mfi>�I")��1�l��B70�����#�1�pW)��Ue��w�k��.�u��?Ő'�i .Aۨ��`�D�2V�}�#���l��>g�)K��+���d.�Z��J�z�P�b7�P��W�2]x���=���a����3�|?�[��/��78�%�>�FƠ�mTNd�Y��g�T@�K&�dv�-��e�
;��&�'*V۪8���E���Y�L	������i��:n�R:�Z�}��Z�|!�>^h����eI
C�U1��h���!|�Z��#��J8?�ŭ��tX3r�0c�2%��Åc?����6��`9
 �z��S;�D)痿''�S�<�AZ�%�β���zA:����<_c�C>���1�4�i%5ߙ&?�ıQ�2����e��)���tc��(?r��/�l?'q={���3T���&%)�8zI�kk�b�������BJ�Q���t��Z�,x�$�c^)A˙��Ȑ�����ɨ��d?F�GqG����d�������܅i4Q�|o����E��[��M$7�D%���ܢ:
R�OT`�n�ԶU5?q<���l5^�.4xI����5�-�q��~B����]�m��$.�����ڞ0�*��\T2��:��-�'J6@����#���c����'	�t� �J�������v�<�)���TJ��|��R;?�J֌��;�_�RqJL������,�P�f�g�8�*���n//�Ж9������e�m>�tS��ԩc�M��0��7��{��jX1>�ܸ��~�3Bbf��������"s��Sc#���Gԣ��HAGB���S�#��7�����C.�QC�͎z9>�������c탦v&��=����R擔T䬧d ����4BO��/m��6捪��kNk\�C�*���ܱ��s|��Pl�qV�e_KV���H��������7Y4b�폱��X�b��8v���V�|������Exe��,t�2D3�����&���ܐp~�hI���<�*�䂘�����"� ���#��D!��G�V�w�h;�g�����{�A�/T�T��6�A��BA�v�jn���n�$�n՜f@ʴ#�`_1����X�<����� �]���)��y�Qςo̻Ѿ�m�*^����|dm�5���Ӈ����2W�n5oYX��G �V#w�L��g��ˎR[��_�h.?�՝�zAT�S�
��z����l�y���mb�Kh�3����[�^	ܬ/���#����oAl��S��Ū���6V�=��*űO�I�W�c�H�4��u��<#���Q݆2兤j��!��;/Ƀ���:��>	�7T����I���}v�J2B�kQ��^�jօ{�DYc{��dV�6�}���Ϣ�'�sa,ܶ�����lA��-����;�u3A�*UX(�ذ*��߿���)��N�з`��=R�%%u��B'=�ė�#��a���1��8��k>��X6Jo��iN�|TC�ޠt���S�/Z��B�i�^C�(W��M��<��=f��bF�,ۅ�߬�0>��_���A
!!
�9���q�ɋ��O���;ϭW.ú?'�6e�RϼlƁ�᪙)w�*�3`��jQ�R��.
��l[h�MM\�)����ȧЄ�T>�;Z�do_� *%_`�q� B�ؠ(㪌\?|H�NfG�����.���(���tYe����/�=�F����-�,d'������8�"��D<΅�,:�G?��f�2}������O��X�X��.G��D�e[�$���߻N�����a;D6�Ne�~zナ�X������b����3�W���Nd7�N���#�qMm��g���ְ��&$����{�hq��Mh�a�n�ɰ����=��8�~��ԡ�2�Rz`
/X�&-��!�>_�7��B��Q�`�BX֘{��ʑH��ʶ��/fn-6�|�q�5�Н��ٳjZ;GF��;H�8�Z���hY%�K3�ik���4�X��@/7�\�B�/z��E�-Z�c���XGp@�S� �Wm�M���W3K��#�JK��sb:��v�_c�C?z�� #�R�g^�\�D��$�L\l1�+���ƺ��
��H�@��NDgʀ��p�"�<�5���õ���%y(�����S�Za#��wk�Y�#���4����w�����(��Æ .u�a<�Ȟ�t݀�s@�2G܀�x�z���T� 'B�bPtק-8J�L�|U:�%���|
0AcdP�ˉ��W��],�V�=Gל�.�"o�)�0��mm��l����;K]�d�N����R�62]F4�Jda+d���R%�"��z��].��������?���	f�,(H���Vf�����;�GlA!�:1��"sk
�����]��U���P����}�Z���}�1�o4)�S�OxL��Mŝ�]3���x�a
Kt5�fG�9��X9#�V;!�Q17��P��xhX���y��\6oó�a�"�L%����o����Y�T'��?������p��Z�Ț` ��*6��4��*��1Qd[�9�cj�}�Mp�H7:�_�������G��ņ���Oz������W�z�V�g-z������<Vt&�ZfuٹE��?���� �i��z�Y-��5t^w���sL�G9�(�t9��=Ӱ�mй�ř�h�ƾ��A����l�-�Dt:�;�^V�"!sػE=�C~��-0GY��ʂY���C���,5��/؏F�Xa�o�n��b��o��=" �X�o�}�;s�c�݃�&��#���fu��.+d?�P*FU���kɏ�Эs��z�^�`��D�A"��m#0B�^�8��Hp?n8_�sm��	6��1y/~���o�����V���!{������ΟVN1ݺ�;�{��qm�b���*��n���I}���$W��X15'�.DZF���2)-LN��֤���\��� #o����4��W7Rf�
e�8M�ɵ4��2�lk�a�AXȺ��'?�lҹ�,��Z��Ū����4߰�5� }�@켐Mp+��U�wE�>��4�
�`N%�k[��M�'�i��_�5庛>O/+{�'���t��/D(RA�����<��B���d�T��c��\N!�E
�Xp�n�C<Xՙ�{�0��o�b0b�d1Zj���n��C�m��A8����{XzWů�~9��@��c"$
H���| ��I��}��6�9X{n`|6�Q��9���n�����i���ᶚe��̼�R��e�-��R��i�)/a+�i���7�j��Ԅ�s��C�k�
�^E�̀�Ӏ(��vu�+�eD}�J�� �mK%FR�o2�2�;a���w�Ϝ5"�\7�V�gG%f�'�3�Lj&���LiKC�Gu�cE�~1�F
F�V��?���K��:%��nU��I��6�!����Z ����2�{HrZ��B��R�=J$�@�᣻U�YN������$��ާ-Ur^ �2�̮�uSO�?�.������˳lxM��J�M+�Lkg��$�q���F�S��r�"hBq�1(�*�wf�o�tut|);�Yu�����cj+k��Oh���86���CjFZ�A����$ć(���5g����PY�w�9�����aqd���o��_�[�����f����1�jIsYG�;��b��ki}AB�ϟ_�������>�a�V��gfا1�5����*��+ƿ�g�N��p��-oߦ���y � 6�l��k�0e��B��[W烚������)�d�(\�Y. �$�J��e���B�[FF�������4�r?ĭN��*�|��}c��GY�o;S�\�*�:���`HTs,����v|��RY��Y��bL��أ���E/c�W@�z'�(ה�i$��4�"�oj���j��;"��<�ol)��g������(�3�IQ��$�|��L����Ka��ʚ����h"
�b��۟�[$*]�wou���9C��`v��l%�Օ�VG������R��Li�� N��н ���*:������*�Ef��W�DB�U?*)�v�����wM�\Yg���*�I��G~5�ZoJ�,����|[�t*�D�&�I*�ci�A`�.��j�f[��<��tK���)���\o�2��֍U�a�!�5��l�YV�s���In��'����ۋ�0�����zw����"�D0}PJ�\V��_��o5��m8�H�g�~:2S�h�ng�/�f�<��?��ΜV�~�9	%e`G�������8_&`��F�{J ��K�s����ZXC�Y<�R�cm�]P�nPK�	zm=�^��t��!�T�c^��z����wq��-M�KM�����S�#�̜9�����%Ov� �`�׋��X��b��/�6��g"�O����nP**�t,��4}��Ш+|ڌ���+�Qr<��y8L��i���Zۍ'�Fň���@��Do�$���h����+��ٻ���t'دXl�P��Y��Rd������Q<X�2�_Lj�y$��SC7��PI��9�G=��d5�5�gC�k��s^"���l�Y�P�	M��f���g�k����aZ���;�),�?}!ȩ�ثu�3�ot����/��ـf� 2��׀L:'��Iڍw�vi/����q(���j�wC�zK��+�z� 姴�lCC��GayE�E��lb�9^)�5��o�_�a�r�B���h�>.�Ư�����@*�����VDͅ���3���`P{�:�!�P�2<����p���(�\��T��OW1ycqG*Ө�O�Neob:�F;��tƳ�P�x�FE�� f�)REz9�� �9�3��p4o�|�i�mm��6�J..�w�13D���ߤ�����X:�����S��X_��3l/
�d�p��}����-	�<˥Rց8�^uc��6=��qRg���,{i�ҫ��{Q���L�W�e���z�����:#kV(���( �e�ڊ\��\�Z*��ȥz0�9�[v���ƢQ�qN0��N�����@R��IE;�^��z�����x�+DS����#g�P�k�:�&RА��j�9����X|Ź�|�$����0����׮2X���{p��2����WͰ��}�(��)�gxdߤ��
^�d�+�����^:�/�Ț6��퓁a��S!�?�rnh�sNk�b���'D���~o������@ͷ���=z
JPLŖ�M!h�>,L(��Ǹ��}:�bዊ%��֏dh�����""� ��w�E�,�y�R�b�s�67db���b�E��Y���WF���6��8��g*��[	ِQ��u�a�:{�밴�U&�O���-�цTT�;��A_��1�2P�[#���[H4�7�%l򪫊����<ĉ ց�U�#;!|C���F#>�����Z v#�c��Z�_��y��?X~)��C46h��F�o�$����:Ä^R��l�y�4�\_ޅ/�8��ܣOw�������ԣq9��BX4���n�Ag_ʳ8��x;�*L��֋N��aX� ���<��;bM�����:oG���y�L`%6����J*�01IEQ��KmM^�8~�V��d�����o���h�ej��<�;�y6���0:�Z��_�q=&�]<��F��1է���)�s)�#��d�	����I��/ụ��k%2�2rW���_}=_�$����yrs���Le䱼^ݶ`�v��7�?͍�
���ˉ��9|XyV�x�ak��ֲ���],�-��(�)�C�T����D<ݺ��ycJ�Lم#g��'+U�m��>����/� �`�~^(!~�)w�2�5�� r��Ơ�}�����]<��c�J�9T�}���x��^w�D؂����xݗ�� p¾���$L����5�䠾�ƥI�߫���0����f@g����� �|��p��(�C�K�K9��l����������+���@�|���	[���b�A/q���ObG��K�%�c|�E���_�f%a�~��#t\���eŤZ�N�-M��������	Ω2�!Yjk�|�=�*�!:X���X3�\w9b�@XT�%J'Ȋ;���씘W�������6?'��DF
}��u�	�����6�j
��� �ע�8(.���*��M�� V�}� �=�6Ie����Z�kp�.󥇗N������\��Y-��j�"���:B0�Cݾ.0Y�t���W#~/ɷHx�ވ	��kz	=y�B��}�x=h�2T���b�����#T
&@{�Sʶtޞ���D�X���$H_��������G�,�y��2��Ն�r>�&:I(_�8�Qr�� ��3����֔%�}�X��_�U�(�bn�$�`��_�Ay(���jY���Q�2�,��lI.�{&� �RHs}��T�&$�r�dΪ��_4�H����u9&:���ϯZ�cU�bO�)��C�hң9�����	����nѦ�^_pnЯ�#���=���|�%H�bѵG�d��E�)�l�Ԕ=���%��̚�:��7o.e}��\k<!t����:�(��̀2b_Z�
�_��R��EO�PDr��\�;4E��޾�⷇s5���Ϻڌ�>۶S=�?H$�X�z�2e[���g#SD���v�3����Y�iS��ER�,�}-T���?�$_�!���"_��
�A����������JOfJ�ٜt��&�Ë����(����`q�]Zb���Z��N������� #�v*�3�;�����+��,BTk,�H-��l�)����� �#aS�\��㿅�h�Q��H��}�E�i�[ф`�Q��6O��W=���&1�	�R��v��Z�\�������_;
��6V
��=�azN���c3$��t��x�)��hw�\�spv��Ρ���4�KM�ɼ^ߗp@��8\8Rn�g[�����m(H L `��­K � {�76�S��4jh�����J��-B��mm�JC���T�Vn���K H�5R@ρ]��f��avO�hT���m1�M�X{}sU{*����n�ۨ��>�ȟ4�;���}+�J���������S��}6�i�u�O�!sg"M]C��D�����q���ȩ�5�{M�Tq0����O7T����.����p���zI|��%�|'��s��
>(��9?�r lŨvŜ�d�\�㙄�(�I���L*^�9hE��� ໇�L������3��H�8���[>���O��)x��c�{���ӻ�
�����Ƹ15`�v�0@��
��\�u��x�1����i���Q|O��K�ҥ尵����DD&�A�2���v�S��g;�y��y*ܿ���z��2��@XF�v9����i���&��Y,�?�Kl@��v�;4�QhY���Z�wk(�p72w�����I��lSi�������:���W�f'H"���Z�����I�V��}���R�F�a��Y��C��u�f.a����]f���6��@N� `��piX1^��@����F4���f��`���ܼ��+�`�rxwPWCԞ��1@�@�M�m���*D�a����zT_�z&��p��m�ޢ*+�p�Q�\��D�RBK��'�
�0@¤�P�����څ8)�y72yb��-��˟��i�o�y�A��q���\mN9D~o�k��yT�j�Y�ϸ,�ƪS��N���Qk]�*�#VBу���8��T�q�#�f�����Q�mP�/�m[�gi>6�uh��VhY�S�un}_4z�d	���Wg%�Z��=�AC�㭚�4���ed��G������LJ�欂Pg�6G��*z�7-�٣��{�N��;�E
�l��Y��!���~�_cI$6<߬�2���?�o�R����V3UH�"��=�ӵ�Vo���R�dջs�����)Y}|��@X�Pq�3�.|��2�1K�	4��Kb#�/�i	cC���K�s¯���k"B��ڡٓX���5�x� �9{�#ߴ,l���:n�����N��w����9�m_���iS?A��O�!4r�>u��������S/�y%<R�W��!m�W0#�8��q]��8ⵁ�D)��QT%V��~7��B?�`g����$(n�v�:mIUk�8i?/��닄�!��������bl���߰Rky��h����BJ&�<$c6��0�a4������㭦�B�%]Z;9�I�g��\$}K�����]�.��x�E j[��ߊx���F�^���Y��ǋV�(JU����H�wm�F�1:P�H���b^�=߹m`5a[zHȡ����0R��rOGDk�V�q�����`�̕�N�t�>U��0���;�y�U;�"�uiw첨�i�n,>��Y>:H���OBV����ޟ`�k!�*	L�V���P"��M��q���b�y�6+_��Km����H���Y�N��i�f��)o��4*n�,�-�mEĥU4K|�w?XW���'F)(����0lW�~A�t*�@��k�^�	�F2�YWy�|#=X_Z�U���JFuM�@�o����ãJ6*���%*D�:�pX���������o�E�e��bO����[?q��Lc��';����Y� �J[}m4!j��"��V��z�K G�G�I�|`�gE��Ӛ�Z��2���
�Lr�k2�B:��b��M@�U�f�$�	� ����o��	Tߩ�é��kؖ��U��o�*�A�6�=���R��������/5ݓ�����Ϟ�&/�m'�8���+�?R����ɇwN�
^�~N����y�-a=d���B�F�|j{qQtH'�y�ۈ̧� /���'�Ÿ�@����`�I\�1�YX@�
��mI�U�^a&m5�M/`-�-suT��X4T�)��X� sVZy���m���/g�ebXx�tlq�5����vxb��?�7��PB�~�=�8��B�"�=L/F+�6^h<iUz�Zĕ�&P��Rv�M��gW��fu4W�?��?�5��*����)�=",-M��v�P�7�D#�US|��u),���϶&cM���f>HÀ�ɴ�|jRD�Q�R�u��
OW`}�=H�f��p֙"�Y�a�,9{�Y�8�D��0L�]�dQ�EI:D$�S}�A'N�7��mY)��1�؇�@�쭦�r�I�:�����j�+���'~��<#'ܺ��P�����Oc�������H okE�����7H�1]����l}�G�uT��S�Q)�<(���~��F����{J��5�n���&�8L^갅�5���d�(�������rW�(���,�st^���W"6���hM#��Ly�C_�����[1<[t�-6����J	��w�֌��g�'�;���I�w�c� �✑˿ a+ �����<��-�λ�_KA	<^���p�� ���9-���ܩM`�T��3����BC΄��p�������a�4���7	�,�V]�>�m���Vm
����_�,#s� �˼e�$r�)#q	.۶���^�Y�`���B$���C�N�z,�=��v��I�u�HT�]��D��>w�lRO�'߽A���x{� L����4�WϖJ|�H�e��SM3O���2q�O�Q.��xr
ͱ%`��7�W���jj��ږ 3���b�.˲4��kۤ�	c��E/��<�_�qC��擊 ��4ҫ*8}=�J��JN>�=�r�RD�f/r��h}iM_Ӌg�(y�HA���K��)�"���w 9�{K��L�ʐX0/�_A6�yBÃ�̫��}�bt�2p�V%���od���� jb<,��rY���9kq�F�,+��I�Y������ {Ki����0:�"Zh��r�>��l�'�_3��p��4���=��<u��#��"�BZDϽ�w/����C��)��8�\��\*�h�H+�@ ��ͬ�P1d;�cӮ��tH�͒�DM��cc	��_�l$P���'�Q�����`��҉6�
p��5��R���4%��-��"ҲT4Pe\-
i��y��rr��B�[�`˱ ����'��^�5؎�^��+b#�gL����)
��>����|'�Rą�A�h��;s�`�*x7���ׄ�s�
�L��(�IpsȬ5�!5F[�B���-��Lz	&U6����O?�c�V)���	�T�b:?%S,F���xdn�ݲ��ƫ�^S�������wv�6�Xu��� �I�aD9x��O����h�j��ٶ."}"X�ӽN��s�OJ�3��6ԖQ��|4$RWϺ� ]OE�s�^�p����ϳ��b�g��g+v"�H���6vm�8��m����K3J�v�kϰhԩ��/�ܿ�)
����Hj���|\q�S��9-�k�ױQ=kX7��"z���Ad+��|�K�0K�N�u�J��O{$�t))�Cc��v�CX�[�#�����@<S�⒉F�A9�A������