��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��U��ee>Lی�I��"�Sy�#!���Vʘ$QL�OԈ��7c�ð]�}$N��t��zA��R����-���hO�
��{�T��*7G����.��E�t��|�|Q+��;i��a!s 0�Z)f�AE�T�4`*�OvT�&�4�����1��	�'o(��4�Y��Y\�
�%{0qoW4�@ �Dع��,�4�1Cк29�2�|(������n����RD��+_gec2��jr�UAr��!Q.���|՚�f_h4���t�^��4©��R��֪;��GyI��6n���^<EѮ H���7��U���1��K$xH�^g��L��0��C��=��>'��%*���T�])��f�dfl�	?��U2�\�?���s���V��V���+H�%!9K>�h[O�>Jc��OXt�Pȣ&݄��n��4Wc
F�>\�-�l�S0�>�����Ff���/�#���'ǵ_N�(��>Φ�詳"��EJMP~v���ɵ�&��%:�u��7�ϟ��븿:W�W�����@=c��j�U5�ۦf�f��5�!��/�>�N�s�2�u�ȝl���Q�溅�7��*hf=1��1����@ ���I��4�C��e��QV��R��R����A�x��,�E�.�  P�D�	s�e�`U�/y����4}���_���HC�CIu����s�%�btؑ=��3`���:����-�,��aB���9r��<�F���BL�0$��:|�?L���O�c�*S�A5 ���lƑ�g�e�C�����Z���B5�f��h)̣��^��T��Ed�W�(�����K��p��-��f��''�&��u��fz�V <#�Z�:8��c#}���w��k3�����ɮ<�UN����y�O!Ss����)�'bȯ�������]�=��j����;��^w�-�'ظ����s��"" Ow!���}@�ِ"s�4�9I��S�x�6>{Թ�B+�a�D׷U��T��r�E+��5��?��(*��iwCڛ�Tj>,�r�l@g}�������>��5�yD9�?�f�$����:����=��Vh��FM�Z�*렪7O�H�|��MVrzo��PY�8(l4�Oܚ��� ����x������c���M7-�B��}i��xLd�p�����%@FYaZu���nJRq,�̚���3���g	��hX
��*/�8;|L���]�h4�|��p� �ܝ`*������`O�8�P{�T�oZ
��A $0$��cB�4lq3*��P9�kk@O���X�o�P���y/�E͐��v�>:�H��e��Ysv���7��
6��uC�o�[+;���5����.��%��#�	x�H�RH�	��v�c�}.��&�۸��Q��|:���:��f/�ހ��Z{����
8�(h��-�n�/\��wJ9�5o7å��D
.L�m�c�m7�1��>0qC� �f����������5{B��r'����?�tV�=b�����W�vG=Ȼ��Iz���5��8NDSq ����"Lt}v�A��������wU#��1,kݮ�Q5�D������>���KQcң` zEK��x㘰\�	��5�`�/�����W��kb%J�L*�N�1[ ���p͋�<��sr��p�΢��B�Fm$��J<�Y`*��������h�Z������3�R0e��0\�U�"Y幃� �B�HI��.�M�?����c{��X	l���d^���ز��S�M�M��5M�i�(��#1A9����<�b�{�R�+^�P�Tý7���:`^��Y���5�1d!���Gt��7��P"4�qw�n�^a�X0E�`��Y�ε�c��L���Gk���`B@> ^%2���A)��
m�"Y]"���8G���札��T"��?|Y�2e?;���)�q�m_�LPdP�}-�uq^�XRX.B��GI�L����F�u�sf%�׬��]���*I'��+\��:��!b'�(T�t(3��J/Q��<֦��&�U1��OXu�\�Wp����G�lE�w�5�h��¡S��?�����j������	����'�[Ch?�Y�9�{����5�x^�4���0� ʪ��T^%�$3@V���]=º�}��H�gܛUR&���A��>D=Qia�$�� X���ъ:m�T
����`�V��N<S*�B�R�P��O���@��n�ګ��s��g�>C�I�AZ�I�i$�� 삔�s���~�Л�96��#�ݙ��������#��1�JZ6�|�L���3�͡>zO�s�U��;zۀo�=W����y�"�`�%�hHFy	�z�a���x��hX�
C�?����F�jD�r]^�Kq?׶Q�-b��2XX7���n=j~��,��t�o-��*5XX���;��V��g��;�����G��Oӽ�{�Q8��Euy2�Y�Ǜ���sdR���Ѵ?�r�=��2�H&Щ��V`YMP#!o�
ŗ��1Ƕ�%^�u�����̕��cj�E�|O�~�cr�n���ݨ�'��WF�����ݑ��㈧0����o����[��B���
B�����J����Pv:��Sܡ����Ƣ�����Л�'.1��b�p*o�Kܷ�L��I���m�	!�t�̻@���oi򛧿`�{H"�cd�
i�S]|�~q����VZ�����K�$_�4B/J6Ҁ�_sS� E������# {B���c"~�)+Ֆ�Q�G�$����L����4�P��֯.W�G�*��_�6=k���������=��\w���Z������5z�U~%��H�j����Tt'����`.�u+Q�7�U��2�`-°h2Zϩ�VS�v�R�whC�c<FM�A�i��Ŗ*��d�>�gBi� ��s��g�#���&��P?Q D�Ϋ�����f�w�3�h��+�H�i�f�� �g7X��Њ����2�v�Ɗ�"ͧ���y��;~ZR�,�**�(�R"d!,��xL}Q*���?qv$�y��~6��m���:��#c����xF!�dN���E�����(7�3�aH\�$�kT�^�E�u�J���,ޙ�T8:PQ����A�D�Ǘ�޺�<��b��7�N�� 3M�Q{�k�@/�_�~�m���y�^���aCs�ͭ9"�L�N�dKɳ��g#��I��\K-n�<�Ad�В���N����N�@� 
h[�>�J+��T�Mi(�g����e����>"y5����\���4a�ӳ�O��U���uLQ>�5�吚{�������<��u}�j�вxY7z� ^=B��o����:T��a�n(F�A�^SJ�m��.p9��������K��7c�r;AF�E5���?a�	(?D�J��`#��b�ŵX� �2�f��)�':�j)���/�*�3�n��R m	g���x4�@nx���װs�8l���-�j�ө�c=؄������Ǘ'J�~�z&�j��.3h(j'�,5<
�&������#U�%'�����+��p ��a���6x��洖)�cG#��_�ݗ�Ս����?݆}7� .Z���k�D�}�<�>�
Xi#	���Q6d�G^,�yDdWv��!�&X1$_dA Hʮb���9jiRV܉�ơ���>��%�F�:���EC���)}���O���ޟr\62�V��L��z��9�`:���S `M=q�/�!�2��
C�uP���SZ��kǻ8書LW7��)^	|� *�=}֔��ҕpzL�Xී��}@Z�h		E���B�[�'-�'�[kLָ�8�5+!c��a�c��t;r%m�.B�H�Ć�O��G\zsc�2f�߉�3�+N@#(�N�յ��+��������&A�	��΄9J�D8ϔ�����1��'�����%Q�C2�O��?�	Bq���Mҥ��u�X��WQ�u!�r�T�\�M�J���ۢ�?6^����O�3n:r;��O}���B���+��RH���
��~�b�U��e���4W�e��I��g�Kv��n�I��7H��N��aK��P������bO.De��s�y�B;�����C�x�����"�F;��i�ԩV��8"^PP����"߶�8�2��(]@N�N�r���[�bA=�;y� )����P���&6O��5���s�����ߎ؍%p(�9��6�t���y��.�h�el+^W��|M]��p&��Щ��݌(�&���U�� �Z�H��-��%��t7��*�Yb-�~�D��X����G���fD$Ǭ��������7�n��p�~���y�oh���W��f��Bj>)y5�匌��*s�Bi�gv��1@%�Cdw���L���2HI�����>��� ��z�ፕ�P?Z����<NTwmDw`�2=N6��K&��I�k�T�C$Ż(��T{ӵ#.�|�E��*�nM�Q4��ukY*3���>�UN8�Y��A:E.�f��ǌ��V�Q�<��̃;�T�2i�ގ΋�t_�N���ã
U1���l*�r�k�|�e�e��6Cv_bx�.o9ڱ.��l�~/$��H�K��>�k�Ń��I�Nt)�&�k��+���Z�&R\��Ō(T�l��Hp��I˻$@Ց<ҋ������V,A;WB�#�0Ö�|���-3��	 �M���c28��h�eC(�[�|d�_�V��y
E�1UFA�B\�WP@����_6����ҝD�f��D�FyR�Q�������O�	})�4���e�'�碷��Z����N5$q\��3{��f��C�5���T�u�D>J%���̷ߚ�X���=��Mu��ۋ����ԕ�(��`]�t���R>��Q
 L����^Yl��u V����Ҵ���ȼ��;��q81��}���$	M�X���b���M��;���a����]o��\e���$�O���|3��H���	��F�˝�`�B��BD̨�-]s@r/�*�l�jlZ֨K�t)�k��
�[��#�O�h��C['O%^����3 B]��ۿTK@��ZQ�$�<͒L��"��V�@C�ְ��^�X����L�#�牝(���.'<C��RJ�6�s��e��*�
L��Cw�͌V������?C�=p���e���؈5+vd��fRA���n���~Yl��ww��?��°qL`�Ww���u-��cF�Ҡ����`�$�n���d@[���u�~|.E�?�9C��[3�#m�r��� ���:I�\quj���
�\\��5��,��d�dg�&��-��JcP���y9��Ǿ��*py��z��}�+y�T��!X�i\�?��מ@FS���-�GG�ZPv���"�W������G NQ��+� ˂b�
�|Ո9�g�z�J�Pk���&����eoV���W�ݸ4�)�~0��U��Q���� �l�[^���Z�_��S!%�W�M��W��[��e�ֆ� �$*��"�(�GOp&���'��3����_������"��vw�
�8�4����C�nFT�� T�T}ǡo^� 	�Hv�D�E<���[?��u������p�K���]�"����?t:iW= )���V�9��s�%jh7>]� ���S��RWz&�IM�@��������ꛪ�m�>���Ck���Ιx�	��~����y��cf�������I��S�S�'n��1�mz��j�:d�v��#����s'�u�xE�_��<�u���I�{�3��%RtՆIӃ�'�{��,���D�s*3u>R�>�yP�f8��cJ��N�|i���(7�vK}5H�����5�T�u�{!�:Q�zr=�@w��O