��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>�m��`K����;�U�����wh���Ո/G:b;�x�]B� �Uص�u°T�&m����Inx�F��|�uR{u4��GH�xh4��9�%�\x�c_v�O�h���i�p�����
�h�����J�L
��lA�Z|�~����1�=����}�k	��XV�Ŝz�4�)�y�3�a&~&���'�dlo�㖖q��D���e��I��������(�oK��+G;a)K��=c�[�$�~�'��u��E�d�wE��wFlN���e��-s���p����U8c3�aT��g�����;��P����H���L>ί��ڲ �+�67+ܴ�,�g4�z�<�!�.=��m��ǭ���'a��\����Sr�M�v65)~�+�{X��n�C�\PQΠ�\����G.vLr�ͮ�"��ɐ������2�1c�%@�-��I}7WN��q&PB�
uI�FX�}�1��g6�s\��8�G�Mm�}�F,�
�Gc�!�R��-�#�Fj�~�r�%���3/��Ry�� |R���!�f���� |\����P����0�dBW3��y�w�-�Xf;��D�5o�Fcs/�j�nŚY�s7/��ӷk�o4�p��Z[��Ha�j?���a�2�����}�@�'�q�g���
3�D��̺�g�~��\f �ߘ瀾���b�u$���b��v{ ͹�am���}x5Z������?}8�bU���,R��F�_�1
y�\z\���� ��@+-k�`�M�_��M�{!���n�[A�LjK��� Q��]����q�3Iz���'_���\��2E6�T$s�O.�%Beѵ��Y�Jv��;E1[��F��5֢�+W�)㥀�zXb��k�`p�q������?��#�[y� ���UB\��;�뉖vx���8+<��}6�^�S.�@����|u��R�E'ÑdW[Թ�֧ȼ��rfqmr�Zi}!7���ru�8ô��'B �E�(��X^�.��������|w2STKf�F,���c�L/5�ٌ�$����imƼ��ǈ��;�������:!м��)̰Ƃ���7"�,��]v�-�L9}�A����3��f�i�h����m��:����Fdu��>
5Q��HU;�cK����v�78��J�Y��c�F-�H�&���4�U�gj����Г����p�~�E�n泰��鍴������e�`	���f�\��ěBcU����1<�9����s\Պ�YV@q�Z��M��'�c����d�rX��/�}�NiF}Uj��ܭͬ3v�wv�&ͩN3��4���T�K��H�$3z��T�nvά��>�*�F��� ̈́���L.:���1a3����5��ʼ`^�]����	v����2qUg�(B�K�[R�qbl�x�,m$��]>D(�q�D����Ji����$"��a�����IAZ$��Z�[�4�Բv6���VX�s���'��]u�qI;J�B�LVl��d��r0�&�����Z�A�eb�O�Uֽ���j�0���{�X�f=��$ڠ�w��fw�u7[������w%�9���L�E򍬈?������n�toϣ�?$����:���W�Eh�K��U�8Ϝ�@~oD��e��YWA�n����t����z�FRD��[��T< Xg���kF0��g�l�
K|=�F�s9[~�޾Ϣr�6o*����	�G0ގ�F��̬�y��Ufs��z����+���_�
�ď�l��٢/9�j�AZ濯\�}�cٖ��}�ߚ�	?� Q�r��z���3����G{�H����h���m�D�1�榚���a���)j�T\1P$��S���
�@y�;�2��[���W�ԕW��+���������n��<�o�G�zَ�|SJ�#IWz�'Y��j��s�r�JT���'Ft__Q�NKb#_�a�>HW��b�_:V��s��?�XBٲ����1����i`��K_'��3���y�w�j۳��&�V��u��6�P�Ϙ�w/׹��\��J����kק�a�aK�d<lXRƊ�<�S52�S�B��P�����b<��$$���!���h�m6L5/��HZ����OXpIZY���)�4���~0��@�.��o���\�E�Ӥe��]tSFޢ�U��<hJ�n���B��� v�l����WvNrS �Ŏ�[<� �*hh�e��)��_I��k�؏�%�&p;(1�3x쌹�M(䶯�v]��=dsN&�h��}g@�{�t�q8��O�3�Z��%w��(�=y��Q}>��`�b7h���_�-i7b�HP3^���W9�5%a�Z��&�7��4�i�+v��O�#I�HF�7d�PIh���k|M9��iR�	]��}�����gQ��զ���M_�S����[�o!�`�igN6����H��`�L�3nL�dp�Y�{!�*%����V��z6��ϕL5ּ�r̥J��Щ��"���<g6�����I���^^	�����Q���!����-(L���!doZo b��\���������b�|Q��aԘ�s��A>n-�'˗���Z�6�%����0W���)����;�@R�5Y��<I\k�=oZ_H�[Jmh8��F�2�h-,�)��Š���)�R����D��	����ϻ�|۽�P��;�$��� ͆�dUvVT�x$̗�ܯ�bI�ȡ���:f�		,F�gN��i�e�	&��e�ioH���*a�T�a=��vi:f�0��>�ʩ%��$���uf�p�I�:��t��#�S�i��jf��V����e������Rg�
������ij�K��!h�4q`K��~D�J>5�3;,Ux�e�;tę�).���8�D�A���_�9��k铈#�k��U���c�"�V�8��7��V�܂��"Q�Nf�='d�T4Ƣ�?2i`��J�����kwP����x�a�|;��yU��v$�(~@�x��9��϶���;��R��{��1��Х�n3�����=���4��J?�؈�\���.�Y&�W�2e���)��^�w$h�@|��	��c����@�w�w⁛v��q��⹠/�e|�*��g�Piü��\ل<�b�Os""��E�.R��bL���sTd��xK��圕q#��)TԞDG���^ �P~�/�Ԥ�v�ұg��v�!
����UT���PGպ��>o���� W�����Fy������a�,����S�W>�`Z��`�>����?p9�����k���5��+�JJ�nF)����'4ŔfA���S���Z/1|Hj���-��?`�㩑