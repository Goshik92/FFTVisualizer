��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�6��y��Q$�Q-�
���耑�J����Q9*�@TU��H�0������YՖ��3�~ʙ��\�Z`�Da@a���0�T�ު�?4�����9�W�88-��N}.2cu�37�l�*�u��aR#@�/1?�F�w���"R�t���w�A�bW�E|������}����l���)i�魒Yk�[�м$�*��sfj�őp��{��J�"����#]����CU0[�����D<�0���G�1�����4�H�o���enH1��~��c�7ٛ-���������,EKxo��(�b������X�ko�B�jHVی��m؀� ldg���U�z6C�E�M����*����mrg���09�O|�=��L�w2A|�u$CG�	��ὰڬ��>ZG�8��A�&`�dq���v<ҡj
Rd�g<Sl����9!Z���m��S�A�-�
��E;۴u�mڵ�D�����#�`�o��\����5�	<&���}'t}���o��3����\:���~����oV<~����>WdT�c�uS+�Ű�3��|�y4�h�� o"֣f�tLvG[B�#ԯ���r~�Źh�(��n�0a��h/_�jD�ĕ����X�|�3,�>}���$�TI��n�+M�yQ���ˑ������]*�P<�ěm�[+����f�P��])��u�)�!%����ɛ-V׶���p�aR���[pS����ԯ%@=�-�i����|���<?4����������o�~mGm��A�Ti�p�Q؟͎�*�^�Tz#�����w� ���=53a���$=�4_�
�hp��$�Z��Qv��4�G�eM5C���� �+�9/:�0�|��s� �'Uq�܌�&�g�̦��j)���{��2b�k��@����L�5_���K�}עo�zO��~��Ф�zZ_)�v\E8s�I�8
�yߧI��#е���e"�YEvz�R?��9��U�_�g�vxt�<�Q�O�teR�}u�8�����R�PԘ��
 ̂ F��`A]����6K<�}F��g?��w@x~]{Nma�Qsy|#��pv�[B;|L����/�� �W�'��jm]�����	�z݀܎�8�hݹ����~��/��%L���5�$ C�7�:E(�C���2��s�;yg�ί;��W��~o�*:�����������n͠�LJf�B&>��w�z�9��;��D�����X�|�T�Ja($�.m��&x�@�������d�&ֆtj���t��R����_�S~F!�ה�(�j;7s��T��r�|�o�z.���{<~�2U��ט�:^�`+��<������Y�3����u&D��G
9���k��+(#V^D��@�q;�e�K7Ә�>/}�c�{y��9�i�m�C`��_�OCu0ߦRi ����^������� %�	xU�qHI.�����x&�D<��7ٴ����F�k�P%ʁ䏤K7���)S�ZWok�6��'K9ez�k1x6��Q�'+od���T��ø+�<6����i}$�f�ʜZ��Z��?�c����drn�[�=H�ɸ;�J� �}���+�!�C�S{�Ͳ�� ���/ln�`f&����:�Eo��:w�Y�M�ͦY���\�{H4D*�S]D���v����#C�0�Ev�4\�E��j�^L�6Zƛ�~]�_�<�s���4
�˴���������}����S�Vt����{��Hsu��馆ָ�QF���o0�5�m݂��x��ɡ�P=�#���L찠먠�z�Y�,F�j�>�z�W�s��z��|��8E�]�ϴyL�������@�V�#:��H=�ٵT�&F�p��$��r��J����c�Q�_�|Ϝ��Kܛ;�d��NC3~SI)���vH�"�N��=�}W�n��;x�YE��8���`�?�%*+�&�&&:�Ic�O������/���p�O盤0"f��ɺ���ŵ�-��m��+���E�R?�w�+�g!�aw	}����k���=��-�������Z������,v�B���I�bL�� rь0��Dn�S��{�D��&М�&�>�Y��N��mm�[�C�{,��ꩭt�Q�wӉ�-*������ΑZ6$�PU��͆p���k�u0���$�Mz�\w}6	��zk1���ZY�/��Fg?�t�HҀjP�N���2���RA�H:lZw�;p촿����帳�9Q fs�����m��s��'�Tq��Ҳ��,����f��{�'�`s��?��&X�C��6��[��%����p�&�c���+q�E��l�EoO�
?��p��Uy���pR�9U�3BK;��N�(��C�8U���2V�V;'�e�x�����mP�8����x=���.SՐ�	4?d��A�����N�l�@�i�0�q�_�[ٙ;ě�	Lx�b=�U�pW�쾆إ#��=���@��q��$���N��3jU|�"���w��293��$����Z߿�0�4[��3��%�}��3\��{=�ĕu��,E��Ҟ�/��*�������+E]���S_+�p��غ��^��Le�;�MG��?�����P����ٝ]bJk��f'v�L��;m�}h�2v5W�,k� �`�6�M=�*3��@U����b���<&}B�2�Y��	��t
ۭ �U��D�qn`�ц�#�!>�~)s՗֯
G.��s}u�ҮH)*�F���7����N��n���:+/�~�R7O>Y�r�XG+��p�U�\�Yϗ��]MH�U3��M�"�~��Zl��T#e�-�B��R3�ߐ�i�/Ed��7�>v��@��i���/f^v��r�,qy�2��@�t��D�:i�
���UE�A�*��xP�Ȁ�\�bG|ɰ92)-�'t{���׺;+�xS$|R<�E&=j�@�� e��9�B�x���GM�PS��mg��r�Ϙ����4
��`��#��p��2�~�馯�/Q4�~�l^�/��Ѿ�c��	9O�:��]�����R�c�yMD�O��^��r	~�3���e���
W�����tk9-������Q2{�A�	j���n 7P�{�r������ ��͎��*q�����Ba1����2��6���C�]��3k�?d�΃��-����TCY/�f��X����^>��4��p�7E�LOt.�^��c���E}�wŮ9����!Vá@��^��c����B�3��%
�y�f���*$/�?�q���aB���[WL5xt_]-H�`+;�~��L�b��B��/c
���:]��z�P���їߌ��U�7�q�������#.�d�>v�f�M$�]��5�A���[V����Y
!����T.-�-���='L�g5�Ov�������! �[���1:_$N�&~�c�8��������������(a��N�f�$���̥j}0�
��E [y�ƴ\����߀q��%J��5��S�����@�H��>p6���%j��F�A�N'X��T�#[�\�s�ϗc���H��ئ(?ضϘ�	���H]�\޹o>�������-�^?��t7�"���O�_���G��H
��aLge��u�������f!���Ë�U
mɑ�60>�@�T�H���K�g w./08!��/Fe.�ݚ��*��m�!wV.�P�#'��pxζ!�Ocm�����)�����G�\F�j
|8�T(���k1p���oZ�n�<��'��u ݾ5���K�W
����ȧ��o9&F8_��Ȭṁ�;���O���	ԗfv�F�wM��eFD	)��0�:^%�.Cj����?�z�Y#������p헪ec�X�!�VS�%�$�����0(1��iSp
��/
';5��j��DK�(�sj -�>��F��ZP���VVwC+��FNjQ^��r�c�;3	~W�h`�����8T�L�����WNZP���k�Gu�=�i;��f;u4���_!æ�+�RO�j�|:=����nc��qH?�a��ոR�C�#���!آVPQـ�(h���)SR�c�q�BO\�ɹ�.��J�.��Uli�m{������+"�8<CLqp�Ӥ�[�l������:A�(�e��o��\�&�+%��yf�FW�DQ��`�;�kXbj��v���B����x½
%��*���Շ���C%��/�M
��h��(c����06�jګ�����2�2N.�}@�����:� �d�%��@� 9�l���i�O���+ [�F)�ns�*��n����e�%��R��<2snr����<2B�:��s6�G���C��|i�f�7��R�1����,ci7�\��!���8?��m����xFy�E������0��n�0�% ���1�
+�j���`���%�9fYp,vF`KMK�75�2�I��|��X��Bw��O��a9�� ��T����fU�D�� ����s�5"2,��mV�H/�x<�Lp�K��d�ri-��e�,x��4>� dq��E�-��c<A�m�T�����[�*��9�i6e���z���uk�i��UN��x��//�h6C)�	df+��/�f���$ ����P�b�qI��}K1i�1�%ݙ�w��Q��۩���P�=da�B�D07���m n�z��,�6K��^�����a(��VƬ�D�B�F7��ꡝg���(3����7°���������O�k1Dwg^㛙�8�!�4�@8N��=kƯ�Zs��M~۶�{�W��)r�e2<8�Q�C�N ��Df,-Q�G��yR���7�55񣸰����J���,=��	bsb ji{ >�e���J�0h�
�Pd�8�KX� {� Yu�bc����+���-�o����|iZ�(�\c�+���W8��_U{8�_�,�2��}$2x�0����+ﾰ���-�k=r}�%k����l�9J;5�+w��!t��2�g0J�y՛�ۀ'��S�h&�W����3S�'�G�p�%�� WW��	���6��¥���Jd�� i��l_GT�����>�D�y�A�A��G!tmP�-	:�O�f�Hc�� ��Ⴆ�S�4�+�� ��ޠz�*�\��r���:%@��=�e,ƝQ��@-+v�Wx��}I����� �s`N_q��^���Q�9���${%�/e���ޏf6;�XK���L$��ȃ+�!��v �BuM����WW�Z����=��\��P�������W�fH��&���_E�y?�'ݘ��=r�%��x�-��d�'�B�V��*+0A
?ea�]�������1�U�7�5B%/oUC[B���������x=�`fM�e��/�Ĭ�fh��� �*5�����)n���z`����6�k�LY��.�޴a/��R(0R:���f-����g��= ��h��$��N�N<��+�2i�tBw2gB0�h�|'�"$��yW��t���9!R�LwA�iD׾8��e�1h��%I`qt�^1<Q��L��K?/<�
q�O[���ԙ>䥞P�����+���I^���Cv��2��޳���A F(��],�W��*0���fZ�H@�=�f�L� 4��u�2�#����'3����cn��wm��o�r2������)��*��H$fUE�]C���Z`�v)G"w��9I�&�f	��� 5���t�ϲ���Ɨ�w��j���ʅ���%���!8ڬ�_u�8\�*���c�Le9�_����f�n�QY>��b�ZZij��%�~�>'g����TQ �")үæp��}'����P�����&�HH=�����S@óD<�8ʆPs�F�I|�[6���Tp�0���[�-h�5�c.I9�b),�˂�ޭ�c����W�k�kg�C�>~��7$�Z�<�Cc����3�	� <�Ͻ����&�����X�ۤEZ
-�l���K%�{J���wD:7'ˁnf������u@==����v6a��݄ʓ�@��$�θ����:�`���e��:����ꓸ�*��è&�4��� ep��H��]�<�N!�h�,W�����sw��a9j(�I�0�_�=Q�̱:Q�ճ�%���J3�k�e���(X5Y՟��c�m2�C��?�hY����k�����0�v��-�ӝ�+b��S��hH?�ц��B��
�8=���
�"�m�s ��M_
myQ�QU[�_�ug��jp�\Խ��\�T���M�Skb�5,ж@i�?G���-Wet=��nU��"� fo,�VK
40��|���O�c���<��A��s��1rF�?�cA�=C�~L#/�ͰM�.�E���'�� :������S��Z" āM��Տ�_�%]o�A懧��/�
��t8��6�����5>z����
8�7zs�0��X$�H��¡i<9��H9��8@����+��S=)[<�D��~H(�`4��\`Lj�Se�_�2O7otꘙ��{[BeO55�:c�m�p��]>$�e]�`�������[�~b��_����)�W<Q["��oHQ)���G�PE�H�:�j�V� �a>�Y�>�Zo�f�.0X{��S��mԿ���"�*[���%��=EV�-��BE܊٪�K�m+��q���3EU2��r��끟�q�t��Xp6q�{��*�m���2�B<�9H�b> c�fb��v��[�<ՖĻ���WB��X�bS���IY5^�؈w9�a�6��l&ٖ��@kL��������� ���M/T誐�g,�m�+'$�W���W���h��A��2�U	�<��)�GB�'�t9�Gk���/y�	��d�<��4�s��g2že���7!�\��t�U��[��<K���O��%��&5!����d���l	ߵy�&9�$�Oz3[1)��1���DZ#�2~TtQ<������/��6"�$���|�!t�AU�--S�M/��QԵY�N$��Bae���0t��.*9�-K�¼b*��ƅ�~�1�z�e����i�'�[Z
��x��]t/����^��>s�?��W�}��<�&Dn�
�.����9ylHK3��(��o~�
��?wba�=1��]�G��_����Q�UҌ�q-���\IDM�8m�8�܏ C�c���)�IGg��҃��V�0��^�xK[�2�q{B����@��C	��	i����f��@6i����m	����J�X�Vy�bHƻV����y���rqP\2'о�W���=2���4�+03�N\��y��|��$�F�����W8$!P����Se��vy݋.k�:��yS�aȅGv#�C;�iܝc�ʗvÓ
%C��k��lUG#3J2dN G���M����+����E?��(�	�+�5��V2��M�'�,Ut�����9����n���|�Q��*�.L؆��ˌ:�φ?x���
$Nɟ�kx��ت<��`
Ƹĩ�7U5�i
p+�"�ۭ�++1&hu�<�fI1mw�&��]�;�rčD���h,��7�s� �kL��n��7"�j*�b�A���'G�Z���� �>M����S�k�&��3�,���V6Zr6��4�[���kG�>j�����p	:�/k��Kg߭x�?��~̓�y�:�j\�i�hQ�fp��Z��[D�@�&,��p��=��B�P[�����+�F��}��K�H��E!��2]ފ܉�]�����>cr_��t��c�����;L:Fg���=)T��1~�	mK�՜9��⾌�dcчp���w�s��Qv�u�����A���H��
�>�.�,Ƅ�c��i<O�I@�~s�K��6;��F��yo�H�"�<N�C$���8�,J$���0p�B�)H�	��D��Ut<�9��;�WE�֋G��_���߭6��m��b
�)�6�V[+ T@��l��hp�լ�� Z��K��l��y��n�Oj9����tU�C�M|>�g��c�*1��Uwn��)R�6�i��ҙHb6n��,�WZ�!�Q�g��O ��a��/�$In���7��aW�
m�KH��/J�Nl��39	���$_�D�mX��H]�e��T�dns�4� �,��Pv�C���>�e��T-x��}�@nu �{��A�S�w�Ͳ�����D���8�;��j���/-��9��{,�d>��Ҍ$xp�{�QSO���6�3uE�iC���|K��R�
a����n��6��+��1[�woƖ�?�ϔnқ
WpA+�>�������Q���7&��ށ+��Z�߂�|�S��%�nƙm%E��`��И��E�º��~�|Q�L�̔)ۚ�i��-��hd�E�Kr���/X����SG?�ϻP�L������Z����u� E�:��=�V�ȴ]���&5���3��*;gM�z���N�h�G6J��{�h���Ho΍�}�(=�ŀy���Y��ŭ���%�K�7�Q����kR�-p�ia��^}���-a}��Z<�y�0f��6pO���D�]�k�� ω�)�0Hc1͝Ztoq[b�c�$:�; b=�V�¿�a�r<�vw�o'L������Q����-	Po3��9��=�YK僰#R��t���{�ް��Z�Ҽ �q*�U�r` �OL)e�o�cs4�Dm�8|�{Z�h�Q�@c�dP��S� v=N�Jc��_B��i)dݔ8!��f]�rD����'�s+���6TzL/��J��G󥤀�i� sT��+ˑ	{7�{�?�m���LÓ�:���10�$���k�.��_��L������g�X1��&����Т�p!w�&�h;h!p�rAd�ry�
N�n@yO�h�<���w�x�X��td�t���]�\M�my���/탺�Ƿ�@B������l�ΐ*o�|L�2$��:�=�e�V��Y���u2��,�1㖜9�cL c ����=~�n��	4��FW���k�� 0���:7]��y@ơb��2K!��E�"-�T��qS�江��;=�/d�N
�#�u��<��mVYӜh�!�ҷ$��je�~D�с�!�F�"9��K�#
V�!��K�-��_V�Z����.�۪��|G2Q�U3/�[���i�5�E���n�9}Kוo�A��T�vF�,�s߀��J�=�r��Xg�~��6�l&�Um,�v�;�v���v֤��	�Iو�]�7�(�hD\���A��^K��`
�<�٢�iG�w`I7h�p��C��G���^��âYC���DG�]���H1�R��t�J�0Wj[:!Þ�]^+-�f���!5%݈���%E��g4�:E�f�6�=�biPW�z_#����=��;5{=/�h�F;��)��K����D&�G��{<�\>�6�L��Q��X���G]�vL�����S$I�K�1�S��gn�d��,��
Q_IE�H��~ZcJ�u�h<�A��su�$���{�1��-F��f�"'�3ۨ��Uu��-�(;�Jp=�c%�-�����FQ\^a�z�ǵ�鎖��3A�˺s��[�
0o�8%����sf�p�Fl��2`ɕ˗�2]��f���R�nb���k���V�Z*�0(W"q7��~6� �c��hY�О(��_�	�J:��}�
k�HcߍP1~V�!���5�,w�3�������B�r��7p9&nd2.r�L�>(o����y���a���m���T�qȯ����Vv��?&�I'l�
7��7U�5���f��@`���xB�8��5�}/�_5�8f�H��|�Ls�Y
5m�e���Ge@l&��1ؿ|�m$�x��������f]~P�YR?�ޅ&n��pV,���I�<(�a��Ɗ/,Kc퉂�̨J�����%�5��n�7���u�Q����ܜPD;�����Q����2 *���/c(�o�6nX	���.��A�/��(�*����eIy|P��Ǧ%�}�ߏ�������
[;�]�^����V����J��;5S��,�򨎈p�ϙ�����4KA6�*��1
y��ڼU��������J�6�3���y%h�m=m���D1@D�+!�#I O{�uj,h+�$A U���0>���\�{��%���d��͠�3�:�����2$8��Hk��c+ĳ,���6a����Q�?Rh���a*��	V�.�o��đ�0|Z)k�>�y-��)��
m��nu͇�p�Ў����{�lV��J�w�
81��H�5�A��_�i^���s��o�Ѣ��+�\1�rY7�!Zɣ79���[��
z�M �_��r�Y�S��-��6�!8�m����vi��o
��Tc3�Ρ0��cJ��0��qt���rU��x�,+�չ��)/[���TV �3���	��0����׎��ƀj@4z ���+a��#K�Gz�Nk(!q��7J��|��hV&H �k�W�����g����K����F�����
wձ�8.�1b����I	Ђ�YD�P3!l��I9�Fn�'������:	�����r$��+�6)�{�|���k�L�RRJ���;~u Q��DA�?RK�������{q�Л���9�#����i�E��.E�_�:M����7���h坛����#e�}��4[8_�(w�����3�F*�+��}�:T*�*4v�G]��X2�om�NmL�5գQ�r�d�v֦�� ��31o����7�Ԗ⠔>���1�#���sU�� ��&ˋ��Ω���*l��3�m$�t�����V�Uu$"��S�u�A�̧r��`�$"jO�v�~�oJ)Q�'U��RB�OGW��4�����	Y1ꀯ����'�ò�Sw��+��T�� p�HXi�e�ϖ�"<q���$��CG���Εn{�P��v�#*H�7��W���z�c��I$}8o����	� ��Q�#5{��L�P%�/es(�����pV7���e��m3�~��V��q���{RbRk+,j����r�Y-Һ��j�XU�c*�x|#��g�:���
M���O��ܤp1CX�A�>QT�����b��>�wH����l�G�u:�_���i*L��bp����+��<��c�Q�ӷ|?����ܟf^���0�!;����f~t-�b�3"��x�8n�6ݨ�'���~[���vo�-�n��?f5�����iK�����rO�����}� Y*���ڲ�	c�֏Q��˥�[^G*�?�;U�CP��Z�Ln5��j�I3u�Q�y���+k}0��ݸ�iJ�qR^�Ӧ�r��	LS�$2 ��d���hT�7(�㺿��]�~|\�KQ�M�'����x&����a��	,���i�("�˭-��Њe�i����8Ľov�|�yX�d�\�3�m�R����h�5����'�Q������!�C�1����|�cF�F���
�|..GN���o�U�q�%��X��k 8{9�C�ua�$P��"^�40�+
�8̚��s�΢��DE�8�1ec�	,�޹��%�4%!d����D��(�v�؄�6V�t��]��_�1�|@ �$Z8�։��ipw�dv�
����_{���t/UK�P�� ~>�FEUf�"�|s'�<�Z+����֋�����M摞�L�Ċ �¿c�O
�C#9f�2��W������A�LV�.����v�+�v�%�8ֈ`N�a���$Y������5��`Z���X��J���Z\0�Ha�xׁ�T���Ȗ���z ^?ԕ �R���W,�G����?f/�
[��Mf�%ߛ�$4�dy\�����D�ZZ.+y��\�5���d�cW\���fU>s.���W|k��h��
�ȋ^�ͅIgm����f�f�۶�}Tĝ��&qpF�9c�zSΩ�{�&���!�i�T0Bȫ#3^-A����y�A;s�vS��)幣�d!��SS�P\�EB�Ks1l�����r7���w p�0f���W����%�B"p�NU�F�L���)��VSoƯ� k�r�~ҀbL9�Ԁj%p��_kJ�x ���	s��W��0�9� `�>W�k߭X<u_ӽ�/��m�����ˑB�e<�J�erQ���~�:���?��3�u��C�[������(u�������XUn1����"I�8j ���<�W�{W��Yh:��c}@�a����E���Y��c? y*da�l�>��4a7em�,D�+��%	����V�nq	$��-�H�wYW���eُy+���x�����b�=�*�zםr��qR]C;��zk���_���Cf�tY��Ef>�V�\е�aBL�Fur�u0�y4��;�ā����y��2 t ����a,(y�X{9��2h��n�B����W6"�Ss��Z;���R���v_۾�:T���0�ب��@�CdG�uI�b��
�np�a�QP@�:���k�$�H]U�M��:��yZ%e�@�_F��ƪ>׃NMcf����:���PwĻ��zR5C,\i"�_��!���9kYѥ&�Nܚ��@	��7j�[^�ٷ�M'��><�Eէ�_����Z��`��_v�V|ډ-���Eԋ�_�u:Y��:�� �\j��E�����ec�Ė�>`0�%]���BD�"n�'��1vų�GMΗ�а�a����_
m�#��^0�'Gn D4��YW5~	]�U�CH���߂2Otu���&�j�KLH����o���H��4x�+N�˚n=�lj����\����,!۶49H��-����(���(¼����CT��CbS���)�WP�_����{��i���6.�k���D:&s�B\Y9���F���P�v��{���*��#ͅ	�o
���xx!R2@�N��4B�Ad8K+�àw�S$�G�8���k�M��faY��-r�VΫHM�C~8M�u�Z��N��Fȱ�f�Di���'��dQ{[�y>����p)�R{Wei;�׽���h,v �T=�SN4��k|׊r2��W�~}��b���6���<����n1����Ik�� �>�t\/{+��8R޲��nk�tK߶��&��B�Ǒ�S��?f���*�ܣ�P��t�"yX���9K�SҰ����ץ�D�s��F-b�	��Y�0g��"�;���tҟGpbI`�W�߂��1VQ�I�8�5����
�H�yV�#��CҊ�l��C(V_������nM�s�؉�h�T��#�E
��y�"��W@� �CĀ]�D*���@�d�,R�~)@nfǼ���H��5�1h��W��a�dD{��21�UsOO?��L�?���E��Ȁ�c�E^�����u��U�t$�۸���v�&������:�H}GcZ2�Rq��{�_��z#>+��j��T��?��
��A�q� ���������:Ӛ�sed� ���}���)�Mx�6F�2t��l���3\������pJҜ1��?�}k�tD��@�+g>�{�uy�2��L��++��ʊ����!sk��yA�'�z�ce��#U�"���%���4�B;oY�˒�-��*|��X�E��vr����z��l���ē���@���
�g6]3�b��n;��a��&H����c�jZ�%��a�v��-����lc�3L�l��������>�G�m�Lx�_G Т	�lS({���i�7�*�J}�6�'�1u�f�����Y�Ʃ\`G�J��C}|_ϸ4���i!�F���WVP;;i�P�2CtErw�1j�^��c5k���G5��:�\ßT���|BE��p��tQpfL�"D��] ��`���
�v��n�NL�6�x�@gR�+bf��r#���-?��E5t�D͕���������W�d���H|72x�J��UV1I���	[���#v��q
���z�~�������(b6��^k*m�量f�Pn�vT�6��B��/��0�p�|�ى��[X(	+R��sa�@�B�p��x�v_ݤt)X;u�!��a<�Q�&b_��?K�^��%��ȅ䯄������C�<���.%��Chzt_:����9�[��7��-����s�1k1q��$���j�V��9ᕾ��ŧ�M���=<�a�d�2g{����c1GD��^m�3�q�
�9��t�E��2��X��zm?����W��!��Y��O���{E�5"zd7/���߱�,�"�>߱��[�+Cb�g�e�K�!7��'�sUkZ��f�,4._1�9���ax?�8��gR^��P�Q8�-#TO�g� '+��sl~����{1n��S36�J5=��.������1�Eg�y���[T�K�\='Gۆ���K��v_�jx��kK�]��se����Q>`,�J �Tk��`��-ދ�r�hp�r�����,j�����v7�йdQ��E�ڍ�Mzm3���h^;.W�(�����1���Nn�'��'��#�j��,��5�N�,~�e�A߱>$_A{����[�֔#�^�����3���N������)�}��p��d#2QQl�b��p��y��mg����v������I�>&@�o�?Ac3��9Tx�ý)[�A�������N�'VA��W��`f=y#���ZgJOf��s�V=1Ƙ৘��.�4��y�I�I�'/ge�6���nN�R�1��anG4Wk^��fXG�%[�v��7^l���#��K	̐	�|�A�"Y�k�C���Z��f�ƍ�޳��V$S־�����g�Z�{����yz�	��W�!8�Fy���g�J;x�EUaT��N���HX�����<(� '�����6�<pà#�[	�Z�-� if�OE��{�l��$��M�a�4�+������ �6t�b�N��J�-*�f�Zv_�杓�V�:�/s�z%n�
�w��f����˗�/�=/�����oF�LU9���e�^ʛ�:�c��^΀�K�g��=0��d���k��U�4�o�gX�E�焹����@.[B�Z��U�VM���9��УZy7�"9|tcȢAi"ҵU�"�����vj�x����G_���C˕p@��N�C\�����S�lc��f���sr]��EC<�a�)p*�ɕTJ��+1������eO!Ĭ���<~���V��2(|�#�M]�x7�Te�V������ƺU���tD���A�؟���6=��h�M0�)�q��5T����;�tD�Otn��<;_�->�u	�;��ܿ=����]�S)V��)�upLP���Y-�5�|k�Tw�B6��#��Zl~��A�R��x��Gx���֒�Q ��h�*ܪ�܍4��Ĭ���C���Cb��[��@4�|�P�%�h�ǭ��XBZ_��ِ�a����� :`t��F�d����1�ԠH�Mq��u�]"�:��|�xD>��(7v҇L�Y�&t����J�a���a j'��5����igR����KxlI9�T�J��6�Q�I\�ЖU��گ9K{�ͰZ��ǒBR���;檘�������Y)��٢Gs"�j�>���R�^�*4�3���ò��`o�Vҥ![]'~�e�K�)�>"\G �R"�V���7�Bȕ�|.:�P]ӡw5O��9���OP����eO���5�%ZQ;9>}�c������*C��2�9﷎�G�?Ї쥯��K���W ���8��S�(�h��拢����:_H=��g��g9{���1���`�x�գVO�ϕA����L�Q Oy{�'(q�8��\���)΅^�j[��G����e��A\����|��a�;�b�F(�s6��,���M<�ZD�N|��()>#��p���o�P�	��g�1�(Fa��_s'˪a����:L[G�5/����P��MH
7�צ|bΟw�FeQE{�q��̵]Q5�i�!'ϔ�FY�j�#�ػ	�	�����'l2P�#��TP��*D�sW��nT���.�˃r�z�`p�Ogr���� ���qp�*�%|���S1N�����0eC�>4hh�zҁ0u���N��/����U��i�����ڠ��L$6R%�l�^]b;~�E��Չ4���@�^@�����䌎O�-��R��B�p~���R�	�[�Xl��zB�EV�]Br7}7 e�B��y��{�]���9$;/��S��ȩ��pP���W�0Z����+L�Kֻ�n�����5�ﮠqV[�F�m��t����o[}l5<�Y�/�d�_l�Y�IMb��o����ŀ@������qY�-W��u�@g$�7�!==��2>�`�1�,�`�o��)�"��������6�uĈ4�t���?�_�e1T�	e� ��E>r'�ϛ�a�>��9Iӵ�AKݒr����&�4R�]S}��q��e�1�{&�#~VY�A��\y>iM=�tM�~�㟩^"�ƶ�Z &�������9b}h�Z<奰�n�0i��fM��^G�wɴ��մ��O��۹�U�j�a�ר�c��� ��&I&��c���B�Z���W��ݹ�VF;}����]� �v�]h.%�"�h��q$m��b�v��e���e?e�iM�֨�mg)
m��1��6R34�6���V��,J���j��)������`�B��Qg�-q�t�r r�^�I^y�����$��-&���8�E�҄�޵9)��m,��������Cb�;.N�LI1�������:Ĭ ��a�Z�*��$7����9jY�%,�?:~S�ĩ�r�;a��}���CC���V�i���R��}���ʢ㔄eEr:/~��\��Eg�ӊ�q����������w���wE�vaX�ԑ'�9W��V����1�Q��������0V*�����|����ٔ���Y6�����	��vV�MP�a�ngR�*y�*�r��u������8��b8�-z np"`Bs���qkw3��������؏���oG�I>���I�e��`Μ��s�S��E�Pp�[�B�;mg�^�E��9�
P�^?����A�C�j��>��R��-J,W�e��n�b�`u�A�.7spþ4��Z��g�ܧ�)�n��=�מ�
�<��e���y�IL���db��N�K���[�:��Z��1o��S�ԅ�������h���0�S8! ����.�ힼȧ[�y��'°���*�!M*K�J�>ȹ=2�K���i�����h�W���}�{u�Y,�����N!��6@�����b,0��wZW<S䭊+��j���=w���	eze����lӨ���H2�5_<F�~/`���?uvD�lk���j�W����>Z��+g�\|�I�����T>���7�
�%�&2���ft�HוUN�ˣ�́�o�:�f�z GNMT�	�4�9
���W�Q|YjĞ�T	8�\�i�Q~z�Zק0��0�V1�0���P�[�����Z��V�Յ�FA�7�'	a�H�@���!�+`y�U�S3�j��߳??�{����J��2���P� ����ʋ"�Z���R'9�����*�� ��n���f��+�a�q���w+PA���yU����Vy���C�&Hk�a��B�����h/����g���q���葯)���h�'tW=u'�N�:ON�;2��e~���S�n��Oc���݋�}wZK�
W�ZZ?!�8/��P���_�@����x� �]�����&oqM>�,�^�<)'����Xw �F��u��9�+��^|8l�X����:�� �?��m,F�5�
u�Q��`���;@�H�[e:�?�ƥ����Cl�`�������f=��4hrX	JcƏ�*0}d6��j̭N��n�Wĥ*�a��9{Z�<��r�,~�ڳuJj�Ŋ�͊3t2v�hY+A��&���|���<[Z����ط��Yu�����ݍ���V��(a~�J�Be?�Fa�#�o�N@+gq��S����^h���;���������
$F$��z�p�7�D�қ��`�/����T�(5֗nh�I����D`5�Y-Z��ur+!�RJ��f����T�,��D�R�H��&̓k?��:\���O���xC�@*�Sw<�z�"."c���,�b�q�6XB9��o�b5_��O>X}���w��!\��"�M���!�,���hǧy �j�c�q�._b Mx��fOG�;�2
�&���<A/:��p�k�No>�w��p����w$�
MѴ�a��n:�1��n������v5�#ͯ�]����F
�q����H�߄"����]I����A&��h�d��PP���fŬ�b����9�?�#8�eόjb�w���K�Q�IsL^�ȁ+Ϟ�}�k���x���h�t�61�����+H+�LT%��3�3h�T�,[��q׹�%��5�.�{{��ٶ�R�l��t3��K<_��ll�|����N���H�г�M��K��S�nj-��2X��e�3�����́����:\�$�@1:?��i�]�T��Fe�C��g�Ƚ�-��'퍓����*��A'�뙮�y��c�Z�� �/Q� ���ǭ�'�t�����c*N�jS�^�d*��v&����W,�����S|��o�<�Ѧi��O)��H��z�H�M<�p+JnW�z3����ԑ%��g3KX2��C$L���tl���G���S��rq���,b�A�ƚ��|�qa��'J��T��y��˿�s�yC<����{Բ͟M��|�<�����L�w+)P�w`z�5]_"'�޵����R0y?g �&X��'���^vG��y[P�yM��'�p3��0*�3Z����<n��iNT�Χ���]��!�N.��fc4�� )��mȭ��{� �lS?C�?���9�Z�����
 2O�j�w�2���,�����I��_�o���6 ��M
�2�
HYN�*|\���g[�z�Sx� �P9��E����	5�U������V,D�A���=�pzw�;�+���N'��ZCG)w�mӴ�UZ�CT��@��FU�O|	���Y��,�xI�e��7"�oˀ�u�s}��Oe��1=r�z#H� 1P�Ȯ�І���������9������<w��@��L;Ȱq�h�w�-K��j�R������SQ���@��\���WC�1X�d���LIx�ތ�ѹ[Y��n ������2ŵ�"Z�h�b�5f���8-��y:��� �E+�<&C�C���_�`W��}5Bov+M�C�����{�D��N�X�Qb3�K!M�Κ�v�p9I�m���*h��ݷx��G�J���L���e�,�#�j�N��"M��\��>��ַ��P�m
��o� �o'�=<���ަ�CRzH`
%��$rȹ?��I�!���u�q`�'�q��<$$��ɬ/�Ka�Ϋ�C��Zj���zه$���nNc�V�'�[�*3Csh��Vۋ��x�Tn�}�[���L�!�BVW∾��n4�:]��� y{����.GN�@�����o�+�����!L�P��Ŷ����0IP�6�nK������������-T�-3z�u�a����F���o���Y���`��-�"��a_��u��0�CGo��=��5=�WXK�-�t ���/l����(�!H��b���X��� W�Ja����n���ƘJ�tw:t:�DW"����$&>�u��~m�#S��9�d�Y�U9�AŚ�.�I+q����[�m*���j6b��6�<<0���T������,�q���"*% qvXi���A��YR�$	�_[�8����f'j�R��Y�d��A.��:�e�[��h�� ���L�^�?b#�2I�p�ȰESM ����6�H>�V#��0٩i��L���X�� =�=a�)ₘ1E-2�2p�ܖ��y��92�x'����0�:Q���P�^<1����N��^�����0�V��k�dװ��B��X���]����:��f ���@�	����=�zR�����l�H�<jf�^ ��.�YB�Y��ivkY.��| �C��[<t'�����z���J=FXz)��=l}�|Z�9pQw�*	��*������:l��Z./���"��V��O��ؤb����x2�s�V�;�S�y2�0j�b���
UJ1\hm�.�K�H�be���8�A���Q��Q}&"��٦�1[pnV15j���ݛ(��L��d[��P
Ǔ:x��eQ\�1��m� ?|�أؖ�� �t2�}<�`U�v~E�|�fGFԓn�i�yt��&z��x
�b7�q	l�o�IN�}�x���.���M���eN?ܪ����b��S���o���ħ����>Ѳ�3�W,/� +�`O|������{����	GS��|u��/�4�S��d�'/�ĵ��@�S��\��j83�����t���ϔ�+ ��'�ې�x�Z�5���i�v:v���`貳`�\1��z�pi��ȁ��r��IK�v�=dU�w>U4�6�����1œ�M�`�;W5Jh{o����?�#2��,�#���`��H���Zd`/�C��l�EH3��l�G·^��`��d��$�@K4k�Mu�KTY�nB'�7������3����a~�U\��~P,U�#,�=A�����O���ZʃI��Y͐մߛ>��aZ���?~�{�!������1I'qѭ�:H���O�o�Hԅq���֑����&�dM�Ŧ�G)(��$yh�u<�e�跀j ��U�3/�Dt� .��(��.��J@�xȲ�i�!�?���Dh$�c)M{���-!ዟ����]\$&C>_��]�{��֢<�O1����Dִ�����z+{V��a�jc\'��|��r:r�	32D\U4]{,�*1�'���Q���`x��&lӱW��W��^�O /���K�XTH�����b��F�Pfi���ء�`eǿ)WJQ���-���ω�١��"	f!G8�b_6C�nsXm+�#4�2T���]ʙ�Pq�aX9��F�F�G���R5�,#�j�*JP���p���i�y#cpG�
�c�2[�wJ^�}p_�����V���Bv}z�4�_�袮���w�_�;������˞��VB�.��i�
��5(Q4�;vי��v6A!�j&�#%9ڧ4���2�b�hd6(C�X�*JDҒI���Ԏ�W�?����v�?+]Q`ȋ�fs�+}�����x�`9�Z6����>����<Bj�巚f6�a��8c��ܡ�z�K}��a����>VM1����8����"�>p��+,ѯ�AN&=�.\�<pI�����+2`�:��֪���(@e��@�Ex����[��q}��ڕ�F܎dҨ�9�)P����)��|��tgdτ���(.m�(��Z���m2�T��8�dף�`L}UL���(c�v1n��U����M9�
���F��9�
t���S����^�©����l=V��h �m��SҜo�	�������;�^�C�e��co
O�������e�1��x��\#O��h��s�<Q�;��q��؟,��f���3z��Ts9�o��������v%�˩���J��g �ȯD;���j����jZ��B�#��}�&,Z����7��3y��4?���D��(BZ�A�2��[qGY`�����K)ͭ��wg�F�%�g	���6<�/�ڑ���(���|�׶��;�p?}BfAWI�J���þ���G�hv��E�77��iX��fܑ�U2Ƶ洟x��8(�/&]�)���p�;�`���ߚ� GZn�V-\��펼W���^�]���w�P���L/;�VI��������@�{,3��\~�q;z����`�3���mE����+ތ)s���(ȲoQIm;�-�:C�'�NxgR��${��\�wv���D!�e�����ǲ�~��d=�Voh����l������ה���{o�P4_&Eڄ�w��ﳜ�C�����Cqe�����x�˼�ׄǎ��)@>�@��O,q�VtSk:0��FP����!�.�<�Aw���C���/��u.6|ܱPZ"+��d���߃����gF��1�ȩ����9�u��vT�^��6<4�;�3�QZ{(; DA;�T4Q����ڊ&$�Tu�:��T-�ڝ�-mj�g'7g7]wc�#�8N�-��Qj q�ڙ�������WeӀW�7����z9�w�y?����kYh�#\\��@�S��ڣ<u��jL�Z$w�\A�-N���Ieز����d�*�`�[����v]�j����FU0�޿\�`Z���٤3u0���C��E-���cR2�uLօ@�Ke��|�p�q8XF-�k��yFq�N��?I"ZZ��h$��!L��W���k|c���ޫC����*���!JU�JD��#gDnz��#2C�w�/�N)Q�G�3�y��>(N�vL`M��Şn�s�ܤ�Dz&+d4�L��p���?�����,@�4[�L��=�:n���Kc�����!���j-ٿ�W�����ׅ�\MS a�a%��TnԤS�d%o�9u��do�
�-ݛ��� jF��J��.H�4@y�����,*����6#�MZ5�u��$��vr��l6tĥ���W�8$ӿZ�TGF���O߃&�3n	����+M�㛗^+Vl�]�%�r�%������>�$t�U)�T+�Y8��Et�ĺbz�k!Yd\�|xs�m�e�����=��ךf��qԫi���צ���A1��%C�b�_���\�.4�^�gC��9L�c{&p��4[(��񴄩3�Uw��\�΀��L_���͒jU2ձ�5� �)֟�@�ގ.t�<�gd	�m�kBk���As���nguBX�[(���w��3iY���ٌ�B������/Aჽ9�Ռ�j��ʟ��X*�.���'~�
$fΧh����C5#��l
�67$�M���Y�@�%�<s9<4fQ.�����?<���_}Iص�H.�@;h�<�獎�L@n&�C�S^�35��=��|�H=��������_7��8o�2�B.�C�Lw{���O����ǡ��Cחښ��s���g&p��k���-=%����C/q��vC��v�p\#ѬTW���y:7`߃"�5�z�۵!�;��Z�ϛ%�C�Z������>��Q^�X҉�H�7a��g��*A�Q`
ͩ�SCT�[��j`�a�u}��A��axc��vn�������󳓛d�L�$5^B��Xqjo��a���T}��\��ͬ}F@�̖���c�tj���s�����\.���5G���Sͱ����1-���\�����]�e0@L�~"�m��cG�F3�(��ԠN�t�(ө��Y��Cs���w[����g��H�N�Ʊ������PG�$��p�cno�0b+�eMsj�8����m���Ko(����^���yfk��')��i��l$8}3�g�?C#���uē�P�c�(*W�0,ށ�z����!e�g��Z�\�8�EE�FQ�������n͞ɴ/�Hg7�a�k����-��l�a�0� ��B�l�c`%��.����`�<�'�pd����o$��r>a<T(ub=����?ya��Lf�̅f-e���?��3�Jb"�L�?��c���h�N婙G{<���>��ob��B϶�ۣD�Yw���sINc���BT�_y��WL�w"�l���\�5 b㭜��T0{E� �������t�jR�kF\ڀ[�ݞ
Z��5y���I~���SK�Id�t��-'��t�X�<�ff��FW��PFڇ+��o�nS���,� ����$(�dh�B��r�	���&��v����L+Y�$OZ�E+�z�1�rK;��I�c>��p����T�An�����ƒ�z�Uסܫ��a�P��lcn��2k����F-��jF����C6���V��mw�e͞�eC����ɖ��m�\����Z�Yu'X���qz5��l�k��;��@��.�L�Uq�*�S �����_�6����Z�#��i�P0�3^��˱�Q"}�y����A�س�$�Տ�N�آ<���O5�(��
��+�(�V
ʆ4�Ú!w�5�å��"��c�[��W�g�Vq{ve�H�D��&5Ε�^�
��$Z�"c�͛l!5%Z?$���Q	�Z;>�������'E&�"Ih�PT�oE3p_66%\��b�bWP�B
. �is������&�� ���fF� ����mti\P.Hr�\~��zjK����X%���h�����J86�C(Q7k�9�'1(�}�TG
?x!P������ԶRX �])������|�^)�EOQz��xg%��WP���>�x�5ϒ@�*g���˸�#_�H�7�U����KLri�ax��}�פ�p�o�S�,�*�m�G.r���+j�#�VL��D�~0�r��&y����hLi/��OK<��؉&S?����'��n�?K\�����!��؛Ҟ(�����dm>�������.zq����^LĞl�cq�?�N��'+ֱ氭+�F�l�ݟ=�0��zq��iF�x�hIB�|�g
��w�ES���O��@�s���ҥy|WSח�]/�N�Ԁ��{'���60;o�k����&�E\��������x.�M�U�!p#:��<GD�U0d���:�=�  S�;�JUS���z"T�T��y%�Yݙ�)��2I��r�3u����8����,x�N֊���Z[��OCY�a�؊�Gg�3g*�G�6���Q�Qck�aB��᭼߶N/p�A�����C�0/��,�U��"7�����œA	�)kGxȖ�q#�����ģ�)� �	�q !�Y��V��^F�>���?5P�M`s`��"uu�h�}Wͳp��JN?ōV��8�x���0}��>OF4�6���'K���3����LfӐ[iIS�� �I3���h����[q珮�N�(��m �,Ɵ�t��������r�����5�v����㋄N���iHG�3OZ[�h�lg+�p�I�FՕ˜d�ɴ��0o�)\�z�%*y�h�O�j���3<�z5(�����?o)�c6��t����b�ja�+��%�SaF�E{�6��ގ"K���9�bSh@�Rcɐ�kڶԣ?)�����<׫�#pGT�~��$M�J�,����m�z&��w->�T%�,����:�!*m(U��=�q�r ��49��+���=@xhcʤI�	�~,��m�U��<���N��4J���LSs�+;����]������-�5Y�<��
�9�mz�+~��&����f�(B���}ʎ��I$|CϤ}؟Ї�G!�¸�#�1��86�<�0�	�P�	��-3+z��!��	�����Ù�I��WG=M��L/7)n������~�q(�ba~"��U��G���=���i13������Yk�|�WP��-���YW�b7m���9m$�x��衏kb��xI,@�}$7��N��$��,dY�J= �))����^1��J��e��k<0�L!Up��?�ʂAl���IH��A@��i���W��ě
�7P��0��GR�q��S�8�yl��mp.�J���{�^��|��te5��xY�预S���OxU#�7
�j����2��ȪՕ�2	�~QC7�
>=�����e���B�V���'�ҋ�`_�Dyi]ޜy8����&<W3�$Ү���]_B�;Tg5�9��.�+>��bW��X�mqn������(�(��̨�H
���;�P�O��S��~��C{��i2�MÎ�oW�^~C�tH�ٜ�x<�ݵ?M�{prC0�Ut����9���`� ��r��Ns��H5�CF;k�,����|y�.�(�F��c+��"z]g��b���@��	��
?i�����9��^.U�����m�o�2G���;h�����^}��qٞ�k�jU����4�@Y��7I�V�jQfM ?�o�_F�C�8�Nҍ��4�c9%�78ڻX��y.�c��:3z?�#�He�w`���7�����?0`�+��T|�#_�7goG���H-Y���(�m�B�D�(��cI��!Y���n�o��V��v�ԊX��Z��y��6F�6I���3��E��eM�뼕u�F-�~τ@$�#1�-;:ޚ����B̥�`p�㷆H�ٷ����,Y���������zko���nc�~�=�h���IX� <��	�6��zKv$���Ǖq�|B�N��~2<�b�ӷ�G�8���۴�Z���Qx�Q
�a�����(`���a�՝���Q�@!�h Q��;�Ѐ#)O�VMٿz�aS��e5���y����H�ߖ�����jٽ�9Ƽ�`�H{��c���X�{�1V�t�҅X��i#�f��oP:���ubC��V=����|�H�:0�+���av(
i�K���sC$ӳ��_*�����տ�Qb%�����v��>�r��%+�j��$���OĎ6�o���	��~�x�ݒK�e�/S��LQ�'�D#�ƻY�;�����Uw:~o[N=��;֮��}xX�b^�:��	-B�a��pǌ4rv���j���a^j�|n/%������re��SN��<�:���}W�ʑ�ѻ4ډ�z靟�`�~���D[ ��IǓ�5�-g��{S$M�[A�r�N}��bV�[���1�����ZÉ;\%�%�L�H��)�>�^SX٫�
k�YQ�U^���s��r�2.��Dv�2~b�߆�����A��b��S�ƿ�b�&#z?���l�T�l[��v`o"O9�C�V�L���l�֪��և�ZuU���HU�J]q�M�u	K�����GE?ěϟ���S�$��FT���0Q��,��!�9�bomc��Q�hnݛ{���?j���cH�a6�y�4��՟���:	vsZ��[m�P(��ɾ�B����DX�t���d!i�������v�P}k��I�FR)�7��­�>d�}�
A@㕅3��v7I�o C���������߰�!�s�n�Q�s|˭d�aE����M#�9nLi#פ]������q�]��z�^�y�u,:e�ȃ����L�&U�}`��.%Ջ��e�zH9#?�)��uy��¾W�V�t�'"�˟����"�/�����k:������)���_��Ѝ��@������&����i��䫸.�/��
\�è���u���,3�{��kU��j�d��Dg�T7{�>�`��0�F=�(p�L�T�����k��J`���񏵔|�6= /��r�>��#�j�X}��Eik��2�Rc9�W���pȈ}������I�J�N��	lhL��^ħ���E6��3��Yn!y׬D�C����Y!��ZLl�i��XXҾ�U.�T1�Z��SW-9bxBu�s$��Ҩc����#��x�㲐V�dȂ�0�+Q�Ұ�6%��T_X�{V��$z�{�i=���J�nY�@W���.i@��W2��  ��;�/v��9�� 㫟ħ����g)���	�czWp�
�-J��,��μl85�!�*N���j>s(x��:�&8�x��@G�{�����Y�)fk�Х.�\\�����% �d/o4�z�.����h��g1�~C�x#���S��&-�j�fO7R��׷������������⢩-y
�b���ZL��"�_�1�jp�V(s��I�_}d�����4��1�}	��Ru���0��,�m����8��N��(���g�S8�Ok�����wuJ ��߸�;2��އߣ��&l 9��5�]+���m}�����Z�-��#�6X����aע�ЛAI���}��Dm$�Hب��<4N��%"ܭ�.�5QsE�e_����cUa���#mSX.Aq�;m2Έ��X�j�B��}6�ǡ�v�~�?�[ʂ�^�s���N���S���v�x�C���'�0����0�ݨ5�l@1Sx�YG�Q8�e���P��?N�}��X�XX�����MF��8�ާI^��K���/�Eȟ��+���ku�|*��:	�Z��{8�y�JŌyY�	���!�t���Kj�4����5��8�)C+��H�=�~% �iV�-��|q���9
Y� shQ�!�D��᎛���m*�=54#Zb Џ(��E��xv�Eٔ�,��F�e�(b�.���%i����o�b�p��I������M5#��j�T�e`�W����y��C>`��|ω�p$#0�"K�
h5
n+���M� �y����aQ��Dc�3�G�+zf��Ի���7/�mM��c�q���{���s ��b_k���R2� 
�#�����Q���BI~�e��A��VP�F�V썟��l�&�J\��6��B-�l��Ѿz�JX�``	A��m��pΜXĊ���e�&�9�R�����w�,y��}�˄����`=�K~��\W��`HO���iJ�#axև܊�NFz�Ր(X�ĉM�E��ɴ-�	|D��b§2�"��JV��ֈ�d6���3.��y԰a�,an�n����ڽ�ֳ}�◓��?#���-EB��n�-��c���7�%�J�U5�����}�Q�1o��\-ZV�|�M�g�gg�����Aq
,z~�2~g@Q��ޭ��Ԫ[Y����G�ٶa�lMCtr+�������O-��D�hv���/œ~�AHh�3�@���J^��|��������	Ɖ��ޱz���~�o��ckG�o�hˑ�MZ�؍�w[�Fr%�Թ�\C`��yN������K�&������x��O��K`nbZT�T����5���͜;��U��IXR��}_1h��k͡ݽJЮ�R�|�!؄�K0�B:�$B�^���E�Y]�L&��}p�q�F�8�	�U��9�v����!'�[5;5���p)���[k�'��M
 �D����t@���;�e�=^Z���@�� �/�-��՝��d�,��|@��}����52���d%`x^�*x;�$��Xw��'g��F��cgh]GW��۴�<���/��@�]���$
TQ�W#+0 �M���k�_��}�+��rz��l�B1�b��S��J�~�J�X�IRoK�אo��ȺbR���ő�Lc9>^�PHD���7q���haw^]ĭ�x������!��?�T �J@�xb�����&��z��ɂrs[�펷'��ȹ\
�p�1��>�DZ��N��9�����R�,��_�+��g�7���A��s'9���i��!�����ůētXF�z�#��/:�Z���
5}Qk�<��[@��[�\bz���䔐��Q�T>�=�<�<���|u��
v�ՁJ�"������ՔYV8��o�ǔv�=��"+��G��<�e'"��M%�@�Y{^-\y�����$��wC�fK)�	�a?2J둹��:���>�Ihb��/d�ʆ��Me�K��E,W�$��8)WbM޹�a�Ц@�5�q9X�8�z�ħ��.|0�j��)�,�g�/�H2��.����V�׾4\cx߬�J|��`=w��2t�+Lݲ��!�Tb+��l9��G`;���]T¸����H�/�y�7��a�,�OMA{��(H�(�m_�=��a 8�����9I����YC-�X�]��?��z���1���)��0D��}n^K��c�Ic�[LDQ7;0�%��u��5@O�^�4aL��`O�L�f����K�u��� ����@������Cg���u@�)��FS����s�8@��)�1`h����{�����k�FL��  �3�=C�bҺ{�04��#,G3co�rښ}�z����7�:��\�W�p���;D�>����c`����{�.>�#��G����l���(�?�A��d�#w�ms���,2�.�����#��aN�bO	l�g@x��Ϡ�}��:@3�Al�;@E�e�Tn�$W�.�2Ay2��[{��ΒP��p���Yvv�r�f���*i`�Ekq�ɘ)�a�^d�7t�:%Ӈ�f��ģ��I�uAn��7"����k�b�`�J�븛Uw��S���biB6P���$�V�n�l`���Є1��J_�}|43���M�׿�k�F(!u���v^��+��sr����f 2�_�3�%)�ˉ�QA�ar�Mj�����8Ip|;�o�]jX��e�r�x�3�ى������9�;Vǚ0B?Z����*;�>	��l���N�<3D���O��������x&�/�0��|@�r�,?/�׳��k���rQ�%��[^��[����5ś5��No��Raa�OU��`�$<����1���Q#d�Q��I|��B1-v;�����&����Pa�؊��Z�Yr��4c"
:���˘��B��p����Tc�O͏��*��c�e)��O��3���0���T ސ�C/��E�A�X@��蓲_㓧�	�骷�3Lc�Դ
BܷFAD5}�y�0�!��NQ{HK��x>8@���朇��;��t^�2�s�۳26���J!�eM�KF?����@����7x�w5����A�A�Q�?�j����8�2���xB�F^shQ���y�
XI
XB���C�DV!��-6����e���$V��7q9�n�]�ѷ�O��_��;���%���#H�]p�-�߫�Dy��L����F�(�Ԟ���{K�V=d���zLY�c��}�I�_yl'����]B)w����uO0"5������!�=��6����'��W��be�z j�df�R�������)Æ�,u8G`PZ��D��O���&A�-%ۤ�K��S�ľ�B�w���]_����Zd'�����b{d�������EBw[F�Jm����������ȋcJ�L�%R9N���ԖA�"CxYFV4��t}�o���:���[�Ju
!h�2�\-cD����eqv�+�+a{�tu��G�`������祁�n66�e4�i�����W���j�Z�l`h*�>@ڡv��R�' ^a�����`0�d��g�.	�CwВ��=#P�<��9I�ר��B_�8�\$�k�0�oM�����j��>��t��F@�n|�g��sw�:n�cz���a��,1�#,e�@}�VgY��� d�ڧ%�P։���x��@�R�c˲��~�;�g/�;���W���7U��(�,�[%�Xb)R\C�t��_�g�,D��
��Zf��!a���14A��3�KKQ6��Zk��+6g��l�ЧQ����f#(�ȏrp��ʚ�{�UN�Sѡrp��Ld�����/�p�j���HiI��T����l��D��{M�v��>d�����f�����ԙC_��X���MF��\R�v���j�	e%��E/��`�����F�':`�����YP��I��Fs����1�5l��SLu����',E���ix�X3f7�:3Rz}Y�f!9˿��V���
��+����Ε�1� �O���>�,hX���S۽.<=ߐ�*��]��G��k`���F>���n5�w��x�x�x��F��9���Oc�S���ƿ�UnOB���q���H�،� ��|���f`��@�4 ��	�en��F�r�ġ/���;��F�}�#V`�EHv��N����mkэt�R����`kN�j��l~^>���[X3bC=�[����Зpa�%�r��?��&�?"���1[BC:���M	�+-�/2�=`1jl��\�N�����k\m}��\��d�\��Fٚd�F���T��.�0C��ĿL�q�%�.꯹ �q�%Ҋ���+M#y��ϕ�bV�!��l9���{SP�A�m�-��Ųn��C�-ӣ�R�[c�W�ݧ�g�j�����r��`�R-����[8p�ɗq���F���^���G���}5#���?ȴ��������	Q:� ƫ����
���[ �� ���9��r(��&|L�(B� ��}4�"#Ar��Lګ>�ާ���?φ�����TP����'����u��A�f+�	�O��:31����Dz�iW(\ ���/�0\�Wo\�g�d��r=�d����a`�?�(׵^eH�u��T�d��@q��,�ɦ8��m뵥ǒQ�hb��:z�Sva��\L|T.��#HQ�֯�+-�,x5�N�j�[{+*}�ષ�zh����&����[�3q���&x��!�}�+����t��dW����u�֨aF�S2,�.�`Vpa���k- ۤ���}�l��h���>�œ_�u(e��4[;3:��K�����g��4�w�C�	�֯�b���i�)� �"�hm^o��.H4�9�����A7.<NE;-EsT�VY"'M"���|
�p1����qʝ�JJ^_����ެR�z�m�����c*j�c̥�*�ܬ2B��o����ʶbn{n�@����~j%����!]/Wb������e<�m�!��C_~K����->�f"H�vjY�#�d�����P�����NI�G$�մ�<����w7$��l�����r/3� �����yKI-��jV�z�/V$[({V���N8�y���;Կ�׿�ԓ� 1�۵/�I�V c}��ˢ9tc��N����B��l(|��7��Z�,=���?��6�w��ۡ�GL�fٱ����s7�kbQ1qe������c_튬�gB;��(�pa�De\���x�����g@��S�D�W$$�0�e��
�8���������GFzM�4N�7m\J3�l	���O�5���_=U�:���*Na��5���Q#�|��T��hE���11>�> � Ƴ�M������
}�k��,'bl���bG��{�,��}��n�X�hc썇)�u�S\o����XOU:q���5�Yx�9����(��D���(,��d@�n��?q�Yc� �����>��%~]5(#X��.X,�ֵ����!�p��o�н��` ��e	UTN���{�<���+˭���c4e��M�.��]��v�� ��R˕-R�7��;����{�>��#���qi��H��/{�7�SN����c��*�a�
�y�U(f7��Y^abk=��8Mqǜ-�p������^X~S�ǰ�8s��!�HJ9������h/�g�Sk�ُ"({ӈ��E�׫�@a4�&d���3�4��.V,mt^�e��r��[ݮ�
�a��@1l�$>c��������)0�ȵ(���� ����a���Rqh��IP]k����5=ȭ�)z��"m�x1�{Ɛ�,�7��2>B�U�NDhv�TShxJ"�h	&^�� �Tp�V�2�E+	�U.r�n�e���P�6��)���8Ī7�}�������!�b �Q"�m�i�y��a���ͺ�=R�^+�6�:����ot�u�=�T�a��Y��*j�H>j*M��2���rn�.���X+|��2�Bu���G���2�D�K�T}�
����,�5�k)�����I�<�HЗД_8v�k�a�gw�^f䂧Y0�8'�=�����gG�+<������̾Rû7R�f��2��,�H��"|��5��u�t/���΂Teȱx�4k!�Յ��t��%��>�us�,�[�>���\�V�5
 �M�x�c?}E?=��
�"%���KI}2�.�2�ܠ�V-bDkn:��å-��s��
�A�9K����	���G�{rXx61�n,:�c��
�qw�n���&��v-<yG&��`�~i�ogy)�t{hU��[y�>�Yb>T���fm}����������ܷY� ���ㅾ�\�j�_j�r���u��J}��&�NL��Bf:�{<i�v/��O4�ɝ���kev:�Sʤ:���V���@�s�iIܟ��k���Tw���7*q��b�i�=�1�m�|��l�i�����8�)g�,#�3y��rЕ��e|j_��,��{�}���L�r������ת�KV��%h;
L����-�~"t\E4�8M�P>%g0���W���W(1끽�n��ɐ�l�K4��c[����`\s6�&~�\I�Sٗ�'��i_�����:�.lq�B���'K���J=���L�鿑�����,��'α�`���k�2m����iJ��M�4�4&�?ǰ�� �\V8w���d��grL�Gd,ϱ�oN2U�ְj�ZM޷�Է{��攡�;]wB@u�#��ԍ��zGx�F�k�M�{nl�0�Td���2Ei�V�{Q�h
�_����g������}��� ����i�_�`�-)(��B��^�8n��0��w�/_���XG�s�R����e6kK�Bm�dχ,�����{\"X�f�
�Vzr^��4�C󍉘�5��o�}����Pb�����".�S*c��ef���>���Vdu�D��1���02iJ�G}m+�ʥ�kΥ/'��1߆.��k@��Y<a���&�7?�T/~�5r���0ˋ��a@*;����c���yl�&^;1����
�D�����D�M�"�ٿ�
n�/�L<_N��<��-��(FU
���Z�pܐsb|_Z�xZ�0�17i;,�
���"�\���V�\�2�m�Z����;��ɒ�&\�r+�h�(]&�c���-$��"���
d-T��������}���o��z�O�;^���C{W�!��Y�,;��v&TN�h���� )�	���슕r��bS����>��&����r.����9�,0�8�1�K�Y�&�yǶt�$�n��-����q(�PB�sԛ� �����ua��}4�C�L�&��@��	���H��j�y����ډp��Y3Q������F�QM�a�L�%�K<RՍsk]m�'P�J���v����0�+UZĹΧ�˲��A��8ޤ�)9����ԫ:��x߲8�x����C5���+0aG-�Gx22&Hq�������)Y��,9v��ħ	3����3�%vo$yE$�֤����	|`�O�P��ގr
K���d}�*
�mU;�<�,�B�>�"$2��b�a�a�����(��f�m�aN>L���O�	�"e��u�R�����]����AW��.�{�~�'m2��s��������i���[���><�� ���#��ra�W���$�m�2J�����N�/���r�n�\�5[bn�T��*�b��!�?)��vAv��H4��pn�tb�����&B9���I0L6�}]�9H/���ѹ+����E�Z����X�MryzX�Y�3����d����Di�"�B�T��)�Ը�ԫ,0�����!�%��?w��z����Ïi��$��B���$��r��f�.*&��t�\���=�f�;��)P'��-&�� �7M��)z3mR?���#�`���`���=qӌF0:�,�#��f{WH��!Y��_5�jF���Qqwk�e����T�渗����E�rs���K@�u�@V�d�έDX+O���d�������?�O�׬��C��&��LG�L��:��7�R�4G�O�_5}q�Z[͈	���ɋ��8yҷ�ȯ6  ��nz�$%����RW�<�a�c��p����PAC�˸��. �{��s!�k��c�9G)y�������Ę��Y>5XO�/��$S����Z�s��y�����3z�r�#�u�o��dJLC���,�.~���un1��(�p��~IЄ��5���q��:��l=��j�&� ��P|0�F���2���0trq��J��yr�����/a����&4�K�H"ছU1�Jd�v٤�/� ���Au�F�}7�B���|�(x�b�3�yFñ�_�54ʺN7�Toh�t�r�"�Yμ�]�Rg��4ŉ뉍"�����b����`\�#����݉�3qh�.�����os�d6�����%p��[���!��\��8�-R�JpЮ�o*?�iy��B����W��� ���.Gשd�/ l��Cp��=κt��[e�hmԮP3��%$��	�����f1H5/ݱ_&f�M�Q������H�}3?������]~��K����F|/v�o�n�_<��!��	G.����� ω�T=�Z�(��b�g�]�n��ŧL5�-����NQ��*�lb䫹ڥ�?Wl�7�;1^t:�&j���V�*W%�3� ���F�B�]��O�XWx)�*AtNY�3Fn�h��V�m��Ug���;�����������F�<�(����V�����Oߺi�wV:s���n���gvF�ܓjk\�NFhL�׮��v��%/e�ռM����GI�V�ۧ�HZ�5��nܠ�)�wت�;�&�"z�����j�lc�I��XHP�����æ����H{aX �}��ٱ�ެt�G$��z�gC`gҝC��XہL𔻆: e��?j�a*��m�@}��|ͮ��������BcB�hhv�%�|&�:{�6�����O�ئ
X��Rq�%jj���;ځ2��\�+����lM���+l3��OY"�C��,6Ж8G���l9�57��H4v�,TʓI�6��Wq������q���Cu���{��)QN��w�[���$},IXF�i�&��ґg�oU\�,��Sm�I�����/,9wnn:mU]@^���_��$����*R�p
 �%����A�(�/E[B�N�@�U �� h�|Z�hu;5�D9N9\u{T��_	.ۣP%Np[N��6c�%�H,й��<���V��Y���.�ǟ�En�-C_f8�!��VoQ��6�ISK�&mU�$�ן��i��{bS$�5V�k8C2X�M���5��3��Y����1��Y��LHT��c���*Ld��fe؝���d�Q�f*��o���&ڬmYs��$�L��]�.i��-�s�,�c�k���$	��!��Q�Cgs������OP���L$���'=������,���~圮����a0mZ���%�O�4��@E1����Ei,w��ϧ��T4��2���q����*w���NMNވ�2d�@B�0� ��8s9�hP��L���z�����>Q�L^45w�G���W��j]�§��*F	yи��;$��g9�\W�Db���D�B�?i&Y����T���0�I��r/f��T6��s��Ͻ��~E�5��5�Y���n��|��d��5�kHb?�r��(�e���?ם��QS@�J��2�I�4A:����p��������KA�vu��Z�X��I?p�����?��V�]���%K��"�'��ϡʇz�S�=:-���Ưߴ�o� �K����EdA U+p��j<Cg`םD�����QT-JAx�@�N|�.|�Ԍ�~��$�6�M	�#8[6zf�c���1d��z��8G�	''E`��q��G�-���-�J��{@��L�jV��^�-�dH]���f���w�zp�j�J ���7z���+{�F%����}o�H��S�SHmc�R�|��@^�J���v�u�P܇UCG,��x���Bs���7A7��c@�˸1�����gT��V��"헃U����Y"lX�5��ن؂�F���A�8��;f��$~Ai�{J ��"e#��Fj�'-��=q�T���W�
��^���"߯0�L����l�j�
��7�fQ��`8�gz�A��V<�Z�6ql�T�L��(�'�H�40�O ���<��,�j�lZ{�ښK\�YJ��I��> n��]��R�4R{2��'q�AH�_�+kv]�l���/�AL؄��Pn#�N�wI�:����Q�Ø��QfjkE��.�*�(g�shh(8|>WN�n��5�qH���ܖ��F�Q��r�-
Q��m��F_\$Ji��,勨3L���R�j�>5����VTV|B���gwJ�߰j���Ls��v��=��=w�"u�&��y쪶���P�!�����M5/Y�����l�7�5T)���t���i2���;5H�L�q��}JB�栜�oD-���V��<���gO��R
�uaT�*�	p�8��՚���Ag̷�"x�~�ZsM��GBz�կ��R]�?N$�b1]۴Ei ���
�{8�
��'\~�M4�}���n6�-2�X\���yl��7�2�fg�RC���{��<��~ѳ,��<C8��Wδb-(RA9G�wN�e�&���˱kJ�Df������q�l�i�iV�f@U:}#��ܓSm&F��xj��~^�J8�#���<�C�n6��d���{\@\�3�c�$Xs�6��!v|�2ȵR����Ӫ�.ʥRK�d0z_Y����r��fD�a2��[�WWad���ax��1"VQy8֫
<�u�IO�u���h~�ᱩ1���֡D}����3�SGk���k��q�L,6��x]���������p�f
�����<�f(K_��źt0oe���b�d7X���������*���F�C�ظ��4��(:]*W��I~J})1�?��c.0�Q��Q�<�������:Ǎ���7@���X��yg]���j����;:_�&HT��+{�}��Y����+[>��c�U�/IH�l;QeIfZ�k�On;L������jZ,��c�v�KJ�#p��<�$ճ����ɗ-ݒ�`�����Vnq�LG��|�B@���?�˯�O��sp�7		�c�������)tdMT��(��q����{���^�+�D$�M�>�N��bSq����:S�:���ԭ�;��	%W�m�T��zn�xp�������[�C89����h�)�Z��/{�aƭ~'4��PC��>M%���f�2H��'�v��	c��E�4�4�l%�]G�T�T^jw�?��h�B��%�����5 �0)F�-/�j��1�4K�������C��g�L���S���Jf�|cFE�E�!����\z���ͱ)Z�U�>�B��Z�{�7A>��;���Z3p~�{����u����P�S�[Xۅ Rp,��9 �??�>����>+k�4�w��Lr�(X�o�ha����#6l�f�9I������o�ς�=��C}TĢ��s�d{��L��\B��K�w�gO�{uI[���D�E�Z.���s��Gc�uẠ<���"��ѹ}|K^
\�x.ba��:}�MN���B�!O�:�t�:��������j-��$i��I�� ߦ��pP�,��<�Q��K�]�).
�5T��C����֕��H���O�`�=�n�ov/�aOW;ϐ��&a����//�s���Σu5dLC����&d,z�5 �M�޼ ng$`~�Nh+��'x<���M��Iq���4$5E���E��V���a����^	*�)]7�Iϊ����3��x�0j,���l�	�c���"|�M�k�"�8��A�ڞ���J����}`6�h!��b�m�}|#:b��*�ﰿ:\E��>�KF�q���Jdt��,�q������E�������xMӦd\v0؂�7��՜�M�4ȝtnB��Ğ���v�^d"���.K]����ޭh��F_��U�a*���6��-��7j��AW��bL�k	���ò;~^����/3`N��&�9\7��R	7�}�Ek��`�P���ΐG�ړsy�hr$��@�ß��:��Y�e�PF��_�M-�7�E���C�"�Ohp�Q����M���)5��Kt�R�X+�D�A:����9��:|��Z�����M��W	�۝B������"*=U�oM8rO��^��9����c�YEN�����G+ٙJ���	���Oz�־���&�(�e����{����pl���>w�Pj��2��p���e��4m��}#7�2�;N Y262����0���ċ����%P�w�:�����e�)kF����|".Q�if_W���g�5������7�^ГB�O8�i�P���d8+$�e�,�qT�7$A�;�͂�&!��<��8�zI
#(��B|�����I�'ܼfK�s
|�T���`��G_aT����u➓Q��$5�4 A�$�囨��t��^�"����,8�������O��_g&�_�j�35+}�H^��V�Ė�v��>7r�|���ca���C�?s#h�� ��+�M�+��ތϖ��J���b�US ���^=�؞˄�F����O/ޝ�ڬ���q�KEKQ'jn� ���5�$����oM�@���{-�K:"�E�G��[��B	�94Ѵ�KB�|p�����S�����gA�ʐ��f��z-�f|���� R��[Z�1�fX����I��H�GΨ}����\��䓞�hc��T!P�G^��;�-����q�kM|�C�G��53+?��F�����0L�ܒ'��i�n��o���-�t