��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]����
3�k�?�����Ņ�{{j�|�Ƒ�|�ݸ�x�l#7�VAe1�6�1/�c�I4�b���'X�6�<a�y|ePx�����?+X��gK��f%Qh��l����D�],��	�f�<�ZAWl�g�����4A�3=(۩�W�OC�&NRөQ�Ҵ�#�ͥ�|����S�Fo�'Z\��{6��a�n�F@�_�e�د��{�|���\��1&A��dY�����פWY�}I?��,jGX���>�bhf@��ٝ�,�8n�L��I �/�$���!�0�^�k��5��<�E�Q�#[ڟ9�a(6%�!���ե���c27+J�ݱ���J�_���TYxV���<'B�a;-��+���fM�	<�ّv+^�~���K��q��/�#˴͗a��
\L4�OP��B[��K'lYA8�׀��� v����7�ڋ�s��:���}BR����Gտ꺎�$>��=ꚐȐ�dP��+�&���g�-���8Ůz73J-8�k�S!D��@�zF�E?ق��8��Z���Ss���?���U+0�|�	��}�\T}��8@���ga���	P���&}�ҲQ�g-�Yn����8�V*JnCMv@y5]����r����A��'2{P�#YB��+��d4N?�'ߩ&���z@�k6�^�C���ܶl�����O�����q�bn���1���_8E?�p���K�Y����Wg=�O�FDx�F*�VS��VD�Ŝ��:��`ΒA�ءhIw��98�s彶�nO�ԙ�0!�EaH��m`��W{����	V������}�5@F�-��ɔ�AUEhi
[�>�0�nZ�=`-]TD�h�� ���u==E��A�ny�11(�н9�����h�U/蜂�q�4�3(���0��Mh#�(�{�������rһh���Ȋ��9��SҀ�F��-��yt<�v`�KW��؛ȼ��+y��;���b̏k��0�}��'�;�R�{i��Ox&Z��f��Q3]8�B3�J|2�-bl������A�7EN��
�}!7N܁:||#���-�\��ȣi���'�!��TW�t�@�h�tkT�z�� �^{�)d�Gq���*���sr���z��/�K9~�-�|����6k�>D�-�8ES�ǘ� /�O����:Z�M�2?�"�_^����16�VKS��b�Yy��.+X�eɷ�~5˧ڥ�*$���tFd��.J^�P��Λ�F��x��ÊP;i5.�ߔ�O�lX�`�����8R\���=��:K��H��!��N