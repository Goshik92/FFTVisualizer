��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv 6�$���m|9�μ��:q����H�r�4�A�����ls�w�"�E~���Z�ޣ��IS��K�l��ĜJp������2Q���{
����qˍ��|���e�����g�R��hG�"	�/��,+�J�=F	�k�@']K��lx`Bp�&c�Ux=����I&�ŀ�"fԫ\uaW���B�L�e}2�o��!��%86�ϿG!��kq���m�A�Q��N���_�� �O��C#��r��Æn��Z��_�vr��GӫR'�������� :ƀ6.�-��L����ȋ<�{i�9�"Գ �$C���Thn���]j�ر�j���$��E����	�~2	�t[��ʪC�ܕ6K�Չу|���z˂��W�7�����,��IK��&�������,l�D\������Փ��!��Q�ZRD�)���n/���<��<ʔf��,�k���^�	�[���B�r3���ā��N�:}�����ܮ	0J��Q��dTT��L��g;�P%`� (��_(0�oat[��ڔ�_��{j�&!����̺���Ʃ��$ƅ-�����QS��/�Ͷ��ʨ��Ya�Yypvr�N�3���u�=ˋK�ܦ�rވ�t	I�sح՞?�zy��Y���ޓ��ǰ)�l�Q��K�8�ps��-M>\p��]��˂c~��:2IM�h(�Y#D���}F.C��&��e��D�d~�|�c�\���gD�cS71Iӏjj��ڳ�"�t�a���x����`�t��HO��ڋ/��L���%	�nL��"�g�=O�@@�D����q]��R���$VD�<�s9�~p!Q5r��(���Q�D�C>{8d�zp"c�:�W�@��RaLjD��v~Gs�`�3�-i��.����G���Cy����癖�%����A��O��sq�Mk:�Dl:��y��J���A	�����I��Og,㤎��j�J��x���˜\�f5� �-(�ďw��K��*�!;���:�����ч�B%�ly���;g��-.>����4�߰	�-)�&gA����4ﵴ<�z9$�z���R$�8����Y�.�2fI}:��TAM���?�2�}憧I�)���T~q�������:SD�zW��E����ܱ���:9fH��d�ٲ��1��l�<�\�7��%B�==�XC,���=I���)T�&J&	�J-�.ZS}���=X�-wor$�}8F��2�s#%7C�u�o�={��8���^3�*W�0p���&��Ʋi]����������s{�Ͽ�Kb�K�����oKȡ'� +���K�z����ڻ\<�2�������7C�s�
���e���i��x����E�"n�ĭgtfr�5=��3���'���s$�ɣ�E�����T��E;�S�Ȇ�q{�+Z��xV�"�vh	�N�hZ����t�B_�ǭ0z���WSh-�5� ������������$��SDn�'?�^}I����~���X�?�i即���vI`
6�2h-`�[~D�	Լ/ͭ�*;){`2Dn�"y?^�]씨���_W�\����h��}���I�G�fw�� 2l۞�B��L�2I_4}���� ڽ��n$꼕�!�U\��a?����	��A#ir�ѿW��^䃽`p�2Cv�)�ά|��q�6ڠ(9�N�~c�=8qKxXS��r�w��A��̝��\~/qs؜��V*��b��(H�E�X	�*vV�"#1�?�*?~���{��m����Q$*FM�g�^�D_��o��Mp�6�(�'�]A����o�W�%O�톟�N�x�e��,�M*Ά1[}��x_�Fj��� ���Dt��
�$�q��>8⻃�����9�+U	��3�e��i�M�~ʂ}|)�#b�]vq�ד�THX��ٳ���A��!'�����@9|r�Knhb���G$ؼ�Z��.���,+ϥy'��@�����l���zE�U�8�n�w遺��{A)����{�T��D������M��d��>�E��fe���_uc~���`�6�*s���Q��Q��7�k|�����IB ����l��A�����qJ��(}t�w���>:��s�,f�pb�\���Ց��(�眤��)gn>�5�5/!gU��¹r��$�	�<�L��2���ؙ[Tt����h���B!�M�As��bǯ)j�b��w�G�i��e����H��h>ҵ�j��ƄI����(�K��~] �
��i�ui1�){g琂�)/t�� O�q ��03���g����qOiB�G���h_�3�d�����{,p|=������M�YA$��+$����-�� ~�ʣȫ�H��L�c Ci�$���*R�@g1�#̀3�ߋ�g�A��
�M�in��N��˩��]�����}�֒���(�!���(5J��9~%�	��|{��''@��a�إ�F1fDWޣ�TP7b���Xh���J|�|"��j��W;	�(9�S�j'%͚�6�h�~��{56aZu�GA�����Y!%L%���T�`T��<M�4#g��ݮݱ �=h� R�7	;�m��Q���k�
����h����GL�C��EC|�05.+�!��-��u^e���m���-�e�B)�oB��ʇ��0Z��WjC�P1n�&
x���[Q9%�� ��� n�4�V}��kVG�Z)
z�����;�2�%7᭾6��C�[�W���v�� ��q����y �Rn��k���54)z�nҋ�d.��ubQİ��P������QT��i�f5�`�3���!g��3"G��pg���Vɛ�萦��S���'����p�����͕ZڲM?)���vZ3$';֤zkT%?���8He%Z�B�w�$oR���d6��`<X5D��1���ծЯ�{5W[<��K�$���JXy)yQ�`��d'��)S���J�b@�g;*7T��F��,������o�LB����+K�v[�/�R�)Z&r���Vc�m��D5��%��KA�o��c�آߧ���l�d��W��+#��-� �k�edfS̟DbaD'D��;�Y�LО�YT�]��[�k����ˀ�Jx��Cc�	/nY�ј�7�Q?���x�C13筵���E`��c4w������K�5W��'�L�ј��i�%F�ߨH5�GWKBJ{��Az�Y	"!m��y�(ُ�'���u#`�}����n�`�����D4҈�1�Wej>�O z��٘���=N#�v�)������t����Rϟ3�PUxK7���M��,�]-
"ͬ��3�0\��L����ޕ	o�� /ws�� (z
�\�5��-|Q'A���Þ�&�
N�ƭ��m��(�4����D�D��m�׆����#���*fE$U4�L�"}����=H����"6zM_�6���M�w�u�1L��k?����}�N�^�>�R����[��
uW�]/sR90���k�����ʢ!L�
�I���5`����E�R]�o@>�{[�H���ojKfWb���W���ׄ�8_�Y�N[u��ԏI4k���C�תP��Ο�����{|�$g�I����(mJ-l���ȸ��ט�l�7>�HXo߾~��(/p�z�����_��c�r[������`�U�n�u��D�څ$ ACܝ&vӘ.������X�f�qa�2��6S� ����K9/�/�?r���g��{#���9ͩ�DQ�Α�]�C��,S�Qe�ޟG��]L���C��m�9E��[�z�{�xT������z��v�K+���,�����Uw+k�V�\��ۉC�MYǻp�$_�v�Qgch��}��	���R��N�)�M�p�:�5Dw�z�C��L��$T�`�V��CA!�jnv�����O�iU2Ow����jb�@���������@���nP����fp�����0���7b�B�[�whS4�z���d6��$�]�5:�V1]�$����� �\���/o���@��b�"���Z��{ǝ?yUv1�����C*@V���v1�����:�@0�]���du�h�"�z*���#C�X�:wu(2`�1�m;F����B����T���g�.�Ó�:)7�Gb�[b��lEU]�Y�  ���9�E��(�qX�@���#�:<��R	�^��U��~�󀌯�-�����%����0���(g����k ����=߱���Q̨YX�X��Uq���p�����-�"���Ivm��q�Ǐ�H"` B�qOc�I���p�ZYZ3�<��I�R����5j�^0�#V��g+ԃ�xl�>���o�̺��i���3�Lк	=���L�w��0o�!�-��.��ku���^�]&K\��@n�G��=�������Q�!�2�}K.c/>:"\��t�&Dq����םDp����v�������g������� �*D2k �Oĳ���10��,Hfr��_��J�dQ��3a�g���7�����Ӓ0I��W�y����b��ʿ��o��E��J�C�#yM~Ę»Ƹ�;��YM�ww��Q\�i� �^�d6�&gU���H��dɈ#�7[�aFd�"z়N6~��۷�莦�fKy�6}5	q�D0��s���~����[���N	��j��X�{O1e�� ��Z0��_���R�	.�صg���k?��Շ�lB��i�[۩�Ĉ(%���@��!�f��cCy�\S��G�8C�l�����̸@�y;���iL�-���_��V�,'��6�D����y�[��!��]�ۻ2>�8{�����>�fl����c���$���"�?a�\E+�B��J��W�
��툲|���)�g����̷�;<����0K�go���RL&����í����/ώ�*�r>/Zp x]�����g��d.�j ��:}��� i���em����!o�>?I�#��ݵ�<�݂����Ă�h�I=����L1�η�.��z���B�<%72�o
��ȡ9+�F}k"W�:�������#f�ѩze�~�k8w1Sp��?�[F}��w���j��}�;���)���-	��s�A�=�]�*Lm-��wD;�����Q�֫����*Z튗�Η�����՗]{�bKnbx�� K����r�K�;s
2I�G���I��{a��%�g����b���q!T�w�E9�eL�d:��/��c�8�;����Ķ��@�%�v뤔)��2��3u&%�y���jĘk<�]+$q倩��.�	�jEB��A��e|����y=���˭�b{"��]�4f��f4?����<��@�R�|:�(��h�'��[d�>,B�hv�c=��H��gb��ѫ(�D0֔^﯂$'�]L���d
~��X�����
�\H���h�4sF�����R3��͠�6�|o�oC����=l/�YJ{���Ҵ�SP�T����ZP�a�����UB!�[���.N��\���x�r�O���.���t<�SN,|J��b�X��M&��}���K� ��"�)t��4�X�_ϊdq�ne�Y�� "}�7�b�JF�>��\�u���D2����=.�<R����N�X��`�����{H��ׄC�c�G?c�2JuY�xLK ���wa}����J/W�r�H�F�-b���+H�h�s|Z�6�Mg�S���������qb,�����9 O����n���J�Y�e����Hj����6��^�G���+P>f�Yq��j'XR@}A�����L��;��W ��0���$�%@�!��8����*3���Twr�HcSԗ�rΰ
!�j�K�
_<�K�C��+�����>�G��Y�l,�%��<��������R�I��}$B�~%Y�1E?�^9K0Rf,��A�LRyD���������A�.�GSK�`��f-�l�F�Ѵ���b[I&�î����K�'��3z��Ö��s��F�7��[��P���7Y���6�ܷ�*��Q���B�^�a�����_���X"9�|��P��Z׫�W���Q���=�,�]���j�R��UrqY�<De�}���peM[���^}ϱ|$vA0�)�.���ζs�r��le�s>@���/�3>��" �N76�8�"%���������Ӱ,D����%Y�C��";櫯�s���?$yП3��j-s�oS��k�6�˻Ο.1���g�z ���TN�+�HbxSU�4�G. uW������0'yN���g��B�Y���|�5L���+NI���y�ޒ�ƽ�g|g�F�/"b{οK'�蛚�0N�^i#����!U e�Bǵ�?�7�l^���+B+�I�	�V���H����Kz*+H`&�R�ڪ�)΂�j�l����{�de���|�6ua���v�����e_�S#�!c��7g̪#���lY[X��6M0��Hje��_u�(��3���ӻ���*�ر�l�4�.�Zx��8=w��O3���2 ���}�R�_�Υ�~je�����\�j���B2�>5k�ѷ����R�K.J�%�hˏ��-�r���*��hC��G���(N㿎�
�v��Cͪ*�����弑�8�C��Vb<�}����`�Į������:DF��/��%��v�v���l�´�%�O��͇!*����%�n���h���V�р��#ҕk�"S�����p�u����O���p�� H�S
rW��ylj�l)<�>c�V�����꠬9#���L����[++A��P��V�`��F�)Ǽ��;���_u6�6�JMƦ�I���G����Y�!e�o���A}�i���Wh�H��:�V���>�_�Ue�oí|��V�wUy��G��l���%�A�㤣��]E��PYw���/2�o`�VTzh�%.�	�hՀ
gt�����tO����M�Xe��zj�|]�[�,�Cx@�>a�}��%J��Ɂ	�� �讋�ĭV��&bh���)�?�]R���H�,@��S��4g��mk�-J�˂o�W���e迟Ml�9ζW5����<u|�/9�[�}_�T��3�1G���G2�g�-��ۜ�)iD7w�lY��P���zd0?�A��A��`�Z,M�P-�W������ҳE9��ya|���r)��s���0Ji�����@ݼ��V��$9AK�0z��d������
�9�E�>�	<5�kcz� ��\c��� )m0�:�2�7�m�=E�;o\��Bx�YO���O�bO�Q��|n`yXZ$��6"�i�ם��Z�DF��Sw����Z�8�X'a��K��N�@͝z�u�H� S�h[*��	�ş�ɟ=iL5r5�G����U�$#es�4�R�M�!,u�9Y��PEԮ ACD��H$+��єj|�\��lU0��lR.�RÑ-e����X7e�\�οN�)mF��|e$OLΓ��r�7��v�C��DK�d�s�y���E#2
<����?qe[���e�r{��SV�Y9;�z˕T
�
�a�+3��*Xq�i�to�&��)>��a&�p��x�����qᔴ�a��" �����2��`1�rw2���K���`��a0�<��G
+x ���P�x�^1��s���Ÿ�m��2W�>��Wu��.�P6o���8�*�6��r��diaG<���<y�5��}����S�t�d�!��e-9�x0����钧~/���&���SX\��¼����^G�W���o G��t�+��ϗ���D�z�2����On���P(��r��Ԣ}��Nr���Lb��.����eղKB�eP?��+'�����ˎoVf����-�(	|/�aXP�Ͳ�bx�pj��I�K�ι�QS[2f���U߁�[��{�:�Yz�B���0���Eq�BK�������Rb�μ���n{iZw3�.�ZP3�Z�b�A���u�4��[�ʟc�v4YZ헮���G S;��`:��C�ղܛ(�?U��S�%�6�:�Ω���Ū�@>�k�;���\[����ҿF���$���\��09��o3X%�)������#�.]�I����v��Ӭ;�V��f[�������� '$��U$l�A8T�0ڢ�<!�=H#�)r�@.]��g�B����X�>+#5TX��sB����z��
g�L�����ף͎=�t�g�=��Q�b���}�����ɽ�͙�B�3�P�$���f��e�"�?��6Ƀ��I�l~�l{��� ��噄#��V��wQㆭ��C�讣Slw��b�
:���kے�k���M���h�����h�3�(��(�J���IM��)����G#w�ɿP�'d,[0��yj�WCɸ�0Q�;���x�'������߾�4n@줠����6��`z��A���H������H��p��FD �-!q�dV
��(��g��� ��Ȓ5��F��pun��#�)�TC��w�//�<dj]Y�10�/hEиh�� �?ɓ��A7�W,$�V9��&{��uXA�O�s}���t�.�[yA|�6��l���Oy�F �V�VPf:��V��JO�%��䙫���0mG尞xO�(��D��e\�?%���8�^�!����r�Y�$�e�ĩ���@�<PKe�<�KY�6C�����W�{c$��'��̏l���&����IT�Z�>�R�Bb�e�M1�Uh�hr�J4�ƌp�
O=���h���s5�U
ns2��=ޤBݭ2g�V�>M���}I!�����Y�F�%91�����噗f��M��ei��	��ϳMǱ�ʎ�Y횦��:"�ӔD����ʜ �l����ǉ�Z�Vrr�k���>h�s����I�ט�2iD�X��{�a�D�ȏ��y]jD�D�S�8e!(�pԁ�<>����YS�O�y"�Vq��HN�������R�<�d��?��2=�Q\2@B���f��"�'��H����6<���_��Tl�B����~���M>a0�X�5(��Xy��:@6�&��D�4�+|Q��ܼ��,���1�'���&��J2Y��ِ}�I��W9:@�.���u|�Pʄ*���(���A=�� e]X?\Ҫ�M�xi1��N2��7@CS) 7�ί���CD`����ꏻ?��8L��oCUן¨��ۂ�L,3�]�*(���a_�:f�VY5�5S��)�n�9��NW�5q���ēl/���#"j  ۾v�N�� ���:�D�c<f�Ѕz��'�\4�2�|��i�O��;���X���/S�� ��A�\&��MX6��7��?�K��U}��(n�%;��w����٢C#� u�kK-\,�/xs�o����Q	�2?�2�ۑr2Xh�-���|��ԭ�ӗ������41*�,�IYU�ǵ����i���}hyE����PT���Wm���Ic���s.\�� /�|�� u��B�P�0��b���3���iɣ?촓��AQ��T�ux��S&߻���l@�,ek(��2p��'��x��:��ݫ���
l{us(�~����b<��\ �=(Y7]��j��(6�;C������������[������'{ �D�F/����L��ƔF��jTY���J*���ae��p:�&�Y�zis�b�Ig X�	E�|(�LY2%�!��x/��ߏF�2r?��/�)���e[=��7C����!?b��w{\�6��<�d
N(_����~�\=ڻ�gGc��A�a���\ry�J
$����[������?4^�֧`&4ҟ��j�u�ͷnuE����x����n�tF��X����uo�-%%pZZ4nb;����X���b��7��͘n�Z3�$l��d)��Zt (K���&6�ǯO�g��N��.?ݭF�����H%ө�,�H�)A{�L���[���pe��ƥ��O���rY�=��%Y����x�He�c��A����>r9_3≀ױ~�s�Α���
���(��q�$����H<x��Aba��[�����W����np-ٻ��CP$����K��Ѵ�U~Rf��Z$�9 ���P�0�7�ct%g�e�1��:�hF�J$� ��}����o�.�aL����Wu��ԓfu.X��h�90SA�f�SB6�"�%1�Zaɖ�_a+8�@���Ip
n�0��!Ƅ_� e!Ph�Ahy���%�̣:�u�g��'��a�TҴ޿ϭ(�]�IC̉C��Y���;C�k���_K'�V`�\[q��߇ӹ�`	ɿB%�B͟3=��L-�x�����|m��R$)�`����0#�pB_��,�v�i���jp,H�")J���&+6Sr��(�QO�&�z��땛����>��z u�[��k/.��� �����0N�Af���I�ɥ��I`��~�*��-��<v�J%7���}X�%�k��r�R�W
Jqf�#N�ָL����s)�W�)ח#ή>�5x���u�#��p�����T��>N�_��f�8�Z���V�W]-�Sb"J0כ�s�Tu�o�S�٩RS'2�L��������FQ[SFЈ�R����"˱�3�&�/ =� ������ms���r���Slb���7/��� �IB�VL"��������3��׫��gHzU���'ZQO��x���\�*�,-�5#�#��O��m��U
y}���v8�J^3
� `����(m���*@]zҌÈ�ss�,�?�&��_�i�($"��PƒMIN}��i��_�~ѱ+����
����w���R�`��'�Df=d�>��SЮ���};p"��]�R�M�O-�|��Y��o:Cl�m�!�[~�<>��~�V�3��2��q��� j�5�9���1�n�-�}�W�l�g�޳`�Ņ�Jtxñu�0�����Tj+HS�\�<���,�(��$��CD�T�d���ARUL93�9�1Aɯ���� ����?0�T�~�������1��˧�m�I^;0ԻBt�Zo���Qjy� ���;h�W2	�n�/ct�PI!��=�����bF���?�F ݘ�p0K��g�q�|}I?�,��D�����T��'=�R�1����ʓ�Ԭ�OUX�֪�d�EhpHz䮎�U1JZx��Wz��ʐ���ґ*ń�����ŵ6j�q7}r;F��/(�Ϥ����ga��h�nc����gʩf��uڀT�+�D�h���I���#��������}��vb\�ݒf�%	�+T�
k��(G���
�㟌<.�(�^M� ��(�w��ф.���/�
�D%+���I�-�����ojc�;�a�%o�^�N̬��w"V���TZ��P�Әo͗zlO��>�l�C�2M	�VT^� ��_�n�T�<���%��+Kl#�n��4Xi��qf�i���>C��5�;cw�r��!J#��ly2=����]·��س�{2�J�O�1�*煛tcJ:u�S����'���q3�i�� �~�aS#Hu��,�\L����(�֤v���g�R��l�x���r��#]����k^|���$����C�V�y9�gZ��m���c�������6N
��|��rj	>"��r��񣦒k(5B��_[��� �p7��������a���;S4����`4�� �Gp����I�[�h�`7+����DDނH������֚�c`��p�	eDrPJ���wC�i��m�R�P'��G֗"����`�Wo�s����	d�����=��,&���7�(���0jP�>s�U�ۿ_\c O�-`��R���M�DL��rppIM1�M��s���y���ܑ�5�ǿ~���n��SC"6k������+��H�':�������G�FGg��@��i���q^t�3A_f����b�65'��M|�&��ѰY��ğ4q�MQ�.�`_�:��!�s O�-��U�w�����	0B8f�ϵ��.md.@���%��A!wQ �[�B�������O@�K�=�Z�"t�̢է����1���n{�;4�G[�
�����]��Ѷ8���G�!\UtU=?�_�!����W�J�af��>Nb�JWjaL��dB��҅�LYO�L��|H�K��+m)�K�2)n�Ő+ ㋀�����h�\�#�-�`��c��V��B�!e�J�υ���Գ["@��ئ0�9v���Z9a�=��Փ~tH���)���	�m���#0�N
���V5�pz�����V��1
��A-�� �"w1�4�?_�Ԥ���O���ˡ�HE����B��@��'؁`u9F��BB��wlz��ҳ���Aի��L���#� ��'(S,�iW�a���ΑM5�����K�Aٌ�?(���$+�"ӕ>v�ئ���.}�SH�4���E��ӥ����v�]w��p*F\0¶[o��_�@'_ye�~v�Y���ʍ����[�l<l@<�����TS�i|`Q��������Ț$�u���0'��N�
f����i�@	:�G�8�()�Z3�>	��<;k��}EF�'��]ۖ9��\h(/��%	�+��m_	���|O�(գ���s��-�����=F�XRwPъ���F�J8���-��Ŷ���'g���c�cR1RJ�X]��yFO����}T��|#��gi��w��O��g����?磟�����Ӯ��5�֪Il�B3���0�D��a+���SI��E
��x�O�1�MET*2��KC��:��9@�]��sd����	<c(�a�xU�`5Sy���`�Ȣ쪈]ю�l�_�I'��4�h���&��d�����g��u7����Q*:�D6O�MJ�5|�s<��E������52п�4h���
��m��˧=�����#�b�]Č��
)�Ά6�X�����
�DQ�M�!��S��Δ�B�1��l���c�+4�6��dL��9�U83���'0�t�9r��~1ɽAyх��u������<I?Nc����`�F1d�NC/X�՚ᗜ��LJȮ��?�]1��S~�,��Z���l��������L*q�+�u�;�=ÛW�D�����s����U��9�C\<����co�6w�Hu�����p��}K�Y�|1m���]@�;!�lֹ��ޅ�N2�m�F8����7Nf��a�پ��!ir���A��`{���  :`����O%z	�l���%��s!�}�&k��ֹ}c<U5L���\t��j���W��d[�Uz�c���_	�A�#������]�
�!-�x�p�>1��.ɓ�Ӷ��-��^��/�UyMj�mFUD��Ц^c ;�тEEX߷&��!J3��߻=,B"b��aPEʄG��R2)���4�M�LRa�K�J,'�qEg\a�hϬ|#�1D}R�JU.f�"�o�X�-E4���7NKcFk�r.=�[�����j�G"�����)9Dl�N���`��xg2���<����2���9e���,��|����*	����l����`���?��Be����)����9��}xa���m#���(�X�2�|���J­�w8����8.��B'�G9��+	�}���A�}K�3�C|w#@����:�g��A"�i�̸l�8����Oh�����i�����P/Ћ���)u�DE<LaT	l�(BQ�L�?a!�޸1�fzt�8��#��I�Ojӻ�6���f��E�&�w�ZԎ�&ۀ�zQ�z/��h-�B'E��a��.�͝��f~�_{���Yg�Œ�V,�KY�����C����E{#�e�8�K̆�wR�]�dKh{4���+�l����?#�L<�B�/o��Bn����U�%���'�Y�8���.�l蝐���j�e���f:|�(	76?��z���Q�m\���݋�RT����uQ��hLa�~�pq2����im(U��k7��LT��0_>Gt��8^��sH�Q2ى��Ú�ւ����)~�֋R�t�O�	Tf��_|�V��]�E��|�_k�ɭqn���`S\OG����\���+
{��2P+�C�7���J�K]�9�u��I�
W�=��5�P\�⟃?��J�q�՝�OG�;�m�!db��E���z��n�KZ�O��r�)wrg�ٿ�"�?e�o�����{��c����LF8~���vE�^��Wu\�&�Y�fM(����\���7���_�X��5��_�WO�*|8����f��G���{Z���:$�lp̙.t���6����8����k�A��!�c<2� Kz����w?� �@S����5�� ��.]�.끖1�]|���ts��V�[���^}�9����t��תE��Y%⧐����w��iQ�����)U�F��H8f�	��,��2
�ϩ�Y#W�{��#.�.p.(H��)~�z��1|��@�����T]����
D��x
8��>^�:���sJ�����9�,��/��IlByD{��od��&�aGC�����"�緙�~��Kd�X8��%��] ����b��o��?YI��^��a�J1�
�����+�����m�� W�7�ݪ�J}���<���ΩjĪ�WR�x��������]��u~�T�ӗ��]��$�qG��qLv+��|���u�r�-@;hZ��L�	��n�V�� �����jyБ&����fFU��pyC���U�}����������_,�{��Q��s͙��/`䦳����9j�X�3}\�k�|����=���73'_IT�����]{�L"r��O��׈��&,a*9/с1$`�Ny����+�w�- [������*D�ԙ�.$bcN��� =>�:�zZ$���`�vų����u�p����4@SU��eCӣ��J`R;x|͉Y!�sZ2�q<�����7PNt�Mh찦I���ӬO@�-�2{����7������t� �JҢ_�T8TU=��"6��IzA��.n�Yv�6���e X�~|T) (ɗ�vo�Yv��Du��Ц����j��	��9+z�;Ԝ<�k�.���>_Ƭ?���	k"�i�=��i�2-�>'t}�g=�+
İ=5���L	�K$&�M�@ojtIΉdd�t�n�����b��P&�����8�j6��B4|�A���d=pC4s��$T�*Ac�0�oŰ�O���d�fG6{��]�j҅�e[a(I�g�;���V��*(iƝ=��������؁���*��ʴ�c@$&_�>�,�+Ϣ�~Z��v_`�r�]�[��j����䅰��3���Ѽ�`�FD��O�g�No�qE����+�_��C<�1:6���� �b�J�����e�+�!���[MLఒs����d=�#p⾨��!s�aBn��#���w�ɻ�3���R��{#���>��ևTIٴ񳘠��T��zB>�Ć_��nߓm�u�G�S�\�������[E�!�uނ���d�x�h�R<h�"̓戎�L�mD����F��&4��֠� ����G@hTezuP���Pp yO�{�k�����6	�!�Qd���*���Ԋ4�.��˘u��:��r�T>��N�+�3Oė�B�ߤ�?��*��õ��`��M�Y�Za�L��K�����m��)��ˈ޿1��y��
X�'���Pr�����0��O,`^���\����}���J8�P3��ǥ���53Q�A�����%e�cuc:��ykt�J�,
#�]"�+�GA��\~��7�
��G�{��P���R��+��:�}ﵤ���dR|?�Ѡ,b�"T�{K�9��/o�/�(L���u�+�DHї Qe�	��p�rz����j�0D@K�u�I2^F��MS�7v�/#Yeӷ �{ ɵC^�\�C;x�%�<mR�x��sF8�F?�W�����:^y��6���ȭ]�ڡ��ю?P�M=5����J8���Ŋ�Z��n�t�����������~�q*2g"O�qJ'�+�ĳ�xj܆J�.l�/����T�E:� (���e��&<�Nm��a�"؛��v����Y�^���"e���H���F��H��Jmu(�P'cP�b�;�d��S ���ޭ�<�����ug,z��lH���W�2�Ö�������N�S��t1�$�4�
m�|�V�s�M/��%�Z9�W��UNYt��Kq�̇Lŀ*)�df�4�������nzZ���0$�/��?gWs	G�
#ʵ�2�1ʵ"�!���`�l/�����M=w�9OKւo9�؎N?~���}!��M�#(�5���CpL��tX9��GED�n�\��yF,΃h�X��">� AL��
�8�21��Y������q@�Z�X�ͼo2���)g'�P@����rEe3��u,X�,��'�/{Q�#e%ܓ
�r��9��{*��*^��\���tj��U��n��D�D!: 8r�)�&��}����k���h2d��fR"֏Z&W �V�\�T�[��A�� �!�8�.t���	�B����u����o9�d�<����:������z ��؃���b��|��Ŷv���8Mn9iь�e���Ӥ?S��7v�K�����''L���>X����&�vb��8�^�u�]�ì�	3�G$ڵ��x��o1P] >�WX���7���f0�!� -O7�N7ƫ��OES�&�ƻ'��F=�����r T��y,�"@~�r����썛ڿ<8�nl��NC��g�.�A�*ZfL����3��y
sa�c��˗$���a�~	~2�RV?�Yg���w�6�µ:�x166��jB���_\�d���DS��Ԣ%�������n��R;�>ʫXl֙+(����В[R�1���"1}�����U��V��4) �/�r*|��>O;��2c5M�B�|�4�& �G��"�PZ#͂d��S��`F誙]������){1��~\�����]�@�n"h ��
σ��z�t��{��s�&���`�\��F ��4��K��,�m�W�[�£�d�H�.�t�#�[��چ
(J���U>�Y�|���U#�É��=� �a黑^Yهb:)���#_��6�6�Iȕ~�@���-RM��F_���Ȑ�H���,����3��n6�Հ��m-f���Mp�{9��u�J7�f�\Y\ә#���Ӈ�;)C��N �pP�m��<Fɑ��p<��S{3C@]����yQ������W�e(>KMq�q�'p��5j1< ���Ý���۰�G��Ei�I�)H#� �XQ��	k����q?�ؖ���S��#�Ng��Z�#�w��uU�x��]X�^��.��:�����j_�G��'�x�,^�'�=7����2-Y����=XB���;c}DW�V����b�>f؞��e�[X�ԽVQ���x��vp���SH�R4��d�r���>-_iO��<�F��do	z�<-��t1���ܨېY#]�r�αl`-��9)�FN��^JR�$�{�W>E�mF�x�F���t�:q<�4��w;>�33뗭x��"���*�*m�8�5��q��U�UP�h0[�B4y:hR�#ꆲZw'��s�v 0���X��VH/�6�(���yɸ"oec`��S�X�Uְ{��.CGaf��p�Rw~+igx�V���Z�{�M��>)�Fz��w��C}�,v�b)A�w9���8��`��DAҩv�٪��]R �;�l��ێ��$�Zi*���~�VBӸ��tr\駣�}t����	��=���q�.�J^���t�Y?Q:�Է�O��Hvƛ�>M~38�F�&魞� �*��/�(R#�r��ܱ�1�C�����j9 lQ��$�X#G��x���0O�,ӰZ�4~�-���.��%�g��ޛ<ܲN����f!{�xf��=	�����Qpb���>D�6w5a��P8"����Vڎa��k=�2�Ԩ�?��RRU��*�[�`�"�S��`��#T���	�ؑfLp�'I��[I�v6��	����	��Lo�������7@��7�b�8�L�'�U&���7��+h�)5K�C9j�{D^��/��f��ကx�k�b؅�m�p`��
�{a^��w�?6��n�x�[�n��ī�\�ji�n�'o��5���9.v��s/��b/̖$�Z$l�BP�V�;O�~
*���t,?��%�"��p*Xѡ0��O7��F�"����7.�}�Z�c��~Ϩ&᳄���Nv���~4s��&b�n=�g*7@��x��rR�w��*���뢄���U��R����ά�T)�Ƒ%�ư�҃�M�ٳ�b1&_����s���\�!��w暨[4�xPh�-(z��;S�*�.��b�/����.�>��+��XܳM ���/Eyh��bSN�fb�k
^�Tų����QO�*�%�#��X�a�@���v>�+{��
�iOr	_5�!���4S��EL�lj�շq���{�����ɶ��ߓ;1T��L���]Zl%	\�[�a��U����A�1���x����D����vO*ΐ�E���DgO0��"�h�Q:XN��D7��$}�~�ծJ��K
�;Ri����U�k?�>9ɐL�)��^uR�!T�c�AE�1dy<�\h�����jn�ߵ�!�#���6Zv�ɝos����oC�%�����rw���Y�\�.w(���v�x�>hz�����5J"�x�Q����,㹪+=k1�с74����yf��0]����kO\r8����f�8�}���� ��
f׏��}X�{�`���`�i4/#���L���m�D(�\Ŵ ;�ZHq?L�B/5�[�������h	��*�����5	���.���@�����.��>mb����$�M��������m��\a��HhuA���,�@w�-�����{�#��o`�B�d_����趗����hK������jx���N��0:���������t3��XY��}.�[~���ɏ{{i�gƁ|���F �lO�(���H��"�����=��J��d�Џ�L\��Y>
#�C������	�EB��n{�f8���?nQF=�`m]O�}-qgpd܋L��S���*�)H��q��L���j1՚Bg����:=������.i	i�7ܵ��l=dEdX�m�כZ���$n�)q��Ź�,uB�]�J�B%��d��e�0������=J��5�ۃ��!� ��Q,�b���+y���| $RC���v}ʓ@�rQ�IRY���N��cׇ���Ax}̷�7
��A9*���jL3m��tϖf>02	`ӂO�~��1��$��>Kj)x'���H"���łrXr H/x$��:%��W���8ɗ����|��{ �<ĵ����E�}�����8��P���
��X`'�^�t1G�L�F�<j���V3
�Ky@Dup��1[��el���ŧdd0l$ؐyO��	��ß*%��T6�g/�H�D�^W��C�vQ�����f���kv�(�����|�w?��ͩ+�6.�3����C�ë!�'wM�N�E����s��dފ����ZM(;MI���
RU5�<7��'�c���t����԰^&�9��4�>=�ҥ��.��Zh0c�:!>�'�v�犐e2�^�C�\�-��jB���r:������йɠW\�jbT���|�^ ̈́l�<d6��er�M!�����Gu?��1&��o�O<�͟!�=��X��T�������YU���ˑ�*nǂ{����9*N��/�wj�Ǻ��+�v~#�����5u���Fo���u��{��K�Y�kw�)u�P�k����Ƥ˨���P�� �p�^�I��<��ȥ�(�ƻN3b:�j��I��R�y���Z=���@�����������Ωp���C�6H;������	��6�Ac���0aO��p�0BOT�tŗ+����C�[L�Noy넾QҰ�췖�\Ŝ� 
�s��&�-v�ex �n�X���q�)���@8Я�#录��`��.�F�{C_�WU��>��i�82*�gCg�oN��O��hx�U&�p2��ѳ�)&�Ԙ42:�m�]P]0-7���]��]D~�΁��$[/�P�1bI��|�B����Z��+��O:�=hp��߃�.�!AR�E9t3��"�}U6ͥ���=X�zU��.�k�J}P<�q���/�5B�3��1���G���y���@����ٹ�z�^��l�'���^�0k�NgW�	���ʄ\������?��ZW��ԍ<-A��T�J�8�L���"�/� {���s0�̈̕`bp1��\ᱣ�ͳ{�*m����6Vڴ�x���9�����,�VTJ ��Q����` �:����tC��8��$��8�a"&K*IC�)�ĺ��K
Dl骽�bY�h��O}Q��.s�fH��z'�`�*i�>w��
�>��S�����<8�h���k(��Uҁ�&���?j�N��7�?�K���Gq,_g��)b�8��yY0X%k4����f�ŽM�'&w���Y�P�l%���		��y�3:)j��=�k�{�0�ҽg l������۪5��_�:�=���=�����T�a�Q�_�m���g�t
�>�0�F<8�H�'��,��X/St�� �ğ��vo���y���t��D&�7��W����i����H	��<���rt� �����7xM������`�O�I	W�.:K\܊��<�
��v�����;�o�ou��C7���OW�`�_�$����>]�X�.�3DO���#�p;�s�~�C�����\���c�t�u����|��H[��Y�����R�p.�j��#���j�n�ᶆJ�x����=$��G���͟;��jV(q�N[P�p�����eɮ���a��$IUBo>+�4����3���*�T�"_�P>e�;ϟ�_\��V�M�����P�|�����d������q�W�����1���*(��#����e�o��猗���=�!H2����҉�#I%'PB ��ĵ��V�����Z	�|���6�0��݈��}Ƽ�̓����<A;!a��|���?������!c9�dk�������ۮ-/��WuT@��:����B\!���|�yAK�ۭ�u�'	�����O�R�g&��5ݱ�@��Y{�w�Z��[���G�B��Ku�&/+�D\��b�N��B��D��͵������A���y�3���řtL�$`?��'E���P�-�%JM��<
 �h�ߡ{Er���&����5�?�u�Z�E��]��o5��Z��2g+�f����>5�-5Xח4�u����Z>�]���͍3����৵��YR�dXٽ��*0y-�t��]f�5�og��$�/�k��\}K��Rs��@b>�H�����.;"X8�e�����3p?ff@�-�줁��J�����w�ƛ��4�>���	�U(["<�� �R}����E���q1)������w:`���k{����0���`N�*���qe\��������"��8�A��2�����KC����,�pu�ϥ�w� �~�)yG�ܷ[�o�%�A�k�iH��; ��)�,��A��Y�F0�����j�f��Dib��J2����֗�!��J��o�X r}t�	�8,¼�����V�~R_X�w} ���ߩV���)�]���r]�r��x7������!�H�߫[�9h^�lK� ��V�� �
:*0�xJ�mob��je��)\!X�U^@�� PM��c�ݐ�P$$�
~�yGx38�����5�=	�i0@��a@4UK)?'��4�1;;{.g,��z5,�ψ�E�1���r�C;X�
M��`�m��n�dG!Djf�`�vT_�j�m�I�|�������=7Q��^���Q���Ub�6X2I��S����ɩl�df8���ϴ:�<��O|��YEZ*�0�g�"��{�8�g_a���	җ�sR�/u����Ƙ�Z_"���c���L	 �Om7R�����@T����,0	(���=�ϣrx.Cy�-��b��Q��a�1~���A�����tj��&�@�V��Z+P<	�zN��E8�N������K-A�DM�����V�%��e~R�mLQ��O�c7�d���~�*8��,���(�$@���v���'{a����,(8m���v\r���0ƀD�tP#ֈX/��n��^���zκ�zbz�6G���Pvz ʳ����1�З���IOfm�
�)1?�z�imY���R/<�X���DuN`