��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�L��58b�Y��u��	>e3gB�8��![�����1I~"�
7�@�@��;�/Z.	��u�w� R��b窫ٰh���%G(������:ul��&I���|��DZ�#z�Y�^Fk�@$)`!1��.t���^���*_�'3.�'�I�ߋ��Y�*�p&Q6�^N��Xw+V�H�և%���C~�(���+ػ��Y���&Uש�F�gմ�ِ+-%���(\`�����q�FM[u:K*��qDS�*�[B;s԰I�1�AݙE��.�w�d�ñsA����Uw1$�
3n���

.�?4����%}S���*����9����J� }K����KZ�;f��S�m�4dw��E+��g.C1��ڎ��s��`��J�F� �cՒ���ͫ�3��L���^ ���d�m�ʞ��b Y�g=o�
�!4���֑rH�{A�I��i�@z�F�&��*����+�� �'.���H\$��ũgn�_M?[�sy0C�A<K�&��	��U%�l�)�(�<��F�V���oƒ�ø�=� ݜDq�� ��?��z�Ã~0�f'����;/�1uov����G�2RL*�^mmq���Z��8��)��Bd�<ѥ�K���F���?ǁ��`���BTNW!�Ƞ�k�U�\yD ����b��T���+��+L����~���'�@� �01������3Rv�K�zG~���B<�#S����9�`t-- �w��,�J9��W���\�{���^��=!˙	xb�I"hx���u=�����>�ّS+�s�(�������K��V!����u'~*F�'��Tp�V5�A�r׫����UkZPcy80�@Z*��O���B��5�s�ʦj�+�iF"�X����rW�p���$�p��ai;҉E,У�'�R.5��'����ș]�!�w]���c�d-O�1of�����M�e[��]���WJ(�,L��3�:����D��50(.�z��h�7�&$q󐒰4�9T���-�;¾�6Ɨy�dD� �F��J@\1�j����1�~_�؄,�`��t��D�Z�eZ�y<�ط��;���~���|�*�>����!��E���@x���|>*z��T���f��CdAJ��U� ���L�'ܹosP+�b�c�bn���n{�
�;1��bQ&�.��/5�����P����Q|Rᣫ��oB�{��t����qg+][��_����>O':w3!����]���4Q�m�w��+�,e�d~�|;,��@��`މ��G�Xr������	��
b����Z�-���N���͓���?���]:�tE9:���H� ��)(Ш��4张��L=V�#�y/�*�K����04��žja���x�ۜ~]���ՙ�T�����`���0�iѕ�r��H��z ����[ 3F:�SP�R߂���Tؾ�Ċ����0����Q(}��PT��5(�{'�j?)�%2d!�����O�����,+)haS&�P�����
@AU�O��S���$d��7K��05u���JN��V��T�jWYJ�nn�.V�昽T�FCO{\֪
���(4��?�`����j=�@�x��Kv	V�D	�dD�P;���(U ,`��e������v�t��tK���������C
*`��$}�"Ի��C?B�E�0|�Q��nMD�i�d���Xs�+u����w�Ux�>� 1U��H��Q���:�;��*�`�1�BW�A�h�ў~��+X"���>K���; ���Adc8�q�3wh-Mj�;#<�'��f�W-�HƓb�+��4����_죠�MΒi�m6�;f�(8���/����	��]�(#ڌ�j������#�7��
�g�1t?�Cƙ�~�M�L��ɒ&�ȓ�FKAc���D�I���Љ�9�3X�?e����uZb�D��mɉ�3O�f��ϙc O�@�~��W)�4�K�m{Jy��җ	ӯ:�m�VF�[f����j�s`5�z�ƞJ�<�ۡ���o��?�ħ�h��Ua��V��B����d$�1�j�ӐK>u	~f�6�8���;D"�q�qC�.��	����X��HO��Q�)��9ш�N�"���xx!5������'>̦)�7�c橐d�kts��@����y����0�L������I<}������%����(�|	1H�g[�n?�I�A��XګK��gԅ��/�P	�g������B�f�<n~�i`���/�A�Iԯ��7���JKM�u(�8#�:�[~[+ Q��?9��O��O��'����*߲ԥ����N��҃��;c���^,2�%\=K5�Y!�����u�a�}��$��2?6)v	�{�*��4$߀N1bk=����BZ`��_�7M���]3	�F�D�8t�8����E����k��F�=?�o5˘�ݭg��g�*V�a��Pu2��c������#زvV��K��	<����e"�v��ok��BF�4��%��p[��|�0)�iR��=�o�c��~{�`#%�N�w絶���D��蘾5�/d�������O|DuCzڴ�d���:��#:�*��G���X�j�1��0Bq�C��3xbF�:�BK˄��M�F���%�с��	�
Y���X+���h�<��2�k'Q��1���޿��\^.bI
��B:�r�E`5 20�F���`�h�~�f�J)AyJ����z�Q8��^Y���h<o8�4��J�i�zu���k^�0Ax8�r�n�$�����>?7��=p�^;���u���c�Xi�eIx���R��P39��{���_����#&�&KQ�ѓ�-�\���k#B�s��J��l������h�D�Ǜd���voçri+������:���S�^�~��y-���'e/{��O�%�H� �?�����@k��F���p�k�C�s]#b�t����xu���g񴔳�~�Ij�p��7]̝7FE���zX�i���	GTV�k}E�ՓL��:���^wF�����8wMQCE�3�	+�@�/~;��ĭU1W��u�T���!?ޭ��ށ���h������{��b%�;�_ba��cB\�ܡ,}�Xo���3Æ��#&q\i��u[1`�������׀��N�PY�BM?���J;Z&����U�ׇ�(z�p�Z�69�⨚�w$e'�5A��]s����i���n6`@@/C����$�����&����Nuq�s�\�;�-.GKC�lˆ��1[b�f��y<_�Q�}���Ѕ��۰{����l�(�5\�L��b9@i��LR]�F��8�m9�I�wm=�3����v�k9�=Hq\A�
O�醆��!��F��7��7�|��
��ncB!��l