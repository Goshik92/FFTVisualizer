��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn���\,�Q��Z��N�S��k�OdQVl���Y���;*H�H�B%�1�RM&E뺍��X���6��K���L�:����C��r_5e��:m�7a�]8ܸ��i4��2hp��Xd��]�961a_5��K�1B���uX��	���S�|���^o[��d�'����۰��@�����*�)� Q6e]i����ڜ�"��ͼ�b�m�Y�vմ��'{�N����\S�e��%N�¤x��U+�����M�d��ݿa��:����lt���8zL��}�Ɣ�S��
 ���w�zّ����P�3�}��~�n�f/1�3��:�hnS�C$Z��˕(���S��o��Z������UrȐ�ʘ��c*��\���9�+{.Ꭽ�C^���X�ƺ]وқE��z.�8q0�p�K-�~Vڳu�J7ŕ��]m[����=Fd��d���^G��&ҍ���=�+���Z8U]��İ$�����hٕ*���Y�/���S��u�ݻ[�7>��[S�Pu�=s؇���S]�|GT|f>{z?�)�A�M9���E}pلG�^�OV��(p��D&�ǣ��J�#.,@r	�k�م�l�� ��$G�ݔ	���sRN�!��(��!:44�la)��e�Etp��m�sD�C����<YSu�4S:osw�|k�𶓄�j����*|���ͭn�8t��3D���^�t�+�����Jp��"?�V����Z+�O.UfoZ@�zTNɈ���S*�RSc�砖S�K�8.
\���G*ǐk+k9���rf�������a[�o9�)����ّ�5���<X-;��ި�FLL��1�%�,D6!%H��������^��u��d]��@���5}`
����lbv�m4VZq�|�f.��Ŧ��� ��ƏQ2/?�/�,���ou�?)�J-�-I�"h�7ڈ��yCqn�M�R4�����߼�y?�_���l����ݟrm3'�[������p�z���$�.<,<ʥtCd�E���Rg�a�����r��6X�Ϝ�8
k��K�*��u��	��_y��v�򠇺<�mI�M8�v��k�<�jq��efI��/硌/+�)~��l�o����
�#l��۬G��M��WDv�{���Ĥ�ed�����i> �'�5�-������+߻�.V�y��?�uz� ��h��ڱ��Z&|� V<�U_�Z�|��c��$f�c,W�>�@���W�s�>4�-9H#�dT�w�i��js���h����1(�:7��p)�A��*����	�������lA�b@X�O��J=�zadJMč��}���Z]���P�3�~�^� ��uv�|F�v��]lG����[{.��p'�֢��wZ���Ĳ%_�-G�V���.�4>�
JT��Dl�����/���'଍7>������uBsH5:N�z�������0�f�n��o���B�b�v��bD��C��e#�yC�:l�3��0�F���W�9�6/�y����k6xfj@����P���]�Ė�=;��~����O��qG�@b*�u�E��n�:���֒}�??Z��MZQwaQ�;�O��-�3��g�B>�&V�ݥY[��2��J���˷�7t �=��<0N��:Cg�]�W�45t�iû���hb���L�����!�a'����3�z
�zK1�Pu��M�W*�������1���m�tX
pi.�|��x��e�n�����(k+E��0�Ӹ��������O<����~��|��_�e�@nbK�>ʳ>-)]�[��I|ڃ��������ok�Ty#T'���/�Q�<���	��q��k���2��Ak��g.S�c�a�袖��#��j�>W���YYn#��HI$pt��y�(ib��+ĘL�7J%:���{~]�"[�����&|�`�� 
�=yM�1K��II��_)m�W�6Y� ������ 2F*�̈́P��a�_�c����ᄜA�}�
�^��-vmd�']�WGX�W��D{����E��j���L��B��7ǦtD,�Ch�o�b�WJ!l���P��tiZ�p}�4�^8C�A�t�Óp�Ng�(�%me�+�UN��3�/�S�Y�uw�W��;d��Tk����ّ�,I�GyY֒�H�@̶�{�Yگ�Aí�b��(
��������,��L-��-h�p�����޿Ԟ��T���s����P�}�tO�W�[*M>�9���������h�ۦ}Y�q���A�����Ęj�k��]�R�#��}��̃�h�?�i���?�H�ž�5���_`LY��<��K{�*�3�=ecPY0w.9��[{)�$��'�+�ޕ���>���aD�Q��=g�>kãL�J$�C]X��	4V�-��Z'�N��*"2rE-ם����-��:ゃ[=!�b���ܧ �exe�R����6a{/E�D`���3`��J}*��%�d��I2��nP*�vc�m�6�z�V���89a×��*h��b�`��">K�2o�.z�{�2�����&�(1k
G �X ����k�~�h�Ę�[v�1�l+�{�/���N�:
�8{R�o	��)/}���J8>7��'s��e)�*�~)�g�R�):u�Ɏ��F�t�}���/���Iv$ηG����0XRJG�Y���(ܖN2e��Kڸs�jw�����n���)y儋Z'MӞ��54��,���3]sj��sT�)�ώn}��wD-H� t1��u�X���C�dS`����`�l�W�N$��	��u:�Jb���F�e�,5P	F\X_�X:q�bdG?�p���B[m]	��A!k��.���v���3FG�?.��(����mV!�;,F�+s�[�Z������̧=����a��2P--�a��bW������$2���cb��m�D.1�KP�����h�#rܝ��PǺ��� \�g��_ mSG�ʓ>g9T���+h�H�L�׹��{�2`"�U���^pzzN O���jY$k˅#��Ԣ���z�wq1��T�n��<ⴄ�DA�C��O�Ļ{�Q~:Z��^�B�N׷����w?ņZՅ�m�)=��W6O�R��]�u�5s})wŗ�&	��j<�����G$15d�v���g)K�?Q�f�q��͂"����'BEc�~�w�`�[یˮ��ι�"��6����&	��)�ڸQ<� �g-l����p��T�K���1����x�")��/��'4JU���Oc�fE�����Bs������5&�Bk��??��}f]U�(��ѩݲ�w;�>5�,��^&�V
�Oj�:p���ݙ%�L�!�?�Z2�Aj燈��%/���\��Ȑ4)�Il�#3�W�����R�hK��^4��7�Uc�t�/5P<�!b��T}��F0�9E����y��A��]}ĸ��0��EI�p*����q��PFa���L&-��� !&P��5�K�?1Wg)���y �]�d-� ��1�/o��<��r���^�iI�ao�z�֮�.���n��é^]�wR�2�ంD|�0w���LrC�CS̜��A*�אѠ�|�H�m�4�Cɿ��[�jᤍR��/<�a��C_�Ħ�"G��Tݑ�~+<�-���+��
J����)�bS���m�X�+,/ȶɕI�%ʹ��+,-Ɖ1v��T� qDȀo(���I�|8��?.lX^����I�o��P��)������V���$��� 9�ќ���'t8�G�k����7�īXEK�������Q���ݧ��Go0�f0���2tɌ�e�6Mp_X:�<�y�!��=�e����)�<tlhgGh����)+N���yF��g�\氰zCO>���9e���y�����qfL	/CGx�Q�I��WH+$f!��?|�}�a�s�9 �O	�B�|\-������K��	�|���EĘ`6W�Čpt}~���>;�G	�uO`4��}.k�7h�D���4�����h�_�A�Y��S�e��ewr��D4��UO�~�Jyu�2bH<� 8��>��ɘ[����*�JJ�+ݗT������g��87�o�{k�a�=�z�\���/���l]O���}�nT9k�"�w�6�[����M����v�K>χ�#��C.�0�UA}����t.I���#����^S4޹���x��V-�1����A�0�9p"�d�b����o�>;���4��OfAq}��m��C���%�a"�Uaj�}0�?(U����]����,��g��b)��l몬�ô�B��!ZB��-}�mT�c��S�@R���Nݵ�5���q���rI�����۾�@��� �,�«�';*{R�2��Q��ߒ���fx��Awؔ��3?�_k�o����А	��1K�\8�{m���&��A���h@@�m9���rM���v+����U\�| ��B�}����ڴ7��<o#5o�>���M�MaB�1�������k�t�M����^5N}zG� ��I'l�j����W�A(L-�����bX
���9W������C���3�o�� |Z{iJ��΁��̮�5�U����w �Q�x�u�j8Jr͊�_=�n���R=`j[����H��<�4)��,���2�t�Y� u;Z��;.'�hM�Q��כ	��Ƅ��hֻ����4?:n?���b��t����ڠ^*�k�����_h>���@p�_mƽ���S<Ol�^�4�B��A9R1�cޫ�KZ�g�۳T�A��X�~�"��m�zO�mS��B���v�܉RAoL����w�r /R^?���/{Y/�5�)l��
`���S�E�Ļ��$&��?�C))��v�C�����!m�%ӡ�?,���*��!=*��_E-v�����^��(+"�f�n*�݀J�<Ih�,�{&ѵ2	��u��.�Ꝯn'�E�2|�\��r/���Aߢ�;<8P����TXОFvNiK.������*Ϲ4�ps�t3���f���P5��c��/����rs������7ۏve��ɓ���F�4Q���ƒ]�/\:�̧��
 �$o���[rl��=�]1E�O0�5���?�dTE�3�ؠ��>ʔ����m�'�nP?��?�L*Q|\���p�굶A��בo������&Y����ꎟ�������h�y#a���MI�wfP
]عB�H|���;or����t��̙� �?z�>��礍�=L����ov�Z:�6�;rJ4G#|>��9���+�y}�O���N��8%����h�;xS�S�l�@e��2'<&	Q���7����D�=,�;,���Z8��O��$��Ϣ��W*��Vj��ǉt�m&M�"�G�M{r����[9��{�\��U��<_��'�
����a�`�����v{n\~��C�x�AűX�eg�	���<�Q��ߴ1y[䞐Jpz>p�d��?�U�|��'�~�79�a�D*�Dj�[��0D�Q��k\�n9hȺ_�A�DIINe� l�p�@у\&5?�����
�����T�9x'��z'^��>77#pI�θ&xh':�;�ZGD?�+�!��^�b�Wq��}
s��Q7� !�P�bt;	�ҋ��%|����~]%�Ȼ�T�������n��������L��@Q�:��V9�"��9,�=���J\��Py���T�����һ�K��@�FYo_�ѯ	^�9��|&_�����A��D�L���p�/�󺩏��''�)��9��[ʺ�4��A&[	̗,�*�.�W�1q?$A��,�Vmt�¹����Z@y	�4<N��­���W�D%�l���ӱ�9�<J@�}Pb�b^I�U�!9��=��R�c�H�.��!Z�Q?P��f~/�U�ݱ$�aa�4^jo�G(p������`,�q�F����,��x�!q��?�]Z���b���m*%|.���B
[\����P~J݂��)��b��j�����J�>���n-���iP`� ��7�]H����qR���+@�E�l�͌�g�?V��	U&������� 
��
��o�$�8�	g����ށ��	�Y��t�������GRǇF��٠�#O����OR��sc�3��!�@�Fl����Y^��z�s����fO�0揰�@u`idS"�V�%0��z����C�����U���H�$#P���/jm]�b�����`l�M�4f���$�Ňk����Imm?�ז49�5#��9��R�<��6"`E�p1vj2��oN��:s�^S�#͑-�0�9Rh���A�Q��Ԕ����g޼ݶk��!�x��B�k�7������Z����鬕�tBQ
\b�M�N4�u^r���7��2�Ȯ�,���P'�Tm�m����+��Lԯ��Y��N�;�nprTZ����Ǌk�b��$]�"�!���@�Ci���7ԲI��S���)BwqI��8�鎻�
�g�e2l�QqDE!���J�Ue0�d��h�_𡜍.�ˋc�[��Udi$��[E`>�#%C-:�]��� �2rpQ?�Ȋ�"���e]����\�ံۆ�zHj���ٓ�6�n��x��DK[��5	N��M��d݌!nrTb���I=���  Y-n��ޗ%mЍ[9�����:�Ȥ��tDMϡ� x���s9�L:�K��pIM":o�������3	�	��e9$p�����W1iշa5���A	%��ǡ�1�D�4�e���tI��׃#PZ l{Jed�\��tS,&�g���c�a	ܺ�}g�.�|�kG_9�d,_5v�,P�g�k�-��Х�ѱ���f�S/��o�hs�@1���`,����sֲ�m��"f@b������v��i]YG#��*�������5�M�[��Ɛr\"�T�Þ����ȦI�L���I�ZX.ò�l��hI�j,���J7��o4ힽq�h��,|BȔ��`���Y�1�`��6�m�G���ƛ�Uh\�L��yS;a�������GPa� �C���U��9�J回�'<&\��q��?�zls��%�m���ќ�Š���.e���$H-���Q-'��2w��G1�<5��`��9B&Y�o����7.{{��!�N�Y~�D�1�QRd���.7��pF?��Hѱl5�s��E����Ͻ���Y����ޘ���� ~1Z3�� %�e��׻�
)�Q*1�-K���芁���������oP��V���#J0#�ۙw+~�7����M2Z��V2�H�[p�{��g�	<�&s�m�ծ@~H~7��y��_h�jew���~�4�Uw�Ě�ٓp�h���y����w%�ˍ�J�d�(�ӻ�fY��4�I,�=r���gb��£芸xW{�`���3��^�{��:E�F�w�I׵��q�վ̸G�H�z��QԲ��]�*�������	�����y�_%�rڭ�8M�~�c:vy������"r�[R����1�7_�He�1Fx��PO���G�����=�!�\GFM������^3� �d����N��4����G�{��.=���:�<J���Al����t=ٲ��*{���#e���Qm��j؀��h�ߐ�=��(�}���eY2�=��o�J���m�����N�d�<;�}�^y1%�@��[H�����0C�a�Q'�/�O�[E�3�r�'���|��O��I���c/i�P�*��LJ�EÁe3r�k�1�w)0��C����c]ڎ�Q��-��7�:�����<'}��2�)�K��w���c��^B��.�����L9!�v@^sq��!6���k654�p���5c�X/�n���{k���I"��I�N��=+�+�B�wk���2�Թ��:�e��0}O�J�6Y�}�ºj���b�D�u��V*�]�&^�D�[��g恋l�����9�"��(.-k��c�����Eh�I���s#0s�q�B��qD�3�kp���V�jЪDw����8`K��LO(C��� �ߗ�/_#�*��O�5�^(�]'l�Si�?�%�B�gE�]qa^6�]F�>�ڱ�mh�0��
�:�Wu�YW2��D�$��
����;gH�(;!��� �wA�Y/"����Il.��wjg�o9�
-��L�X�:�I-��vv	mD�R��d�S�'O��-|~�4JTA6T�O���*��P��[GwGw��
�g��Z�����攘���c��H���t��4/1�?���$����a��q�9�R����R!ڧ�����G8�n��H���8�/����!���X'v����>����Zm�M�<
#�$�Y]��N�#>�!���<W�b�npJ��OLHp�OT�i�6/�ܥQ�]s��d�o���P��ۼ���!_��G_Qv�e�S����Y(ؐF%�} �zq�Y��ҹ���������׍1�B��+KqT&zFX���B�A�th<�����%L*͕I�1q��J̞�ՙ6s����[��:-�Ӂ�f����`�I��1y�)�l !�Eλ<�i��wu��߅�%���=�hͦR3�	��՗uB�Q�4cK+L����5�g
���5h�\�\	_��Sœ�10�(xybG<ͺ֣�є�SX�����}"�F$�[��-mS�����@$�O=S� �%�4,0:�@�=��b��Xt�{��Y:�� �O�I�KP�}������n�:�X�),��,��M:��ώ�!C��o�v!�`�̯�ރ&t�*�m���$#6����W���ʧSjk�4W�_�6�U��ꑛ��	S��]|�0N�I���Gtd�>�̈u{�&(���V�|�r�6<g��g���?ガ��,΄r�h	��5R��Uq���ߜ�`ș�+Zߒ�P{�Cc!=4��%nU��g�ڭ5I��~�S�r��I��p4g9qE����*�JJJD����5a组�8���v�7��vЩ��[VuA�0�	�\K��I�L���f�ʊ����� �k���٦~=���4�Yf���^Hw��_��C�]j9��&��[0�����j���av�_R�����Pp�[�� 0�0��2���g�K2�𘟁l
�k�YQ��:+j�����v��Ч���A-"_��P�o�0����K<]"���u6Q������P����`3Fp��
߯�2�w���s@�;k \Y����6B�ӭ���ۓC�O�`�Qщ���>n�=��C��I��h2�<�f�P^�]�C�E���v��ހ�-��Z���_O0�'ND��,ؚ�:��@r(��eX���M���4c&_�m�;���x´���R�<QD�i�Z����624/N�Kv���*Z��%!_�G��p��u��:I�={r!ڢaIM���B<A�� �'�~"�Rw��o`[���\�I��P`��N^��QZ���|�b�c��C�@E�]�3�j�{��RV8aUڡӻd�X#�?�D�%҄�bpʯZ(�1ӷ��Ww*�E��)U50���oп��c/�Em�N���l�3�Z75���|�D��?)Á��5�R������;�A���l"��̯i�k'{�$G�K�y=���	�E� �j[�oAR _�N�*3���е.��[�eYu���v�F�I�M#t3�¸h��٬�C��j���8 ��R>_΋��>t�2!����&MS(�� &8�����h[���.��%�p�	R^���O�"��5�ؤ�s^M@�!ߪ�xJ�m��[�<+*�S1�j��n�Vmc����T��&ڴRj�� ������6:Z
k�7P�_V��3? �C��?�-�h��6�'����r`a�`Y3����p�[vZ�J�[��]�RR���z��'���I<}#W2���^D�1CgǨ��V�绬I������`�5T�8	�[��z.��N���y��=ō�iQP�`�.���Y����h!&��bG�b2Q#��:it�������D��>���N���T�c"����
4_h���AEn�A+�w}�Y�2�%񣚓�0�N�����%�Z���n���h���x�UuzC�fK�������ʔS5(vE�<�IV~C�����y�)\y��F$�
?�y�K���/� ��̵�y���=�3��96�U��K9�+��ƔX�\F[o�1��{��˼�(�1�G��`�B�|5�/"��xx�GbySK����l��M���؈Y�M�Bx��.��b$��M[E�hJ9�(l�]ؐS��)��L���mcni��Bu����ٖx��ߡ����'�pCb{�ť�pB���P��}�d!��e�C%�=�Y��dk\���Z{wl=������l9gd��P�m��zR����<D�����gd�
�|:�=} CO�k�e�ϝ
�b���K�8�\���4�R<(�4���ۀ�Y����+H.���v}#��h�G��oPGfm�͖�������l�� ��M�%J?��5�8$��	�?g��`!z�#e��4$�f��j�9�{t7\0*A`��K4����l@�1�OB������V#p0K��f��
�Q;o��*�{`�+�������z4x��'F
Fa�w'�)tlQa��y��a��`�'����>-��@7�o�"�n�W�^����^��K��=�x�a�f�U��8�K� ���q��k(E�9N����F�>ū�D�������$Ƭ��.G��x�[����M��<ݠt�C�9q[8�3�q!�+7>KF��C9�"� V��l*B;B^�p�H4^P,$�W�@	�H��]�m�y����]��hd���2Q���Qcn+��'���)��P�h n�7v�R��#z�2�ޝL$�2����-V�Lk*�����I�>5���.�5�J�T�-W��cMc�2U��lm�=�P�[n���@��w�_����j�C�+�u����4�-_��W{�h?^:�ܬ9η� }�4|4(Vf�{����iݒP������;�����ɥ4�����@��\;���Q�X��A�Q*��fԝ��l��ei��ř�	���m��be��?�����\�����b1ڂ��"� �G��H��$��= �e$,.	~�A5�{�{BZ:eɐ���=�6u��NA�p��Z���.�fW@`w�����!���z�~ߨ��J��Fn_9m"��y�@��s���+�!.�QCJ����t�*�+�Zx2��{�	:~
����<���-^�O��ϽB$�Z�mV_񠝪)1���`�]o�x]�à���Z"/�O���-Ku�~D���K�\��y��;wHr�Ї$ �<$�P� m.�������2W6f�L����w�٨��[�0d��ED�9�'H�~Ĥ::s�.���8����ZޭR�,LΒ	�Y��[�S��ǐ���F���Yh�?�\pȎ�yS�� �5����PQ�e{�=4�Tɛ4,p&�ƭpB�{�٤��ѡŹՙ��nY�o�E��a��VG���Ϭ����V7Nmzz:-�~����r���-A�������2��)#���X���~x�9}���7�dƣۙ��g^�\������$�r�1���qzr�t١@�g��0�s���!8|�8
6hՓ`q[�������}�R��i,�SvF:M�����e�uˑ�X����f��R���2`��}p��������iL4X��K������_��hj�H+׎#���I�Z�Es�s��h��^p���"Z��z���\�#.�ڀ�i�
����{�	��-�'"z&g@x'����qN������q\�/[���}��P�֊U���˷����R?�@�����V�
}B;�}�/0��h~��yL���G��DFz����RW�7%;��/���i�g ����i�I��r�-'�(X�pqɳ�� v-�B������|_Z2f̥�Y%����%%��cLg-��2j���<��y�G{��� ���Z�:����ZXAȱ�`3�a�����K /Z�j�A����+�����a�{+�IS��RB {k�e�[���đ�}�8NqGD�5# ��ȍ�B�V�/"�L��b�	�IG1<~#bB��s��<���ǋ�ŠK��_��w�4�_H>�u�`�	L"��2W�WkkW̿i��C�++��䡷�ߊZ�i�6��#q�}uRAᮥ
<�b�?��:(8���ކ^u�o#Cɐ���uq����5�6D�*W �oc��H��~�nP�s����P��3v�ȒR�!Y~��Ԉp�R�<����bV��{F�_�����>؇��Wmrx�����9ӿC�W�Vt�"��jK�2HN�#Q�9��&���th�𳶨Il�5����X�V���gEZ�I:�:�\F�����ev����ᬺf��$���Zؚ�z��ݨ�h	��j=���L�o@�m��@�M�E'�����>����n���}߱8����ol�Ԛz�ƹ��=�U�"�<�\��4��������h�:2=�W����:ײc"c��R{��
����:�t#x�z�4�	�%�/������FRgߗ�6pe��TH�=	�����Ure_�0��;��d6G\[�>9�����@�;�s���$����2�Cn��i���vB��w�ϯ�B�^����ct�u�{��1��0�=���3�xos�N!�!-
����U��z$/�7/��3u[����u�ˢ1P��Ћ�.�G�ݡ�P����`�J�Y����l�<[�ŭْ޿��"���(�lY9�)6�ق.�O��k6�f��-=.)��`���'�%Z�)<�WI�v�`-�#%f|��t�l��G|�qb ���@T.*L(���}�>�|�*�x,��	V*,��dq7� �x�Ik.���1���k����>�
��!�H���6��V�x�4�v�b�k@�6h�=SQ,ڶ�3�W���2K����eC��l�$�t��� =
��T�������Z�ェg̜9���X��N/���x���7롬tK�u"v�ɰU�2 D�ߜ��e���M��+�!t�?�*^�s������i��R
�(fl�&&.��)�P�����ټ]�D{M�;��� �7\�~VnNS�F�[ô��k����]������\��Q����,�5���>�F�b�����.�s0s/�_ѭ�Gb='=�`�7�p����Ԏ{)X��s�D�C�#q��F���~^��V�5H4u��νK������vx��R�w(�Yt�8� =�N��nK�SK�7~�����:��˸�n��Y�zEY��4j�:�ZUm��D���O5Mxb	87*G�jf�� F�S�!�+�8>�:�C7�5^U9@fo����l�4�RP���6��_��q��U.���� ��9�}��h�1/�i�@oX���,���\f��S��3��'��],"!ૡ<��$A譞��$r/oz����ġ�c^8��a�PX ���[��[������N���/(H�<��^k뷋3�p��\g'�[ƴ;@�mM�u��@�fl(u
u �M)킀��|*L1Pj,��t�2'>��qMӈg�j/R�Bw��3Vf�#H�v��舫}�pzk��h�(��*ߪS�M3q��,�c=���3��F��<؇N���w��f���W���c���9�����x㰉��X��`|Sv]&bm�T��T���1��W%�@�[Ç����9�YDV��ضz���ժ�����:ݹ|�T�+�K��D��:��Ю3ڪ��S%��豎d�6�,���#��o�@dY��m�.�,3w������?Iɵ<W��f+�V���,���m�3������z3�8i�B6��A8��i�
~W�������H��˻ *����
F}sx~�7��3���U�������lW�,��^/>�IKH��6d`���s?�:dY��	ک��[؅�[��l�O8����Vy�k��_�晋�T�� h<λ�,JY��T v�}�n?F D~z{enbok2P�I�;J��f�E��3W}���d�(����5���#���5x�^�<N,E!%>����/w���$�>�����~����Bs���g$ݺ��{��H��|.�a@N>������2�Ez����R7��%��CFUR&-EY�d��*����ě��w*˴��P�+Va `��x��Q��΢��x1l:�)]���_`����_�1�wM��&z�o��4RL0�w��MS�䆴�D�'�(t2@�&�� �VD��_n�N��6
!O�S���%��%r
�w�hIk�l��P�p���Oz�aA��/�ֺ��;i���?+R�$Y�u��K!��PM��@eq7���]�hj�����
�B�l�.����5��I�`������<Y����\��Po�6���w1ϛ�e�~k-AMȟ�s��b(t�=��`��9I�|v�4��1�� a��SG.�b�n;ٴ�b~����sa"384<Ra��m�hy��j&8Ĩ�����fYa�n'!y"�P��i�??:�o�*��X�N1��ҧ��0�)țA�C��KX�����˺oe�B=޳�WٝC���l��i,A���k!�i*�쨴c���	�tn�l�˞X|������E���LY�k����l�5��{�J�Yc��+u)��Ǝ%</Ɵ�)WDb����w���BC� ��q��0�Ġ�&�D�C��܆16��FL�&��:��S�����ç��Ju@-UHg7�"9��L���1�w�K:=�S���q��wz?:Q�)�=p����d6�fkk���6���g,fX2!�ʬ�;�l�x�Ҳm�Ѷ���~p�[��"<#��Z6\��6=����0s��T��^&�j�Ay���,���t�E�p�w\�1���j�^�zV���v����I��3Gʪ��$�$ B����� ���6�C��1H�QIx�9�7�5��e��Z� 9�4��k�j^?�_��ߔ��x��<g�����a�s��"��Φϡϭ~awʕ�}��ROX�kN�������\ԢֹMzz�8>xg[fꍛz�W[����!��P;��Gl�*�С�n	/}�}&[��<N@n��+L��aL�ba�V>桄�S߇G�m�0^���-�ⰷ� �:����L�!�Xa��y���P1���ݴ��2I��%�_ۓ�Ԩ��9��f4��^I�6�)w��dI��r�(�CQ�s6'(=ӫ��t���bj�Ut�(��]d�Q�YLD��f�@�!� vjx�&��z`�{���" �aq�Ԟ?@,i�'"0o�7o�O�΢���W�)ʴO�
u�=�͍z7W���·ʐ��ED���T�z��F�?�N0��Q��`�˼s)!9�Bw�/C�A�Y6��~�f���9���,��G�в��1sjhv�	*�'@ԅ�[�)8�얌(c!��k�QM=I@�����H��v����8��!��è'B�?=N[�۟�\���67��cRә�븠�t����`l�
�I����T�X�������-��n|���EK+����M+��&�6����3+*6�%��)�L�-&�|�*�|��y��C���N�{
L�L-������-w�i-}ti���q>�Z����w%=Y�N��J�A� ��I�5�Y�	�Dʭ��뉳-g:AL��C(��Zg2O�B��-��� ��z�{�w���ܼ]&:����՗P����^��wQ*:1��US+`:��ǅ��.���z0s�8pE$�hs���dǟKR�)��4\����dk#���b�v��A[ɫ�^Xa %�}F�^��"�ui�¬�񘾡���Ы�I�쾘c�h�zmx!(�-V&|���_G�*Jr�U�M� �����Z�`�"d�3�����>��O\���C~����z�UG0U�x���6�}�y����B""{��nՓ�z�fq{c��1�����Xez,!v��$>D�it�h�홊VhĆ!���z4�P�,;�aQ˽��e����M�'�>w�����Mg���BȲ����h3�����'_�(�6 26Tđ�G�Z=d�=-c���T�,WqQ���h�0?wѮ���J��`of�yh�z�� 0"�.�Fs^�@�ãr��/ {�����к-슇s޷�?����h��'�I1%h5��W\�uq��0Hm�PH�n�f�/'�dբ�*��ِ�Q[ט�W��K����esSc5�kM��--�����>�A7������.��T�~{��&�i��Kk�;��O �ʭ�mn�`9FB 0٬��4m�s;(
WGK+�P���+V��[g5<P3}Ch��O�_mD����l�L��HG6r����W�u+׾'�,4�����7����jRv|nKБQx-�Տ	�,ܠ��b�^ ��ZV����f���HnA<V�V
2�`����]/�v&�CMY�(D���� �[��}��D�4�_d/[�WNܝ�X�!�>�0��b�=w��&`-7Ԓ�G3����y�~me�t��|L�H��.�$�"B�s��Y����HB:ʲ4:	�X�U�i�
�3��`Z��=�����Sy[�a!�0�'I$��3�Κ����J��%|��륾[y�����w��W��,�e/���Gl��'�w&ɢ݊�'��NY_��(���;5��#���/�+jQɭ7�����D7;{?aT)��^l��M,�P]G������b�L�9�V��OW�69�\�`�Oc���9�V�-~�Mge4��C��$?#�R�X��$hb#�+"�;H��~�4q�,:>�y�ß*���������ek���5ؙ8��AJ��~�4�P	H��d$܅W��b p�"Q*���?[�`�B�uQs?��z�L�3��1��hu�K����幞?�а�'Vv���DP�J��i��<�k`�^,	ijq�D�/����)s����������4Ty�r#�˱6�g�i]��kESy�~�C�+j��]���W���I�SVƿY%�Ή8�_��*��<bP�[����Uu�%���	d�=p��ڎ��8��DE�4 ��t���Yg�N�yV���VO��4�/+B��Hpv���/A�2!��1��ȥ�`�⍛�X�� �V� �_��s�^m�0W �N2�Ь���~}���BQ |1r�˹�bhi��i��#Ɯ����+P,�4��������U��g.r)%���.��!>h��NMS�
K�_�Z�%���"�KE��;����æ��Zo���f�8š1I�W�?$��]�F)���_`�pp�_,
k_o�:�)/����v��^�����!��!C[B���T���&�v}w��������x�0��s3r�����Mdv'O�G�����K� �W�i�3�0LH�7'W��D�~1��4���H�mku��FA���US����14k`�օ�I_�s4�)6L��_+N��)���4.y����r����=���
��B� z��zo�����?�I�z+��� I� ~ۮ��S�M%���| �L���,�B^�ɒ���o����~��#�x�rp�<UJ� b�����^� ��úH�K��,Hc�h�5�#�Q��w+c�zy� �/�=%J�"��#���3��s�ʶB�v`��<���2�9�w�4f0]%R�5�e��bgK�� �a'�L.%�c2��a&�ܢ�#�	~���8�nQ,�L�������q��%Ɣu.��=f1Fd-=I�7ؒ���s�5�)������y�sο;4���N���׭�OADQ�Xl�&��2�VA��gPB��티�X"�j�%��$��7���Bz(L�fr�Z�~�q6S���ՠӒ2�2���s�&�Ud�D��y�����`Mí]����vZ�B)X����3����z
giF�NBb�ؔ�5���=^6�c��%�1�Me��}k�$�I�@���8�+���j?���P]���C�e@9�7$d�h0~H���T�a�|`	����|%����}ޮ��gV�b�ii��=؉�#�er����	�����b�7�R|��Ub�Č	�?���[��oH)�<e��v~���_pf��q�)�
�^��;8;�_ܦ~(@ :���>r"7�3��m7-~ڳ��B�9*����\�a�"��K�bq�Ф
(����%�s`�m;��e����HN�T,̗i�<�4,�":Z��݃���w��?�m���:�^&Ta���?�h����������d+�#��CVaڡ�EbŞ'�� S�V���T~)�E�]���!��+1�i��%Gj�5��k�omo�"�7�
��!��dSJ�i�I���ߋ�We}p��"CD���KM)�3�y�lN,t�(ڟ�������!N��~��l:�M��N�����ui`a����A��I����'� ���1����N5�b�$��)�ߵ�v�� �i�1Mi�u��k���U���~���5�}[�/�HIj(��9`<�]?fB��^e\דJ��=���*�؂�ϩ��Ml�}g�\���"U��>#�tq ҭT�Iw�MS��rӶ2XT#t�D3�~���|�%�w���y�8���*��y@�N��#0cZu����wh%�G�`�+CJ��Ȭݫeh�.ܨ���k�I��x�8%�!����'5K��Z�$tZ+̝9��ݥOz\K��ݓ���X��g�n:?e�̕�o�ٵ�U�R؋��@�~y3�0o���?w�>��3�����j=B��~��dD7n�km �b��Ű��h������h����Y�.��.���l�1/p*w /_���%M��i�F���d��j���$��d��ч�'��>i�Y� =�@���w�"�a��RIw�W%n�>����X��q�n��J#\e���$���7�p^�a�m�:���\�9[+���~�%��� ����Xurp�>�((��ȰyX�����lah� e�,Q?I_\���פ%������B��r���.��Bj�����1	�����1]�&�A.���=��0w!���G
C�S��T�7�P�%B�q�T��"�D��T���W���v� ���>Z*�1��j���FD�|v3
����o�d·I��uV�K�����eq3�ShXq�/C�P�?|��O��G]* ^wǧ&~R��Qr����D!5�/gB/�ϳ}<Y�z����_�ȫ4:.+��\@K�L<�r|)gц�뉩�ڃ5�\8�J0�53����!L�k�+�DA���(��"<���Yo��U� ���$�RG��a��=|�F_t��ﺵצ��C7��kjf'�}|�u���T�L^]">�P_�])9�����<��\ZT�scr����*lY���Ю|��?GeW�%��=��d���Q_���j�� �9J�tZv�	2�:R����jC^��Xc>"��@ys]�x�b��K�%��H ��W���7�LY�RU�w�6���ݰ���=�6S�Dr/^�\¿j獔7�yo�ۤں
�l=�,�6Ӵ���$���V0��Ym=����}�WZk��w� �;�KY��>΀���ùjJK��"�T�^���
G��N#:�h*q�e� ��IrR�qG�5B4�M-�a�h,� �v�$�����m�����0�:��5�п�R�����)��
N���g�ՙ�$��a �B'Dq&g�L<a ��z�@��Ѩ:*d@A�wT:�`����]$��z��۷��V0B9����"�ŵN�dʨ�6$��!�.E��\�S�h�1�o�*�O��E͙�|�e�
H�Bv�"s��X�Ԏ^O�0���?W��V��J�d|��YKr�xM����+oR��t7��k{��z�%i΃��$�|>uN��9���n�Jȿh~�2.rπx�̲C���bv�2ڀ�nz��IƇzo� d*=�m�b���?#S?7e��5�]�B��o�ѧp���6�ɠ�r��=��r룤@�!���y��4݆��Y��|��L����7k���f�'�h#s-�����a'̠�-t"k�k�b3rgTܮa��c���f��1��Y���-�$⾳�|�aU�pʵ]$�zq�UY( D-�
��9���������)��x�+)U~Q�O¯'���
E� ���ؐ�T��)=T�����d(8�� ��L�v�ӕ�����t�Dv�����Z�wՒ�V2�&~hW�7�p�f寫�5�.�4��*Q�К.�v�pee��(�q�5��*Ue`8��������l�S��ΰ��Wn�>���s���t[��_M�c,��������f��0���%�-�$gA�MP��꿣R��9���m�z-����&�_��9�޾�?ç�M���z}Q0$)��R���.����et7�Q���i(k�\�x�4.�do��&h��u�3G�d�����l�ꗈ�T�b/�&�[@�:gM�!��S��ed������f���~��j����MB�<����B
���8����=��zT����5/k���S�-�Ҷ��9z�U�A��W�h�;�&\j��U W�Q�~�J |"w���5���Z{�SV��pɎ�D�8�_q�]���ѹ����jy�Kb�u�z�y��]w�����H�S�����Q���&�(�	�M>ܳW#�?<쵋UΪ��^�Ϙԧ�͡���s�w Y�����҄R$�,��K$7q���
�%&g�������ڵ�շs�e�e�Nd��4�)�8��j�Yʈ�"UC�Z�&�X��"f�+�Gh`R,������?YD�)����	I�;��T=���l�vU��*�u�=*���UW��l� ��Out��V-���p4�/�)tV��wL}�R4t̪��W/��m0[=�#�<WG�����uJ��3o!H݆�/����� 1@�8O	����V� ��Z�Zg���|�B�� 8Z��s��b�}�B�e� ���=�h|��h�3��R��z=����O�DV�J�9�a�6��w��@v�[�~��Ƥe�S�9vS0��Ϭ����7� �t0`P�PbW�W�$��r2�?�:��|pǯ���k���)��t
��?���0�8�����&���vcv��OhR��y�\����R��n����*�k���pP8�eJ��B�Wv�ah��u{`$#\����w�`�� U�^��u�b���an�P�-��6CCDs��*<{ cZ=M2�Z��Qo�Nܵ�S�X����Ă�\p㌱'�kA�k����6t�A�_9��}-�)�"�_�F��?�Hʶ ecP	'��<3�W���ΐPs��1
`"A*�?	�-C�V�������Ɋ�>�ݨ4���NRG���7�S:/�d3�=��r�^K�r�};v�i�H�ґA�N��<n}��@�2���TK	䡛�J��}�T�%�4Ki|���l�?���IX���
�[��Y91[��>�JAp��MHR��9��Q��%��8��+Lє�[�cQ����j'��������]�JLTlollXyNyկ}��H�W�����tQqT�~ѱ`Lr��(����܄�f�(mH�)�=��w~V�4��x1NV���5h�W�^=Q�q`���ɴ�腀��ͦw�2VMN9Sg�GN�����s���e��^8M'H��T���=P:��g�#0~֫��V2:��5R׏�x���x�u�Y�'"#�G���k"��
血6����'ԣ]�U����,G���Sr�w�U��=�$?7x���xA�r�]e&<������A��w�D��\al�����*�x䱞��V9`��P��޳�����10_��Cѩ�4�� (�*^����k�x�B���&E���Ӆ������U�l�yuE򅲒T�a���Qq/�uo�6
86��#w�vƳ=6�{��D�o��e��I��2�2ݷ&��8�\!���G��P���$j�k��y�//\I#��d��Cn�k�Ԡ}[Km+�2�(#ћ�B�z���R�ڼ���"���\��
q,�M9�'1�Ȑv}Om~0-J����{�X�R u�=IN|��E<���=��ȖϿ]Nz�_G���au%S��8������.�,WEÿ���/���6�1����!��N,��K3*������ó�L����
�� ��-"�\U���G�8�����jS�ztEG��o��p?��b%O>��SY�I���*�v�y%j4U�.���ovxt�I�&ѝJGA���2R,�p$~R{V���V�@�R�F�I�Z5��h3uc��So��"*t��� &�g�;��g(DS�>[J�\딴ix󕪻������V?��0�t��/<�ڋ�Si�M}$��&uW���wf�T�G٧3R�VV�b.\oO���歨���cS�t���s*��l��8�U��5��9P��=g!Q/*�:`��m1ꢛc�2u��|��@Nb�5b\��fΤE�J. sЯ�R�zM�ryo�GU�����O92�KꑢÕ_�Yau#07�f�Yt���7T���󯃄�z����uûO��=W