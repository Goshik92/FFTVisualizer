��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ḱ	I*��=z<��t=r��,�3u�:�S�$,���z�U��U@��z�2Mn�������1��Կ)�y����>�͓�$Rb�T�ݩ>,0�J��|\'�������}�fM7�*{]f�/)1�(�S �:Q���4�vS��S���/"��s&�F���XY�|R�ƨ �	Q�1zT۪Η;�߁�O�����7���K��熏�2�%I�K��$XS�C�6����/"�S�+Y�R(1�o<,_ߙ�ʝ/��7��'z�| ^����9L=t@U}$5���3.�P��B3�
��碭F�w��:9��0�n0ٺE;Y��K��2��J[{�^�h%w�B���U�k������.��vL鄰t/�8W�"��G�V]�X�;���w$~ԝ5S�n[��a�����;�� �u���0��|Ϛ(��� ��SI��v7��D�5�+�}���u��q�Wrǩ�?(�E�VU��+���^bz�ʿP�
������dz2����qQ�I�0��YB&`D�)��T<vɟ�u���ͻ�;�rp4!On��BK�a��ݺh�t�TB��l���y�5i�O�%L^��:՜W��0ΙK��TS��S=	��g"����Ꮪ�������5��p��cE�D��?!DH;$��<,'}��lJӯ�?�aJ�����t��S��K�����%�<YJ\H��}D�wl`�>~
ּ����>�@�e�`�/�.�|i�D&����O�����ؖr�Ɠ1?�Ζ���H��%�iB�1�Ƚ��Xrx�p���:)�WG���U�S�ݑ#�����'V�E$�����q;K1�3�9����3�\z����i��S�Ac�-�Lz34qa� ���ӏIN}�J��8V��F�����Q" E��][ao�5*;b���}T���2�Zr��oԽH�D�{��;ȉ�di���b�١�3���f�\2�HNmL���:�kdg	T����>���p�>�@���-�������^	�_GS���6?�6-��/q���(���}����|��Y-y��&a`M���Jj��v�1�W��\�M"�'�����H]Fmͥ�r���CD�f��P�o��;T���<k$4� ̲�����Q��a`3�j<O|A��K�!�����/��v�}d����&Rc��9���fu#	xv~��e$��dFQ�c?��,E?��fP��	r��/3��{]V��Z���ش#$}'j��"yB��t�d� �'\(�%���(^��Xj�������1I��	�+q�Z���O�A*�r�a��-����[>���C&'O�J�|������'>�T/��Λ����Y�!��/��?k�[ъbtn�/{�Q0/6~+Kvi��?7 ��&�>�{T�+[L"h���j�/!4�b���޾�	?���"����#���ŉ��'�f§м��a��Q|��f����%ti&��l��	;�KXn�/�����X�sLT���)�˙����-(��
�aD|�\�HX��:��mKn�!��Ϯ�3-�#ٚM1��h(���G~��*hGs5�->�@t<�hwj7�� S�(S
��L�'aH�4l�y��!j��X�Bd�h�_�n����z�N�:k\�ݶ͔�(���H�}������:���}�9UG9�.����\Ax�&E��f\�<�U�
����:��4*�#�ߨ��6Dq��Or���еZ�9WTl��`����5���[5�d�ir� ��E�3)�| <��Ca��X�mT,1@�ٛ<d��7<��� �V��)`6��`>4��$f��m��������C	��y��ttٗE3��u5r!��Ғ�q�F�]��.��'{���{7+	p��2�������#jZ�&�@�*j�Dc,�	X�s����B}�S���9rS�2�2��;��1�G_u���C����/cE �o�T�:7j:۪q�k�N�5����;~z�bQ6Դ�'�榍�40!/���=�%y$��8�lyڂʖb��;׽0��ĕ���e��?�d�
��|����SI�e�8B@g�ॎ8�WS���u;��:R�݁�D���"�����7�馾4o�� �"˶��t���E,�������s%��K�I�F3,`h��,T�I�>���5���l��(�c��>���] 1a�N�Zy�$��h���c���R������-�c�����
{��E�jK� x{4���[�>��G'��΀�u����AC �8������<�U�S�"�ɉۉ�V{�R���V��	�(�yeh��1�? ��� Nc� �SWn�x�\g��1p�e�M�=n$�+��^�릝A�/Ǒ�:�,&�S,���F@@�d���R�8@=�tF��%�E㱦�[Viަ}��F)o�T��C2������o<�{L�Y����o�n�?�I��<b�*�1	�7kx�ٿ��H���z6�҆Gؓ;����О� �lY���En_����C5ï"���n,x��b�!�U��4�gq�*�3�&��$L�������i|���;8N�Գĥ_!��
��u?]��A�Ȝp��	w���_cYĒײ�UT
D(B���o��E5���>���n��S�3\ �����2kea
ˆU~��F"&��Dqթ{t#j�����$�g��]aw������P!Kj0ݐ�g�)�q��W�-O�*\����ێ�t���@R�����Q�"O٥t���97�*P�v��X��BK8^�~�[��*r�{���I��߼�>)�n��>/'�¯�X2Z_M�~#Cw�(��'	;����&�h� ��$���(Ym�����Jw>T=I"b�	'p��{w[Ry�޿f�-���:��c�S�r��!��L���Q��oA�?��x����z��vY����	������G Պ�[��-`H>�N6�uO�?�fu����I��9��h��(t���co2��X�*ͪ5�x�������|��i�j>ʞ�}s�b���9��5\�3�����ٖ̽���=����/�f��j�E��X\�4T�[��\�tî��{�ϟ����Ŧ�h4;n��E:Դ��b^"^(�T�Kkw�ع�j⫪��Y�j���wJ;J
ە��hߝ��{X�t
` ��1|�1�N��!�� �����,���lN͹�E�\�>�(���ϊ{j��L5��0m�MM�h�U#�"%W����"�LQ��@ ��ZR��6�.�(a���>�I��R+��U�h	�@7�������%�!�r�C�l�_�L�c���%�Ŏ�,�{$�w9�2�T�2p�M�\GH	?evNl~�u�z�ܺ0?�X�l:> }�*�BMC����e�0�]��w?�H/�,v����/v���lb�e5�_�ϞR�'���'?#���R�c��ShQ��t�of�ֲk��u�at����ZL��h���Y^xT����i����Yne]�KuJ���bߟx�0�WP�0�������NϥǪ^ �8j�쭊,T	ޯ�#��c��M�qz+A,N_��zfS��bXE�k+���A�E����r�*�1s�M͛p)X�j�ӜՎ���}�~)��3̥�*���q�FM���+�	�Sa��q�4Z\��`3�{',e��9�~��l|:3��VW��NE�ѼŹ}�xa��fF�u��X6x�_�F�C^�[�l��V�J`�d�H����kr�p�N�˫�N�)��*�d�M�]L���e#W�Ǡi`�����*Qg/!����*<�#0�CF�JvzlR��zM�@���^_2�v���b}���6���v���Aq�5|"*����,n9:��p���;�d���zh�A��npm�K�ye�^W��>V9�74b���Lm2�w�+\X�[�5����9�imD�n�5�OѲP�s3�ŻQ�o��q,�=O��E�
���  �$�E�R�W�y�BY�or�$���IHŉes����q/���J8�Ҵ����<��Z7��!� q��ӌ�d^C7��eT��
U�������*>���"
1Pd����H��R/F�����_f�C0B�3}7�������TW�%�qkݠF��[�GZ�eL:����
�"7�e~�c.W�/�$b ���	X�N+�C���#vl6�����9)[ȼ�_��H���rP����Ŕ���Y��!p��c(�a�x����3AK�<�s�=h%S��Xa�Q<�����w�R�t��FF��u�GGe�N�u GMv:Q�3�B?�B5o��[���� Pޮq�[zWf�̶U>Ƃ�����	v�;E��/	e�x�8�}N�Z�,���P�`R%-d�3�莢`�{%)X8���j�W�^|�|]�9���Ԯ��[���	$���h"�c���-c=o�FPs%0zKMD�B�	��+ü�U��yv��m����K�_l#�kR����
@�����*͢쾴�	��>)�K�T��ȇ$��2����;�__���ޗ8�'}��c���wN��n&���ʟY�-��i]8
m�}�I�6� �d?4ϰ&�|�jp�lSbD�0,�]8=o���g/��.]�dG�.+���Ԥ�N�U:Q����@S����M]��w-�����a���}:B��ޏ�B�&���f�v(T�wo��ř���h����~������4jo��b�Q�k�k�z��|"ꢎt�C�`�zAva� V�Ѹ�ս�({b���$Mp6
^)��H�E!�p�����a%��W�2F��L27|T;�}E�_��I� 3�|��gD��4��u[�5/��|�<���4��ɲ��b��%!�c�P�P�*��J�N�L��~�Ӽt4A� �l�oPB��]��0��l	��K�6��e(i�:�؊lp�ޯH�K�(&GE�$�a3�S�۔�I�]/s�B S$��jsu/uZ��0,�-Ō�R�<�g�sf��¬���f��I�1!��r� ��b+jMCs�\u�f{������9��(�פ����KY�gA2����Y9�ۙ)I��7��J��-ؘ��e�&��;�LCY�y���6����8Y&��2!�X#��ڮ�ܾ�������9����w�,0
���,w0�>��@��
�c&\NS.��v���!̨���+���@�3~�����}3q���(ɰ� wp��u�618���p�.����v��3��������3/y��	=��9;��t�7Y0M9���Dv��a �?�P2� hg~��;�y@Q��n�蛓k*�^���9~Sw����i(_�X�5[�SV��Tκm�L�{72�zvvР�|&��u�M�e��
�"���U���� �7�I�h�l�R�O��2� g������P���|V�� �}��tQ��>};�+ބ/!�(�-�%���ՙ'�Q�S�k�:�BW�b"=>E�tU�7�#�+�t�栰��:&J%ԃ�qZ�؀b�w�'�\E�1+���Z�C8=�dQ�x�g�f�+���B��?ҥ��� h�z����dӴ��5iI�L���J��_��=9:���^����m!N���5p~��%9e*��-�c� ��f|�C�1�ϵ�ōi��=}��{���S��o�hun�����jj���/�h 
�s��_M9�{�cU�T���bY�k���X�MI�����St�= R;��𚷒��E}�aK���j�ˉf[���Lե���.��1���1i��"*��nX��V�/�)2�ċo�9#c����E|�:�$& [6�z2���Z��0���O��_>V��D
(�N 2��2�l"����S�h��q�7r��?�`N�2B�J���Z��r�����*F)&�6_���Inc�8�!;-�Ua�<���A�x�m�ҍ�ܒr�UI�P�Z�����7.�
����7"_^%��a��+[/���m8��"R
E�pP'�<�S*T���*	P���)��'�ӹ��tr;�rl��f��4A9���=��<�L��&+��yظ��k�)��ώ�����ߪ%�e��4��n�B�b��)ǰ�X0��u��J#^4�y~ԥ�G�R�Y$xө�:����q�wZ�xY}\����-�n�������T+k���:�?��|����<���3N�Lo�_^���$���H4�C�V�����~�y(=�i�Hs��߄_�I����=|hv�_���lA�I�A8��%W�;�/=)̪mL���?v�Ɛ���[
����~6�sA����;�!�E+vo]�_4S�۸��u�|����	�ي{�N�WA�=�{��7�3{iP�B����ö� U���J��ӯ��6���0A����_/QM�#�a{RCQa�PK�>��S�}Z^��ljg�q%�)�%^��i�>��EF�@v�A>�5;b[T�Kf������-��mi[%���칭��1]�h^B�U�� �I�|��[RW�^��<�!�"w����|$���\��n8Y��q�U,G��&��c��2k�+Z>UR���k �3& �v&��H!(~�q�3�Dmܾ/Y��<��=�$Ժs�U��q�ɭ閂�����@g*��J��6�&��k�5�'CiX��d�h�M��g�>���uA2m�|A�m3�߰�V{UnD�y�"�d�.,���8��]��]������r}��(dL�oe��NkVS$�q�b�ޝ��ө ��o��ʋ_�e%]���	�n�{�p���٣U�(�s���2��j#��=,�"�7ED�晭T�8����Lj�@������͍.&j��4q�i��Q��t�/��q%��u)�;*�SO���~�p.-؞���0��\�8�C ��q�x�,I*�㉽���>�� ^ �{]��iO�/��c
1�O�Ε�:&I5�=+��S@���@F�&�!`ӥ��X� 4��TLr��o��QO17_|�Z-�%9�5��"mi�������36聓ıvdas	!X"����%GQ�[७��au7��#z��-������,�ӾQMpژ~9��2KD�_�v�Wꂈ��,����}g���٘\8.a�2��Z�D٤��}���w�����/�3�N(;�!H`�|]R7�k!�h%�c��\��m�OՅ˯��n*g�!h��v������͑���.����%ؘ^&��A(�C��wK�Tx�8c�k~@��,.�ZɓOx�C�v�\�$J��C�p�I�:xZ��T"w[ɇZ6T2q�  ��1��Ձ�`�7�*��8��������N}*�O`��L.�9��������0"ͦ֌���}.)�t���pVށ;���"V-��3!���r�{5Eш�����L��m�O���B��?���z)��b��V���t��bW`��+FQ��,�ID��:���W���ס:���/�ʄPO��mg�*|�yWpN�k���W����g`k�L��E�Y���J�Q��Y���9��ϣ>��+�W���t���zXH1FL"�
�b��n��߆�jTN�	�&oH��i���7im|��)������ �R���z���0ɴWpF~{����Bn16=������-c�����P�2d��d,jT%AsH�^ۏ�e>����)��D�������9�Z��˖��g� M[g?D�ki��ev���C�.]�f4یz=����$��P�V6��V�d�j�&���O��2w8`����z:�&�(!��KR���7a@S�[�Ky{\�lʋ�Ѓ9T&\��ʞt��>������_��3ou2��)p���7�o$�ɠ�(Jk�=�%(���U�غk�_�SD:	���be0����(h��mS�C��{���:�ŕ��I,�ޮ��6��	c2�t�\�q5$��`��2$�J1D���|*�'O{J�̆kr&~m`�4�w4�6��s�Fp������B�%n���iη~2����",�k��D�Ī��N��9,Ѳ 8���J��/P��ը�率�-�ы�Z�\<� ���*W�\
��f�~F�G��Ȣ;��� he��s��ͱ�ŤL��&�.Ym�mǴ٤=�c�#ȳJ�Q����ti���1IR���Er��K�/!	#IR�h`�TXE�l���
�-B�<��㳄6&Y��{��Z�����%bQ���2�+4�=ܠ�W��6;�_+�"���V�-�L@�W��9���i1<�n_�m�'��+�|�h�g	a�ܿ�g˛q�x�	����0#eF�&��J!{��V�_�.[f&ޘ\+%d^|#�BLp�q�v^l�
2^_���G'��ol�5�[6�[$�E�?]R�Cƥ�]#+l+O���f��(y#|ʑ��o�8|���j� �(g�P'�)�A]N:F	�U����O��Am�ᡃ�s;	H�D��j�mK BA\2���@�����\J��sTԋ�_
�l��[�IV}�pݠ�:���]PUGC���P�E�Sby��b �ACX�������g��h��+M��z#;MΪ�L����Gｲ�?:&>������NG�h62�>�_�1#5�!�W�ؘX�b��Y	�9�%�Z���Y��H❒�]��`��Ν��X�:�dJ����ێ��rM6��_I���%pɕ�w��)[ �v�R��P�㵌;���` ��tI/�#n�T �#��������cJ�5��oࡽ�����ї��_ȋvD�S�$P��o��2I�zC�`-r��ʷn��0�JȮ�a�$+�$Ҝ�u�W�TR�v	�,.La��Y�K�xlLaw<�@�I|_!��RaN7[�BI��	��ɕZ�09�͌�%� ��0�(/�d^4�[��ʞ-�87�_x�R�FE�{��"t+���"�#��͞`��L��6�uy�B�fw!!���!r-��!�:�K?8�#m9񂖫!����p{|1��o�
���=G��%bo���ӒC>i,��PI��T��S��fע���[΀��Լ�?��Ī]�W��[}9��}?�x�3�<�,�y�M�v󀤜�L��|N�
w
X����DT��u;�lbm������0��)�T�D�1��T�[�"�e��q�jT�ґ�4�!4O��=%\̰������[<�g��N�b�o)�>l�ҕ�����_��09ڂ��i[��#^�ꈯ�#-Y$$�C9eY6��p�����z�,�E	Óy�u�=x~�P���[ܾ���]�t��3ʚ@��щ�yˉ��J{?���q�<��q����Yb�	R��pRR�e�ϗM���y�C�%x��\�PF�#~��T��-Ww"����?a#��[��j|��*����y36 ȕ�x�i剶���n�*�� �V��̕�̤�6��ja'�jx���s	��sg���ݸ�3��=J5�'�sY�4:�*b������b~��G&uϞ!ƹ�El�'���%v;n� *&Hm �����R���[������n{j�}�r��S$�ֻ�Q/)��]�� ��w�T w�$�����	v2����FM-�.��ȴ$�ȸN��8�P�*n��!Y��ί��#`�٫����?w{_��(,��~��uJ�P
?/E26G$�wE~�-+Ufh����2b�nџ���!��^��3���cΔ�v]CT��&��Ȭd�
D�ݲȭϻ5�jU�.e�x�
�W���Ж9���8����1��R����	`A��hR��*���#9�"ᅁ�l*i�??y�?���M9?:քsN���F�f�_06�ѻ^z��[�jx�)����r�Tc�d﷞S�ckH	�?7�`�n�����~�v���vdR��X/��re~Rb;�����^� @�#��Rᑄz[�O��c�5��������C���
ɕy���ߑ{��p�q�5�s���s,RT麆�4�C>"�dk'i��F��G��Ȭ>b݅�s����]e�5HWy�,�2�@f�6& �[chۤ!^BH���_��qh�q9�(�$+��%��h�҂u0�b.b�Um}�H!���6&��_�2*LyU�����V��?�uЇ[�x���GlA�P�{��E+*f�vZZ:�O_�9#޵�nL-�H�j=�ת-P_�@*�ПK�
�'�S��d�LW�i�H�44!��Bּ�4fۢn'�ͭy��F����X��E�g6#��%�BP�X��T�7�#�b��)^���k�����x�fa�q���&��oQ�Ķ��b�����������psy��A�y� �0�W2y���[c�n똳u�޴�hT�wT�삫�]F�&Jt�		�t�X.�dn1
�I"ț{h��sk���SN��;�+<E %q��b�A(n�H�1�pmY�e��d;|0¡됂~̨�g@F��d9�ItZ�/��<��/M"�c��F�iK��@�t���Х	���]�>rZbR�kb�D��qO\t�2�zdgW�6�*��b�τ9�� 圸T��qZc�Ñ�h����%s9ee�cJ!�C�p[1��6�NҜ`j����J��!zg��gQc��Y�l�8�#�D�]~&H���C�����Ģo�h�wc�w��i��D�N]wu/o*ߔ�\C����g�e��A��0��^h Bû�+�`����	MRi���@x�s�	����F�ե2K�O.d�aƦ�mEi�������e��؆��̒s0:�׋���r�E�ML�{Y�M.�= �;0��:��Us�ə!�����:W5"��0�jrض�6���w���~��I���ɬ���r9e@���$i���5���z�?��?W4*6�Z���nu�@{���j�Y�s�VDk
=p2P����x3�w5���B)Ý�J$�BԷ�X>��,y|��bҺ�Rq��Q%u��D
ۑRgr2�&�J.G���D4��T��}G|l�1�փ�	�$�3�b�#����+4�(�;J�)㘣��
�H���!P嬸��ƅ�,ОԵ�9Y?�Ud�9T�P��9|�و/�}2u�P��5��[-J��P�
U�n�ʴz��_
q�'m���9���B�1�q�^[pG4U�ӈ��~Q�xq�p����-w��r�B#��,�R V?D�tz�R<J�j9�*�ȟۤ2�oe��0� lR�X'�꘾���7l��A;Gt=D�;45(n�(���+*���c+��C���B"~�~`?G\Y�
�*~��(���$z��b9���N�L����O���IR��0���67i�v��U�+��nvcMw�,ܞ����u�����aנ|�g�KN����(��z�ӹ��]{�k�����B����n�	�V� �Z��x=��g*XS-���"_^Ӻ ���O�i��&;&ĭ��ڛ5������+Ww�=
�G@��TmT��{��N^$�጗��v��Z�ϝ�31�%]�,�J�G�4�a�M�OdT#~�QOs��{K,T��מ!�t�;"����Ļ�v;#���エ_����E�ІH0�3���������l�faaܪk��w�G5+��ݙGJX�rD�c�(h�Q4g5g�V۳~J.4B�yCE�W!��.Y��X�!�����æ���J����=_���x���]�5�a�%�����.6�|Et{n��F�H�<�E�a��M6Sx��3Z������( ��W�M�4YZ����c�,���w-����L�bqrd���mhX�����6[=�/�.%���pgP8Ov;�S�uX�j%�ƴ��}��U�.�]�B�q\���_����'���}]�<���흸��΋��[�NKv��b����)�R0�Ln��^sQ2U4*Ǝ�G�{���љ3]�<[iT�S2�m1��?�5�� ʈ��1����s(�&����>|2.���K�C�;b�D[a�y�YZ+�u3e�T'A���c�p�Sh�/�c�A�q�!h��A�%��Afr�Ӿ@������9Pb̽/^����Y6�&d�ú?�@����"&�΁�ǯFkBz�&������2�&U�\�k#v�����ј�Cx�eе�]y��P�Bz��Nᠯ��D�Y�;@�{��`�v;���N��J�Cc�̻�2��kA Mi�����~��n�,!�Cŗ�]d��zO�V�0�V��;#���|35ޓ�6�;>��k�r%rF�@��=�n�UV����s��s���d�s��GMqO��6>K<4cz��S�K�x���8h���/eXt_��ͶJ{�qb�?�F��ҵ�O�R�YY޿5��N�Br��085�����ힹF=��G��c�'/�O{M0Z�I{%�G�
����g��|�^z�)����or@|(7��g��ϖU�>F�l�}=�g7�fξ�rگ��:���G�ݼiA����T����ɛ�S��@�㍬ߣ']M�k�	�I"�r�N{�

�����$U}��Q����#(�?�@b՚,��7�hο���=���o,K�}�~��&�����2��1�J�_��o"_?hC��Z�pv6"��&p��b�4�`����C��[��븼6�{�6{��S���a��y4��"�w�(j�O����&늆���"�c:x���H�)���C�fi��0*�u�a���s-��/�	�'Qw �đN:�{�NF%�&ǃ�$3�v���gmQ��`�g�/#����2��H���i���U0�f�'Dj#����g���V�1�BږUMZ ���p�_M�s�ӋO��$�F�G�Kc��0�^3�ʁ*�f'Wg)U�>(��r#o�D;��.;����ڀ�EVu4�y �45�o��~���I��)܏�۳2d��[d��.Fy0lm����NCwk��Z,�"�7 �$E���!��ك��u�Gi��<y	G����)����r�.毽_P��);��to8�@i�5�stޗ*�{�)�\*�^��D⡏m��Xo=�9����܍A	�/�f����><�ȏ�e�ԂQڎ�^k�H��Y�	D�بaJ�QKF	ۂ��,�%N�U�D��{��� �kN�c�![�-�1�&�x�����t�}E������psR	�2O٪���k��~b;��ҕ����z؎��v�M���W���)�r_&ݥp9 �,��
��+^��v&����S�����ZKw����f��Oj��ڌ��e�=�������#wT�UF+=�P��<9�s��r��G�ȷ�P�}���~x@���*GJ�Q�_�u�d�Ko|C[�S�*i�6��ĘQrvQ}��v^>��U���H�:T�'bT�f
��evF��G��B�#���i���#�;p���u���L�&��0���(�"I�g����������6nܡ�Q}L"j
]�/�>���o�A�Q����\�`	�W"�����@Z�ӄ�7m�ju�ܵ��nΛ�Q�^�<˂(�`�W��p쬔@��	�������c��N�� ��n؃`Oѩ@���v���i�R�L>b]�~�Y�&aH���P)K2̊K�82	O@S;�z�$���V�ф@���_r��@+R���nW\�����GL�U�rH�t�`'=)�	>� ����豞��FGjOD���!��~���x�������\9�����5Dw� ��;0I��W	��o��D0(9 �	P�3}�;(�zewf[� g+
$c
��J��&��s�`ٙ4a�3�;X�yw@�),�/�����6>Ȕ]��I����2J�!���>>
��l�ڷ��%��x�W�cD�/ ����H�e�4����8U+5�~`�{��#kX8&)Ic�J$��k��9��M$�):³X��!�~�1��?�@?j-'�̉БzK�)(󸚡>d��s��	<F��n���78�K`0��w��#�^S��{�p�ǅ"���i�;�E�Q��}/������=_�t�*��ژ� :3E�7�jK���g���w�'1��Ak��]I�Z�S�L��#��|[лG�gb9<�nq������������Hv�6��N�=��}�f�c7��?�(�ʯv������'�/�]?��$��y^������]�R�zuf!��n�9����s)G�U9��OG�GSL�{��Z�����	����GG_��e)Ѩ���6�G�۔�=.�����s�~�,��@���˯��^c0gxNz/&�Т��b_�hƲ��iϡ"�7yK[�&����m0�����~l�Oh ��uZ����|ɲ@;D�6Cs9̝��v������+�;�����3�z�*b�W�SS,��,�o,&��X�%q}/V��g�>�mc��������؅|j�W�Fgd=8ص0�яFƾ�@F���E�q�M����E��$ (S���	����Ueo=���
Q�p��ɡu��0�j��s�Ǧ�����ٝ:���f�uƎ�+��.ev>\�U���%i����jx��e�C��OR�pd���[V�wӹ#;�,�å�JH<�y�3)F.Z_}�J�edB�Qj�D'�x&���9�"=g�&q
0�J"��-2�X��8���slA�^�ډ>�;�rx��\K�`v�d�ml�
�2
�_��ԁ8r9Du�]H���� � �@K&f��	�֜Ʊ����[ �Ty�(�^��Q��_ۢ��Z+���������,�t�.n ����s1��j�IRiB�����=�hVE�;_�J�9�R�[]PIófKo7r!QL����+P8'3�������	����O~Ȏ$d-�wb�e����M�8�*��v�R�о@���<}19m����N9��j�,]S�vP~��y:	��G�W�2�G~�KR�:t��X��T@� ��č~��$.%�7��;
�ZϦƯ��$H��_q�:�D�z�u�|p�>j��Jp;�ɪ�OHBP��K�AC�D������B̕CH�!��Tƹ-/��lH}�'��[���D�g
:����ߙ��[�|Vt���A�RZ���1�J�4%F�}`�{���I�
薞b3�\�z�:�����/�A9!�?z�j� ��/v#���(�熿�w$y����v-����hl�c)�:�~��C���$76��X������ݤ!H�5��N�j���гg���F6�7aGE.𽶭B	�b����B)��u�en�Z��h%1kPy�2����3AEǪ�?�c��m���y��F��Ȧ{�� ���,��&��$��t�㩢�B<1���=vϧ�Rm�tf؈3s�g��̋p���v9�K��KHԄ��ɫ��?�~��d2�R�%
$���C��`[6���QA��c�fB�u�d!�E���9�o��2�e��CG�b7
T;[_���ڦA���p���GU��J�� ���.�)�h(��&]�Y^[)�Ӄ;N|a&��t.�$����/�)�����0��1N^��R�cl�����bq�[�@��]��TY����eǽX�
������Ȭ/�No��͊�s��fM|�"�kq���2�>.�q��?,p1�?�u�H�3*XC��G|��Q��K;Nʴ$��҄��`��l_R�*�ky�>W�x�A6WR}��9�=:�`��y�#�r���w���!H�z�@�U���W�����&M%�c�~��\w^��	��0Y�6�PBf��.չg��/i��ݒ����i{(����TZ���#�P�e�zt�R�,T/x1���>��QI&VJY�/(���:�-�L�a���M��d���[">�����I�1)1��>��c��v<,����8�H�H�����c �|��w?'ϲ�Q��"!/ �5��`�h��T���o֛���j������1�F��d���"5=��pq>pCԒ|��ە��W��� ,$͓N�`Ѯs�=f�5ƹո��S��.~��YLPl�+�葅ߕ�� �S�h4�U<-62�-W<��\r�ܦ>��v�,�¤Ý۫�wh@:�6H@���F����LZ��=�}��g����\n�k�Am�ͣI��[�q`��(.-�Z���;*��yR!pn�h2�����.r���G�z�]�+��O��<��GǓ�og������6_;aT�Q2{�[�vX��˳KPA=4��X�9p�����	�� �<�@<o��4���'�41�Ie�
��������&�!4E!}$ʁ�k�}0�m����6�.tAӵf�5��#V,����Tn��W�.!L�oLḀ$��<�����d�#-��@��������K����}�\X_�Q���i��R�ܛ�ދ�]�r`���� ��r�'� �5��Ԗ�_@av�|�h���
�xCH�^O�"`���i�'yg��b
�������{�M	���3L�3�l�-�%�h8_[1����R	��ˡG����t���eY`^YE�|�ڜq���r���+>�YԦ���7{���b�K��)w@�������ݽ��I	��B�|�i�iK'�]�YgDҕ����bW1v�.Ǟh�w����~��ˤfVb�g�����\�b�H]�.J��e	8��I�����;�Z2j�
8ٴ:��h�.VǨ��U��R� �|ge�`���!��+�F�����
/��w��2����ߋ0�ۍޘ�`$�T�@�m�f�!7G�K�U���� ���B=^��4c�"���"�itJq����⭃���&���!˻��_�_C��T�#�0�O8/����JT2I<Q3r�W*�%�d��#(h,�7ǘh�YT�W�R��$����p��f�Fq61�ug��Tm^��'e���?�mň��%J�õ�����CJ �a��;������r���A@��2l����{�FX0�E$t�?vc���X�>�2�{N$�E�&����[�<[�\�s�Vl�p��%�����U�]z���妲�&ӄ������˩��0S���T���3����@�We��ЧŨ2�bڌ�5���u��z�ߺ/A����0�b�p|N'zm��0#��B0X�j�9��(7����n������t2"��^��OxK�*�8�5�G��b���C[�Y�#}Td}$��=���mZ�e8���F��c�j_?�Z�r��t2󎩔2<X�y ����z��(M(EM��+���1	�f����tt���p���	��]Y�d_wH��0����.�#J���]��O|�X��*{+§܌בq����p����R �Bt��d���V�f.�`����U�~�$c�B��-���1�����O���qv�h3��DO���&�I�ϴؔpk�_bƏ�<���G���������uO�,��P$7�W�/9��s�"W��B��О�#����s���J�ɫ0;���(��F
�ߗ2��ww\����Y��G�Z,B�<nQ��;����\QUf��pG��|�Ζ���Ͽ��؉A�+Sk�EMd|��LN��RL�OY�4P���#Mer,[J���#�f{h�@�~�n�TU~w+��N]M�`Ra�4s;�9$�+uL �Am˩�i�.ȴ��=�b�������$�UQ���N�m�Z�ڻ�+sϰ����S^{>$.�m#a�oL�'�S���b[ls��e����Ը�v�x&y:C6��U%l��>@'n���Ө�D��۳$2��a� Ȝo%���\��v� �}���rx�C��r{Wܰ]�8՟���&��&����8�����S@�T��	*޹q��M_�B"�՛���[$�z�<�,���|�W}�U��>�+������O0�6�i��| ����v�2�'����7��9��ƧOOG�\+V������`In	�g�h린�06"eD;�g���R�����qu^n���[?�ǆ���?~w*5����i|U�7�$��(_#m���D��� �9�:Vٸ��ŇWaNۿ�RP8�݀Y�Ͱ=�E��I�����R;�B;JW�m�����%���RߞƊ��N	�[䐤��׸���CQO���s�����Bǃ�3�1ʃ��3��0-{��tii���p`��_J������%�
�ռ�O���jB��΅\P��2n��B�>0�+\q�9�֡���n;���١���N�H]1Σ�od���P�����Z��}�a0Qn���|������c���NĻ�ñx7���w��p�������Tǹ�/awTX�6���V��j����R��a�����hj9%�@5C����:p@���{�!��~#ȳ!~o����q3�.�j�[6)�M���}4d�1�X��ԉ)
��Q6Y�&��Ǻ�Z&ju���h>�E���l�f��r[�E�3���%�r`j�������gR�x�#4�������u��q�}jRif�|�7����2�E��<�]k��#\&l��3'��I�`Sm`���D'1������y������!)��N˚NB���d�JA��������Y�����h�X�Bš�k>�ŉ_������9��tMuq����1,]�І�pwW�~�x|����.�ލ�R��So�z̄H�I�F��}O�v�����}�#� ���GS1���4���0�z����e6�3�~����(v<$�)�Z��
f��da�s:a�/���@,�	�usöc$�&Ǐ��%DG,�>�ߍ+�c
�b!����]z��v1P�|r�2R��K	wp��@IV��h	N�!(�)�Ŵ�T)��^}y�K7���l�I�ɫ$U�n-μ"z4�ֵt:����y;7�(Ǫ�¬�=� F�,`*l��/m �Vj�оA�L˸m��6���s���&��'~�������$oy����g���N��nd�3���Qdq�����U�����B.@ʵ���3�s��f���!����S��߶J?Z����U��jO1���v�,��2$�X5�L Z �0d��)��LUg�j�����XN<���q�c1�KMkg��X�d�tʒ',���\����أ�A�ў�a�n�eC�����	���$� z[�QO�|�7���.��m�*�z�?W�[W�VV�
���~Qvv��,с�O h���?�n�������H��O_x�~�#5!3|3�o��H;�'�����?�F�!�Z�y(��8��c���zאz�O�]���L����!��d���&�25A�8YB	���Q�6��Bڧ�(�̼���O�Tׇ`��ݝ����h��f�e�z�
�}hȣM��)Ҥ����	�" ������kSxD��:��':IB��Ѷ;������a��_�n�F� Y�7M���Ə\A��R�?��/�A���u���m�j͝�`��t��`�[f��q/,�t\�k��P���Rw1*s�w-d�6�rC�^����{�{����V$�FP�a�R,m:�RC�Ɇ"�e����ؓ`wꙁsq��&�3�8�Ng���1�7bҚ�rh?ju�`��@Y5��cZ��<�;���r�ƃ����NB䟔�b�����C��7l�C˄��
�x|9��p���?�O\r�xP!��ْ���Y�³V��d0��3�/Ψ��H�����'z�>�x%/u`�A��K`��~;9�ӦO������w�L@��R�J�ksIf�[�&A�^��R�7��/|��3a�㎫���ݮH���0G�=#���2�(�2�Tp>�a�U�2!�j�}$(��_-�sn����e����RU��6@�����*xX����G%D���t�Neq�˯��`7}
7c���*R���?�!�@#�D�Cz���3�ο��8�(�H��K�hL�D�P�@$��wKO���1v)q�������}�.�͝��35@�Y�b��D��/M10e^W#�=�uR����ܤp�0���ԉ��>�'�m��MGhe��B߄��`�xjh�����R�/���ttU ����c����zljO�z�NYK��;u��۫JDT���$[�S�_hw�Y��뷅���D
Ƒϡ�]��?J�Η���$�p!�z�}����^T�߷C��m2�_F,��ڱ��T-��"/��;b�sǥ>Px�$ ��mż�٣յ���s�*�3���9�E�<"�~��HY���q�L)L��$3���gf6�M��+]��y��n;���ի�(���z�i#����G{���Rr����!��V�a��
�@�3�o�&��Ň[�[�m�ߠ�R�y[��ZS�x��u���5�߅�E�ˊ˟% H�~V�z�UN��D¶*�P�)� �Zn?K@}��15�PV_�f��ԏ�{;���);�u�'�-e#�K0�>dx�;��&`!p����g!@-ٵ����\``�E��N����l�%X��2��x9qg	���c�+���K���j�.�݇��y���lzb�M��愲�<uD���4�����Wl���mJ|�� �B���n��A}��j��&��h�� L�yR��[B�s�PoGp�ȁC�ث�s#�DN�(�e���+���_�C|։��c��wS�X҈�WGd�3_��_yJ6��A���+6��i����M�����K�-fTh]���n3��	i���:ɰ��r��[y�*%�Hb8�F��h�zn�TǊ��2�.�O;�}��r�L�?��*}&���)R;\D;�x������j���2:n=�3�%�f��c��Y��7��8��A�wb�,����l�l"*'*)��Iu�
v��{�	�Y�N�������vܰ�|���,�&"�oq����7��La����F�;@�i��bU��&�u��| ��I"	k3��W)�wL�ՖnA|���� L���IM��0���b���kń�L��W��l	'���O�%D���]ll8ب���3'F�*��?С�t��?��M�^hD.B�*��؊���>>�2{�WUB�o��?� �A	��h/"�C/J�˕����!s�
?`�.#`\�f�F�͝�ǯ��B���Y�Z:�7��3[�
�������؞�?�扫m-����(��Fw@	k��k2��2��p$��N�0���6UM��&}���M��؏�k�ț���u��yJ�s9&�}=��Z1����!ۧ��W���X�D�/TRs�w��۶?<R�ա�V!I]�è^��y�"�ϸ��t'�$\G�'�Q;��k�ǳ��v��G����Pb��o!�LA�V]��Rt�����W!#�}�H6�O�(�R���wW��t����o��8I���ͷ,��I|��`]<4����V"O6�2��6�7E�$q�h��T��ݣ?�|�Ԥa��vg����K3��ٍB�ތ�L��H��4V�Q��Y�m�������������~ӥp����Ke���[�zC���vݵ�����N)8���5$�|�2g� �1�<N�IH@ Ź�gnEÂ�w��Z-ps\A{T��]Z=�:��x�f���s��{w����,t�)��^�!x�����r��P�G�@�����|��^���5� �+<��/2�D_	�t�U&�d���	 �����j��ꁭ�7ޫ���"_+"�A�2��S}�昋�f���/����"ԋ$�~T��� Z
f"p���Q����6�>B��^G�>����?XRV��X�<>�7�K���s'�"��<��pe����ݷL��n��)�+�BR�Y�6G����L��`��Cu��z<�:{�f�uu��<N�n�*���yl������둎��I� 5s�)�����>.�blɘo�$<
.�u���_�'e_G:�� e_�Gu���C�F馽`�r�B�����px`���{�l��̽�,D/�@<�!$W>%`aIC���н�P,'ze�*���e� ��d�:���R�ۣ�����y%�R���2XLIP�Q�����ФL�~�t�����Lt��ן�H[�u���R �J?�%a�xoy�1����α�Dz��ßz�]7�=s�#�pi�]�j�5Or␑B܃�����S���o��֐�)Eg���0�H(����\�	:�C諬��Ɣ�ܽ{�z��P�o:M�Q2�1st�����1�J&�NI�K=x�X��%��w��3jq�Ӗ6�oN�@�YO�*����o�8 5P�K�>�%�م7�UR�M��HH&x�l䊽!�0�u�Eob�h�Կ�Z��_��� s0�:�&�N�;`�9&̑6�+ (����7֑O�
o9���v��D�'s2��6��YL��.�u��u�q���#����&��a�Q����Ղ,�����߉��
�J\��-�Pxܣ�4�m����#M��Ap�]p[�