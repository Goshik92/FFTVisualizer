��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�`��ihۨw0�E�3;�_t+G�����orTλ�I��%��R��	x���B�k��+���gJHV&�D�����ݦ��]��k�4��Cʇ�'�>����犜�ֽ�|H}��|���Y�i���+��ĦIʴ��{�^���G>��P[ް��� ��gg�=+����C�өoSWԈ�D�
��j���tt�yE�2q��^�!Lb��:�*}����%��eKb�d�]��D�ڤmp�T�WЎ��fN�-�Ns�,�E�� �ޟ�F�hӹ��M��7I��&��k���t�h�,��e�{^$?1\�9�����4���`9���;fC#h15C��{�W�r�qg}Q����U_6�|�h�2�5�����o�s��F��>5�������]P�Ʋs��'�7!]���v�T1����)����.�� �˚9��cHYW=����9伔���x�"�OdVڄn\�4��"Ma� �+��V�w6z+iO��{�eڊQ���C6��Y����*#�_`~�Ĵ)���jH6f��X2� �,�;T/rO����v��
4^�v���i��N�V卌+�"HTz���}�Z �M�>l�3:Y��o�+�`k��j �mt��!R G���a�p��3^f��	�AOx9�`	:��G�]����Wh�Y��]��0��K���%��W�Pe��T ��+������v|�2��밆�v}�h���A�o�)+P[;a���4�����BP�"�Qe�aK)㰣\1HId�C�����S���V
�?��I	n�#XG�:�N��1@ƣPO����0�d~��I�-=�+�
l��`r�Y���1T?�:�w{Y�6gO�b�~s{�(�ޚ�W\�9V ,�v��X���S��Si佊�`�M	
�Ws[��;�Ʊw ;�#���&�}��y Tq��bԎ$��X�L]���k����R[T�B*��gf����ʭ�"��7E�ky�ǊL'���m����As���K>�a��ĉ:�꪿�#MT��v+�ͫ-!5��==� ���~{=���Rx��(?�H��!����G����҄�&���c��e���d$d&ݪ¾[㘍�]�/�C գ[[cp�� %!4E����	�|'��d*y���S2m��."`��`s?�5���e8bIo����5���E�Tt�����b�t�A��o�G�r��>J��J�捝*?{aS9PmAkH���[�q<}b���fp�����m���T2�~���0��?�����_�̀�G^�-p�7��Z,�1<�f�Y��w�T0G
�!1Da:[��JC!Պ���.R�6��`&S�/��������S�ʫn�0�?�@ڦ)�<���QCǩKBeX ?�c���0��OU�*��,=�`�X�f��[2�C(�Y�fu7c�-�����/�Z�{����PDI�F��B�V�5)O���)��E�lnK�_�����7MH ��O̐y�hjfi�l�,ӥU�bA �s��ٻ�d٭o��}WUi���a��VjRa�|�<��
:ȴ�xB&��G=��g\�8&+P+�L��	3F��Yg�����A���v.vÓ"��L�nj.�2EV�g_Ct�!_�k�g�g��C޲�r����uCvTo����; ��?��Xp�����J����7 �]j�߳�J\~;�8���=��#�2@8Oajo�bMs��<;�g���x���qO�Q :����{���ˊɯ�#�v��LVQL
n$AWɏ�������F��\[F�D�칾�����l>K�m�'�ح�%̻#u�0d��y9p��1���=v��q=��Q1�Vg�fw�:W��A�\�4��0!K�c�(��Gh�~��A�\q���mF��vLnĬt���ޡj���Qj��5b�������;��&u�_�2�����9 :�W-����=pi ���KZ�Y�j�a�������s�bp:����]���GPFZ9�-�u��[c2�G����6�R��xP��ē`ۗ_���T�#��|��o�|���S��-�S��X�c�Y��aH6�=޿�P�K�%�.�n�5�0�'�2���M����}���@��U|����?.�����J�*B���;�`]�ʸ��7B�� ��>�?�BV���; �h��n�ȷK
�%�`׮�t��%���9ƻx��M�D8?̖!!�z��Ò%>_�B�lNA: �>�6��9 e6�/?SM���O�-��y��E�F[D�6
���&)_Ux'����l�W�>�����0����3�X��Y���TR袱[bh��#�HWpu��A�X���pƻZ���������:K	�Sn���g&p��~*Q�we��HY�k�W��[��,�ᢤ!b�8��Y:�MB�@E��`�~_S�q̘�7|�0��ޢ������\�j�jC��x�M����ތE���	F����Mķ�&�(Sl^���:�a*/�<)Y�viΨW����V&2K�s2)�a��NI�����1�B#Y?~�E�{R�	�������KJ+��ҩE��'Q1֥�p��V���{��+�_W�nBx�Eub���C`�.���w�'97o��Up/>�hp6T�$���f�����n(֢´v�tY"��y�Q���o��-���j��vpe���pt�R
��/砕~3=?�C��1ɞ�cU��	�>Ǐo���j1�+��%�y�RWJJ��ZFw�D 쪀,���s�K�˲����I̾�x�9�
A��^HD͓g�;E��/�M��	5�;�i��n�L�y̐PN\����ջ��qΖn�r>����_�)��3[����cU����:_%�},ހZV4.��ҹ":ò�f�'e{��X_ ��*��~5�>#��K6��r2�M �p���#��_���ǿ��e,�m���D�cK���;g����Ik��2��˸/��	�o��*k?z8d�κ���nK����Y����48|���#��6��[,�\�⛃�]�:��߃[@B8��N?�Ddڑ�h�mi���s`�Ρ�:^�xj(������]*7guZ�WFݦ����4�eFd��1�$P^}��f�'���C�gR�}�A#(�@4nX�`��!�����N^_��c�K� s�_�%�ŕ#%N,J.�E 嗛����Dx��d� r%���|tcU,A����/��$��|��%6��p�A\����h͂7�X�B��=`�iS������'L������W����ȍV��>3�Ǘ#q9G<���l�$�"2H��~sL{�	��X��J~/ @��a��+�9ɰ1<Ջ����Ⳓo�\�/�Y���`y�k�m����z�o�n|y�r��:�9ǚ�����Xo�:������r��px��HR�:}g��,�Ù���ȫ�O�~�|Y3��Ȁ�c�Q�'��6è�����9gE_�5yec.�RC��O�1n����F�tc�*I/|�Ǡ�Ή��1aӿ��|&��WhW����v�(�<��|��9ך�&ْ�	a��	�[L<a�csJ
7bC0�N���jR}�'X�!�[{lb�g��z��6����޺��6a-{7�y���m�;�yWǪ���6}>�g�J��D�2I�#�>=^Qa�Ϊ�?cAݐ�'����P�Ӵ%�r�SwE�]�5�O���K�h�)�CGq���8�[��hF��3똤���y��������w���*�y�{�B�M0��ެ��6�LT	|��SwO�%�8E�f3������\�����p���K�>˾��v��"4v��ȃH.j|CsvYOнzE�SZ��@m^U�� ����*!OB��f�7+�t]c@έ��w�Eu�A��p9��!W��I����39�#��:��޿x�� -�!y���b�rd+qJ�V9�^RGNx���G��\_��b9�~�)�:��!���\X�,@HS�N��·��Φ�B�&R���d�z(R�Mu�G�D0����-�By3�\��tD��4[��D�H�r��)���YG)�r{.��Ͻ�֒�)�0�Ӎ7��j���bfel��"tO���~����1������6�~yP��8,���|2p�m,
��2PSw� \u�LcD/\�)�R-����٤����V�-BuL	fT�[#�g�=��y�3��Mnض���6��?�,_���L\H��Yw��nΖ>��<���C32�m��?��	�Rz)�LEN�s����,ԃv�Qz��2`22n�s�~X�(�t�u �{^�T5R}��]0a�p�"~{셢��h��d~�(�N����@�%�3g���5�	�];��ǨqT$�b�b.�å�=L��R��;���S��E�h����JHp�tUW���Z�'(��H�iy��OG�`x��a�4cǓ��d��A#}�@[����Yxh��0�a���2%��5_�eY��eI\�f���H6\ؑ�i��!+�c>�]lw�P�d�P�/v��K��1\j��5��ҫ	���ܩʸ��/,�\s�"%,g�F3��!x(�!��|c�$��{L�.�|Ò�{�jdu�oC^Œ�j|'���&��}��Fp<��eQ䢷���;��c�>瓺��le���;�����m�x˛F��ݳ��v:���fa^._�7���)�sf7m�"��1�''3�	�a����>惌F�Q`�����ChM�<�
�����q�

��Z���$T��j����-}��[�|̱ˤk`r�|�����G
kM�ٙ@;ꓩv�g��X�1sDfRR�\��͒��b8��Eht���A�°B����7`O��D�n�o@��&���ߗT��;���d;��C�.[յ��N���=����ɳ��$��d�;Wu�G�\4�����Kv)42)AvD��y�<�1��%q]zR����ׄŖ��2����+(�$��Eg�z�^a�)���Fq>�;|�P�3R)FE��,��Y����_.\o�B~��TN�	*�[���������Ⱦ\-*�Ftm�4���A��D$!Z��L�&9䯿�^F7.[=k���-3�� �&��#���Oj�>Oo�C���.)~����=��d����]�����U1l�F*�[M�#U�Ǘa���s�(p	���G�G�$Y0�J�V���yǏJ�j�=Դ-כr��Z�]
4\;y���2(~��n�=rV7t0�~�$���C)�����`p��Ar�cz�L��bCc�ߥ:xH���ӕ�;u�O��T�Ԡ}g���(D���� ^�a��q����?#��%��5\/�rׁڕ�")H�*!�c��r�A;qg�5ʈR��K[|ꖼ������kVpn��C��<�Ezr���cVd�eBȔ��q�MkiP���u#�"I�kNښ�b�y�%�d�6q�GZ��x��~��հ6�R��d�sAhW�#����-⪮����:y�}�	<
V�?�m
��'���;	�B֜��0���Ǘ��#[<R��;l����Me��*��~�XY��*���5{�Z�Й�jx��T�Q��[��pli1x����֡zD`��;Z��{�N �K���;̻G��8A]yV����c˭������ŏ�1�	�	�CÉy�r��7ِ`�e�ʶ�����@{����H>Ş������4t-���K;��y�Q�z���+�3�F׸R��7�zc0�b�����V^T�\A+x.�fr� ��sNQA�5lőT?c~��G�K���O�r��j���
��+���=J�/<�<�#�d ���̏*1Γ�F�r�TӼAty;��E';���>g�^�ua�n��T�$oh�':S�<��c�cZ�)��7f&�e
~�4a��]��˥}*d���m�Nu3����TnCV"3�3��"I8m���2x�0�$��j��%<��5�#��V:��}��,`�䰪su2e����m6>���R�n���G$�gc�w�r��ғ�{a�[qJ�0f����	qu��|�5��7���S%XG��K~�Ro,F�' s~m�������^fT�{1J_Ԧ%gڨ��Jk)�mbEoF5��"E�̌�4��(�F���u���w�l�I<W�O#D�k�����,;T�S�����灣.&Z�+d��Y�9P��->b�N�)\�3�?0�	�-����o�D�q�rοQ"DF�Sũ(}x:�R�����%����#�����6}��T[�?�H�Yǅu��^<���Pׯ#i�,ɲ��M2ņ�c�)��
��a�"��{��lo��ع�=�z-OD��O����3�3���� �d ��RӃ��������I�=f��
���c8*�47�.<K)u���@���vZ�'�_��������Y�65T�wی��i]�l�1� A<�?�q]͸����5�Ď��7��حe?U͠�����A�u�[xm�����oH��,f�1x=���Hsi�����/�G_�ب�UЊs�e1����4K�ƙ�:?�s	)�&�G��\�p�>a����?G�ȲC�{i:X<�L'��U��ת�8�S�V;T=�^�}K�g�l�nr�٘k���hc��x��a�]�����ٙ8��z/�Pi�ȞL�U붖�]��ɴ���ۖ��N�k�9�{�m����( ����h�5lL;'�@b�Zֆl���A����F�0�T�F�������Nv�1I �qd��8�L�^hul�Z<(��G���2��Xb묟�T+1}v� ��޵1���Q�қ�S]\�,G�/\��
 ��M��l�3\�a�j��n/3̏GR\��Yb�����A9{y5�QSdl�`�iy�p���G5��t�K]��u%�Uc�a�@�=�T@�8����s�ss�/�?@�������'a^j��]��{�bP�FS3�oe�ᇗ&��
�$lUo+t��_$����*�?�r�(ݡ4׳�����%@\��.S�9�F�ƩZh\:a̓f�ej�ʯ凫���=ē�#��S�C̢l�;�&@�$�����V%P�z�x` g\.��?)	4W ������$$�J�F\t�0��I/��{�Mn���Ʃ�o�P�>�Xբ�!���{�1�k�$^�c��'�O��ٍ��
����z��'l��JL����?idMÌ5W�B��*�8+�{��V�g��.O�bAG�Ld��CJ7H�2��JD���`�0x���Xf�\���a��H�	$w�C��l���C��]�CÅ��(Y���X�Hs����L�S��U��Xj���M-�#rc���&�H���BkΨ"�R�V�
���J�\�����dA�|����J-��C.e|*�jӟ�#][�ȼ�b|����J[�9_�#ʐ+d��a�����GI-���o{F����Q�I>��۰q�Y���A��>̮�3�<H�O[�u9�B��,C��n�B̤7�o&�\��˙���ϥ�u-����>2'�{r���^E�'��=�R5Y�L�� �k�y�l7@���T��ջ��\���_�G��n�!�4L��S�q����ӥO�r�Af��6�9s�^/�Sl�?"r�s�ES��6� \�=�(��)d8�ϴ�8�����n
���b�� e�NUk@pF-l��׻�����3��`PR��zf�0��՘o����7g��^OnA����x����f�TR�1��t�i����������h��w	��P~�<*�!��)�<���0;��1��]��b�V4�sX�p�����hǑ4��Z�'<8�ivFݗ�ވ/�׆�C��U~o�!+ ��0e�$@)5��[�#ȟ���w��9�I�|h
v��k�؏L� &Pp����EY�\�d�:�'k�l��7�3�� BF�(�uv���m��}Z>�}x� ���ri.4H��T;m=�;d�~"֤�O�rK}�u��~�)������]�z�-�
b���w�Z���.���&!:p���P�Ƈ��Ab��H�z�yu����o?���78�V�\��1�Q[l�a��.~u�ji�AC�����ld�k�vke��3��k�L��9?Z+e���瘅saul�6�t;���jV�n��	��cT��D�I/+[���h6i��i�Qm��eԘ����������u���m��e�w��N<7��Q	�,%��ɜsN�T���>:��(`���5�~έ���������3w2����g�xD=�%B�P��%�����A	�O���5���ҩ��
����$ySG�>v6�#D���� ���J�ת�rFOę%�u��ض�Xj�����刾�s��׮t��=�9��LmW eڍ������z���ֳ�!�8�����{r[� ����Mf�?F@g ?x��Pl-M�@�4�7� ��>��.����j曒�RuX8�T�}�m�B7u]/�+����.������kA &�]�	���B/ ���o+�i���V�n�v(�5����T�	K��K��3M�= �:���8���VE��zs�՞2P�z�Yv$���"o���>����iۓBUñޅ��M�\��c�.�� \/Y��~�}�4��k�{&)�S�!���V�1�Oȍ��g��{$�$���3�!g�i�bDVtW�|�a�Ƕ�IK�^)��/����j^�|9ID�7��ޮ��6d#���ggk���G6E��+}�9歫-!�(�Q�z���RB�k8��}vH�n����2�Z�)���Gz& ��S�������3��u�r��:��U.E�ಷh5��L�}�eG��Ҭ�7��#����>���&8��a��<�1,4|x�Ӈ�v��zA�@�]PK�'_r&���$���g��]�wlgÆC�;f�U~LI�Q�����*Mi����zF>{�/��˶�5��b%>BUW��Z��/���Ǻ�NȀ�T���"Gf�OlzM`�e"ʹq�@ld��}����%/�9��>�f���&k���Z/�㨲�^�)EϳVpu��fw���mSz۝��C�a�.(T�}�o��6V����4�	���Y��ⲱ�=&E���_o4�!�*���|��t(-�?ew��B ��zԅ�.!��� !0��s�:#�Ū�"������c��q#��_�[���C��o^M1"�Ճ��9��UXs�$Y@6�!6���Q�,ܙ�@Omn�K�������vRO@f<��	K��'{�r�����,>�0�7�����e3H%GI;��K�(�;�*v�}�'�VXzq��1�4B2B�;F.㑜T�V�Y����2�^��:��[64t�$'��٢�[�\����^�lp���A,��l&�5Q��+L�e�lG�=��t�{6�X�8�o������u��C}�s�I͇�͛��Ӓ.�c�\
o���QT��Gfx���ʢS5�Tl}Nhv�itmDx��m�d�C�a�b,�겂��%Vi���\�2<M,�6l��v˙�gxZ�ٶ�Sհ���)���Q�Z������]�����SVM>~���m&���>v���S۟��������95Yb�Y��O��L��=�G�����B"�����x,A���1u�3T�d�0$ރ�c�!�#GJq�y���<���d�
�����QQ!F��9�nv��A#OZ';G�(J�L�~�.۞��w��Q�����B�j�-Q��6���X�%�Ԍ��ZDq��1�V�vY�6��^��/�3&��������X4&-g�4ri�����>#|�W<n]h;�N��e�^�^��=��!@TF��y�d�#��R=<ǧ�"�'j}��ܷ��.D��=`�B�1W��?{���>8!J�f�{2~H(X[��^��s��#]�:]��:�;�Y�˷��: ���3��2���3����v����.��D�����0����ۙJ��l��}���0�TH��l���S��P���h�O��c�'
��y��bS���,a~��|���l�J��ϖ8��9�b���SH_ȹ#,J��H�q)a�NU%��P�k�B@Ȧ��o{�0(gԯ2u�� ��x[ӷb���a�Z���"�r� 
]ө��#�cgp�"(!v+��9j����/V�ΐ�v�ƈ��n_n��{��P5u��ɽ��?hW�^k�:f�&� 8g=]�������(�vD[ܽO�[�-z�W�r Ç$��n=1�t���;^���26ߚ��?�*ަ�xv[=d�p9xq��G'~�)QB�No]��;��	�����|'��[� �ך޺z����F�W�Wz��&�%�O����7�4 ��8tʮ���Y}Q�������؇�a��zM���%ȅg�p�B�� ��~g�*R|h��HOi�A��}��QͿn`Z�H��_^n��J�' L�P��ĻL=Dp%*wӄ%p�
���[j��H�^�ӟ�_Y�fk/߈�I#�鲻<D	��f��ۣ����G����}Q��5 D�o\dF Mp���3M��]!�1!<�9��?z���8���%yN_a����J����M����ss�r���*���w 1D%�8]�I��6S�Š+�`˝1w=8FvWG�y<0X�Жpc ��)$��
���Ji���q���ژG����k&���l�e��n�Fw�=���i699;8�whAV�$Ml�,���o]ޯN$�A���z1C
�����!�1�����,y�R�ҪV#Z+�����^`_�'4 ���z��aY6�M��E��ʷ[U�|�[�K���^�T~��i[�P�2.Ožѡ�/��«FUz��'z9n ���d�ziM�����0�� ��Q�5.S��F��nF���F�V8U}6M�6��`�������C���~(�y��t��������;19["��&��>���3��及�T�#Yߒ�j!n#s�����m�UslR
̻���}�G��?��h��V�3�ND=q�S�F��dp��eam{�	}/ކ'y=5���~�h{��������V�]��<��w�i&<+��8H٩v��Ʉ�%>�}��(x��F��g���e.�7��<C�jq���Y����±���]���?�驲׫?�OR��a"n���O{�й��2o(��;Q\�N���ae�,Nc�Z�^�/������U�kR>�"��l�p�79�\32i�f��#1 M�C��\�b-0�שoz����?�{b�n��t!� ��6V��H� ��IKl��aڟ��J_�]I��t��<K����ٶh���[)bm�^+��fJ���,� �m�IY�א�k�HF<u��/��mW5&Y(ҵ�OwS��dU��:�L��6T��76C_��!k����S�&��$bs�Ʈ�M�V�ߓh����$`���fAcr�FV�wG3ڲ�?ń�l�����ğ��
�� ,�V#Թ����8
�`~M7���=j�R����)=[^2$8c�u�G�#y]�П�M��x��'���I�>*i਽e��sR�bin�A�e�S�Z���\đ��
�u��r�R�l�t��<Ë�*Dfڨi�V�]A6�%��,SY2>�������)):Ż�x�ܦ��Nu&�n��$���e��rQ\�b�A<Ǿ�6�/�F�O�Pa$�+���g)�B�j�
����:[�
JƅZ0�����"j���U����㟫9�+���_�7N�ʶ,k�i�"g5�XtXa�/s�}5o𮟌���JF�r���� ����}z8VK�+�_��� �;Z�y�;����T��F�ǩ>�F�kᮎ�!/.ËM�~��"6�\Q7]`P�{җe&33�eS��:#�Z�����!4�V�* ����9�tze&*��u|��z+�W񎆡k-`ӓ:�������Swi�<x?��%�׭QmP(z����1yI.K�h6'_q�<���Y د��TA�q��.�фY�����2]>�U��j����nf�&��[0�t���x��E9Qy���1�G�r�~HٸmM��]����[�k����ʐe��jg�
}�����_.|jŦ�b�i	8a0g֒g�"Z�����o`Y���y8�" �����n(��D��ǀ��:L��QWV�u�9��ٰ���� �rz��!{�q�``Z����]]�iŻ�� �"[��}��D�nL�k�i�\��ˏ�קq��5Q�˥�#��,���JѪn�1�	��
����;����9�ʗo{Fe����y�<Q��0�Ȃ�dH��dme4bl��p]��,S��
��.���8@5���3B{��yT>��?�S�H`�x�p0.t�9u�e���t3O�lVGn�{M����.k�R� Wm������-�U��'�X�Lg`��1"{�g�]���cR�����l"G��fwD.���Q'�� �A�l?�.E���j��l*q� M#�\۾�?����@	�Z�@]�{#0�4�#7�8@��ʶLx]�MgZZ�R0!�L�u�l垢�����<N��(`�[,*�cR=(�&��x>&P֞z��9��2k��O�V�=���K�(�p���>��2W OZ �6�^�4ls��5���>���t�v�IЖT�	�x���O�95��\𝰞�9::'��oSj�$+�E<J�Wo ?)�#1d��Ɍ8�N�r7�]c��y��}�'����yO*Sw��ȮrA�+��w�J��yS��l*r�/�Qwd��mTO�w��`RT�8�Яy�m�8J��z�Ĵ�0��`��K�^c��Nhސ�Yx:M�X��S<���$Ж/:m�])��0�:���,��gh0��#��_)���Zj�f2j��ڙ����F��J��bb%�6G�W@{sM^7y0�?���e3�
݈�	4.�[S�������/*�7�+�W#l�>��ˡN�1����;��N�b���"��)�r��,*zq�ٹŁc^B�ǻ�@�]Eʭ��^��~�H�C}@�B����24������e��ceL�W?�3���%�Vc���7�e�Vq�d�d����1�Be�磒V�S:�[�& ր�O�_b���z�	�&^�+� iĻ�� ��'�V_�֢*4\�^ʼ��C�ys{�a�p��\h#/���Lt���e�s8�����x�.4��J�Uo̸te�IZ��JȐlmb`�;,������&�J�x̏��P{@�Ao�=�/�6��f�۴�W�
;��:�\{iyxw�ϥ�JL�3��8���5*�&݉�Ș�Z|˚���p5�����K?� Lģ(h��A7D�}i� �Qy�	#�@
����~�'C�al�߲N�4�(}�G�~颐�3�M��[15��/[�-*��z�c���ƹ��������φĵ$�v}2I?��w?�1� �c9q.�)�ҕ#��е�R���\��BG�\��V9�֎?՞��Vի}s&�X<�ē�b�Je�Z�)O>M���=m�M!;��}17��v�,�QE�Y!B8�}1����A�h����V�z�8v�GV�A �;�?�=Iy����-�~m�uJ��,2A�#���xP�|`�F.{{��<����l�!n�Ө�M��Pya:�[�MS�RF)��>B`�QU�A.K���e�)D��q��2�|���}�U����b�:�n���,��C����������M���w�,�*���.>��К7���vb+;�8�10Y�o@��c����lnζ�9�6�(B�͹��'�y������@V����(ZP�I�H��n���no�bϺ�u7�F��k`v�#$�H�+T���ѿ{���>�u��K��N@�p"FU_�u�{����2m���~;��;#ui�b���S���2l/x>��S\}���#�N[�ŕ5i#T�{����ӗ����g��HBeƠ;0O��O�q��*8�����͒�$��55=Ru�;g'E�")�7���8R�/>�3u�D��w3��lE	������I8&M��n<]��f�m����V@sL����v��sg��y���*o��f�6�k�D����Ņ����[��P��C���+�fW	A�����^(�8��徐+w۴u3R�.C�|��)�:~0��k�!wȥЫ ��H8ҵ�� ��f�m���g	�G���ۅ�C0TT�����|���⏂�N�
��e����%bDI�QD���
&*AA�Ɓ1��qF��g�᥹���A��x�ĩA�V#���3�P��k�%��:�~�8�N������yc�x�(4�9P\{�^�V!�C�V�~���)�g����a�@<�w8����Ѷ2o�c*��bXo��3o��㜉l�5�8��1i��ܣ	�|hgV�;���z���L��9��������궆�XHWN!�����@}��G�, �n7�x$���B��A�Gԓy�ŋ
hUU�BwT��?�� j�ޢv�κv�pEjm#�K�JC�l�o�i$�k �W�O�_��(cAА[ݣM%�,��!1��	���m�d����&�E ����"����.��
�L�܇�b���R
����� �y��	/�\%���6�E���1M�[:�Oٔf�R�I�JnI�z��n`�0{�(CZM��g*Է��`/Zq�������<���:�
E��b�W�G���6�Vu����{��p���d���\���WI�vb8�g��P��[�u�~ec�h�]MtJ��n��:����E6��Bjtn�ǟ�ʕn�)�/j仞pa}Y���ݫEGԋO~�d×��x�`�pU)���
�}�����%��M�:�P#(HSYۖ�g�0�p��u��!p�`��}/.�$;Po����)9o�l-N��,����9�FR �v	^� ��`������cpG�<oԱ�a!�ъ+mH�ͥ�C艻���"�=�UME7��P����P���g�e�7V���ю���?�p����f���I���:<���Gq���:�FA`�˃A�ȅ�i�Ʒ)�������p������˔^_�|��/��x�쭞�';f)74�#]��1c��Ԩ�������ȕ�;��A���@Ǿ������J��1˴qUKu�U��X�8U�*���=�J���U����n/e���)���no�|�2,�Y�(|@9�㘺rYhTQK���l=B/:s���ͪU
C�ƶ��+��ΔԗQ_�r��)Cs=v�i�@����$�z	<����˹E�����լ��:�/�P^�6MLgxڶ8�QR-<�3������(��o.ײ�"8�����X���4�m_��ȱ���f�2ѫE�뛲=o����!��ǅ'K4D�Ѷ���^9y�R>Y�@i~�,�����GF�R-�u�|�G�]��S�d⶜��+QƁ��㞃�J�0	����$��.�w�7��Y6��ⱍ<s�i�4�z�h}��i�M�PsZ-�e����v:�Ӽ_���9�K7i��0\�#!`ٹ�Q�l1DS�y>�Qˑ^�t���8����5%zL�h�1��!�'w6bM0���S���t���.Bں�*ֻ�I��
�5=gB�3XD�u�?�^�旷=/x���^��3�۫��5c]L��g}Q�e=L��8��2ͪQ��Z��Z˲>�So�(U#��r�F�H���6^�yI���D9��T��0~�E�Z"퉰���������2��Fei����/���k��6!HGV���h�%�/�Ӵ	설��_%?yP��{VY�=��M�O������
o���Qvr�)Ⱦ�F򔞨��Ir��w�GJ�N~>V^ۆ_�_e��Ժ���M��ޢ݀�۝;Aͪ�Z(77�f��k�.��,�pX��,r���Ҭ���NO��O�&� ��Ի����,����,)���q^�<�S�a1����q��8���!Hp8�Xl���<��A�cT��"m�ƣ�r���i����L��F�8x����O@�Ja_����!�A\H�!�	��䤢��[�ٷ��b����DIN��]IC]<�{gZ�uܩ�pc��!��7�a���-�^w�=�=����/H��X-�ضX�"yOZĞ���X��K��'�L��~k��9�p��w!n���M�ZCb�g���D�@:.���_�Gi`�m��(\ئE�%sl�K*`ͱC�J\��v�lfߔ�p2��7O<t��V�[Q}i�h�V-1ՙ`?����$4��� W?�#��m�9�W��8��KEL��Շ��a�*D]�@�Ctn}uj/��%�%�]���%�g�P�]��}bO�V��)>Ð�Q����G���cO�A�=!6���u���q�2����6ʓ�6��B-��J�k'�<��a�c˝�c;��8:9t�����W�<\L�T��]99��3t9�����c͟��K1�l���IҐ}�箳��tBQ����3��	z����=d��/�(�J�eL	��g�y�|bɞ���V��%vRe ?p.�}9��E9�����Կ�1�{�4�ս�lP�G��ǝ&3��Yl�Y�|7PX�rCoQJ��s�@G���(>
�P���>n]��Vm%�S�Z�`We�N�T�h|S��������*\;�*T��>t�V����=�&K{�N��ʲo��X&�OϺ �r�g�XN�~�獅[9��b���ș2�CsWzA�.��a\�׽n��z�
w?�pk���C|�=�XÿF�z�r���%+�*�U����/G�-���x�쵘X�b�Al�wS��CH˓�!�z÷��"��� h��EJĽB��5y��}�I�?���	���q~K��ɳ�4�9G�X��߈1,ȿ�~at F������Yq�a���1T�]�N�^�' �Bu�J\� �zI
?�$g�ڬ���e6\㳥)�������.j��]�ɶ��cW��5QS�i��-���\V�?���_���7x�?A9�4��ʀ�e{p�64~��M�>:=�8��Α�%�S���o�)1�󑞤��xi0�0�HYNP��ڵ�K4�q���Ol�+ʷ`B�����s���Cᑮ���7mo�NҸ�3���E1�M,2n�on"��}R�fh�D"���k���5N�D�7�2�.�g��*/GJ=$�x��{R�L��
,�V	�y�Q���뾇���Cq]E��Ƭg������>�AY�`j�?!�<���G����44ay����5�z�f�:2`�i�5���@ioǣ0�cS(�`���(���9ƿ�ow�M�~��Ƚw��_'\���D�s�?�a��g�w�u:*\��ܧE-<�`�%)� g0�C6�n���MQ�ƩH�~��4驪�����t����SO�ݖ<��8�IR�T��om �VQ4BV4��|�f�c��q/��nGa�P���iVŖ�~�M��A���\f�!L�A#���
�=#�@2Qo~Լ�����^ʼؾ=�WO>���2��<i��� P{�s~{m�'��& &������H1�0`5����x�|���.-Otk�`7_E?`d���Uςإ'���l|�Pj3���_����FZB�d/{��l�wS�Ga9���(|�y��7&3����o�֝�v�lh�ቔ���Y��b���ʘ��]��1�E�+ZP"��"��%j��#磾�g���	6�ݾ�M�8b.�ݘ(K8���F ���[�.��r��y��;���I-Mz�&I����س�#ߦ#̡�N�((�@���lt�{\p���	x=r����H�uk�
^�v������rۨA������!�!
�dtw�9W-��N�l�!�{g[$G)͸N����n���M�=|��Y��Qd�_�?w�X��cfK��  ��g��L�����n؁�;ܳN�9����!�]�L<��iM�a���B=G����'y�B+� ���_�@\����3����?���	n^A�q��~=���\,u��c������Y �7�E���S۫Ǜ/����߯���ÿo�w�MS���A���dK���{"���"�6Ysn�Qp+q4(�������vYwr�E���ӇIɏ�����<q<����n�����z&(5ء� ,��BY������IN���0�<�9�3#ɰN���܊���GJ�.�%`G�w(.J���h�(�}V�ޒl�A��������>�s\�ņȰ3���&��k(5wq��\�����������%��yQ}��<.����j�t���N�PL��LJ���y��oEZ�3��R�x3��D�����w�-&�ڝ��'�,U^d���#SP�l�I_@�����?��-��ث�`�0lg��s����,-�,()=f7)�c3'�X���?*�S������o��~�<m�� tZ�_�S}F
~���DES�J����k��`Ϣ��F����P�v�3
$o~�qh_e����C�(H^t��e'�ȑh�oK�c◌P��%�����?�c}2��TN�Ō�oEBw\��%��/�M4?=R�o0��żX[��e�����$�
>�g�������#|6���o�We��+�yH�c5Pr͛äݗ�1�Z�G�$e�.2�_n�Ԓ6�8&�$M����~�H�1�B}Gq}R/���A҅G��2v�_�GA���Iǧ�r���d)����@�!ܘ�-��W0�O�(1��,���+l���[�Zi�j
�ە�7���&��M�?���`���r���?^�H�}�����y�������cm��iaw,J$;
�L����+�z�,�u7�� �?]ς�V����l�_�����O���N;l	���~����K�џ���҈�Y���2���z�tIv��2I^�_yU"� ��fD�I������0�l"5�����5�-�~���ZD%���'��p^H�tܰP�U�	�Y���#�lAƠ+��?�y�9s�5�:�S_�WiGΉ���t�?k��o"�.r�v�& FrL.M{Z��W���f! ;��T[��Qg����L?>�/��JB�0h���2���G���3��̚.kpԴ�����k��W����	�|�˕��2[v������5�T�"t�tmb���ǂ9�|~�璞\3$T�a�.�����-��6(%�A� �6I�=���dЀ���mC�S���ל�m����*D°]r��UG�k��ľ��2�X�:�R��#��|y����3TP;|��.�u�U�^�/!D��?Q�>7�a{bet-�tI�L��(��M��'����$6m�i����G�n� 8ޜLH���(a��J�8pW���7��S@�NZly���o�Goׯ�* x��0��썙��88���u~Z�F���@��p�Л(s#8�'��N��?�(��x�P���!������ֿ���~(N��Ј
KiG�hAz��q�u�w�^��ք�qm��v��Z�TQsژ
��'Y5��w�\
\�va�y�b�jk�l���2l��?-���7�R�A�h;Ze��:.�L�C��f!��]�M�c�,T���4��Wa����N������W qލ������ܥ�xP�政5"lM��M�'Г�����g��9;̧��H�C0����*���0���4f�n���
����Dɛv��1��XH!��h���=���7�)ɜս/M�!$��Lf]�j"kQ�� ]&����J)�>�9>�o)�Chq�?H'�K+� �6�|b;m��������7F4Ƨ|{�&n�8�,�E��S�O�>U*�yn��QV�KW��$byDj�F�%R�e#�)T��Qz��DĊw�����ӊ|[-��S/����x���+j����n��oUDD4����ɻ������	�^Ǹ&7�	\a&��0�*a_�nB&�_`V�k��7dv���Ou U���J����el������*@��9�>�u�3Ҳ���F��p�mJvG�!&��X�ʇ��x챒@V(0�xey6�@�$���(�Qo9|�'Y������#9�ƖGS0�\�'g����lb�e
�+.�:	|T��MG�ȊB�4���w�VV�+��G�mmGp�n�O�%�Q��;
���KQs�|�5��i��T����&VJ��V� X	 _s,�Y�=�`V�{xǮ��f���uzZ*<�B�Q/εgڸ�m���m�ƥ��Dg�Ҟc���/�����X+)���7�_<Q�N�2����H�J6���y�r��c2�Iò��-��^�CMK�m�)�TA�J���&��{��<E�pFY��1�`���ʐ3|�K��!5�8�+>��:�xhE,�jmG����B&��L���X���V;`���d{(|!Ĥ�%�����>卋nABcY�dg���������A=X��g�	�%\��3��6�u5����@���AW�U%'E��!y]�b��dV(�0/2�u�},'�i�G�5�Q��X;tOFR�;�i���2�V�<�?�Wo���A��>�o/��q����|{����q㋅_t�&���F���,+ԋ͇�p]16�|`��)u��Y1hި�� ���W�pc����ګ���n7��$G�J	�����P�͆���l��Sk����k Ԏ���b}l����}R�N���sj�qɭx�Uu/-{3~�!d1����j�.���Eũ�v�vv�q�ҷ)'!���X�[�(��`jk�(-~�N�cW�Kʢ�p�O���S����}V��M��@�;�̊j4XF�s�З#���E27�F�ĲIt����7?����O��C�K�*����q����#�~z�$�g�?�F�]��^�ȕ�$�����[9x˛U���ֺ"�q8����7�[R{�c�B$w��%C5:܂�*��!�$(̆ �h�h�+�.j��&�!E��gf�gB"��/��R��Qa�I&�گɄ��[D�olz[b�zW��U^P��8�O����+���L�كt?w�n<#ABjhsѾ2���?����Mbv��4Ѐ����H6�]̬���	1b��"r��smIy����
O&�)]���`P��t�N����-�Xlɷm��r?�x�/�����K����_D��,����nƱA��_le���*�� ���.a�F���p6�|�%w�yIx�V[�m(SA��2�a8��܃>PďV�C}���;�	�tf�q2�r��2Bե#��oE`��H�A�Ԣ�
��2)0#F����:�^���|��.���F �[����3wG�惑ϲ4N
Uy	^M-��ט^�Q��o�Qޱ'���'��D8��#�p� ؈�hp�2��
��w�f��:��f�{�R��{{�H�GP5󪢀3%"Sٓ]� Nd����7	�!�w׹�tOq�t>%�	F�)������.!`����"�?��_LS't��vފZ�� ��r]�z�&�Z%[J@��Gf�ԟ�/PT
⽬UD��E1�,�t��SS��!�5�|頽��;�t�f����C@��N`g�3�B���"]�>�Q�*���pd��2���1�v���rG����f�F�c�d�M�S�G��l4�ԫ����R1��j���Yj)q�#��H��0D�-;�y�� �7��?�R��N�IB
�R�ՕFOӒ(0�?鲗��:�Wu,����;�$2~��Ֆ��iQ�+�ـWYb��Gx�L��Y�	�-ڻ��>v�Y�;�i{��O�u[��ʓ����~��7��}�ze�T������'������z��9/?���Rn7�y���R�=��$P^�8���8�̧��(�� ����Y��K�n�m��`V�Ѐ�׾Z�U�g��AN��H.9�Vz��r�0j���>	@ ��*�7՜�v�k��5!NCe���Vw6"ް��3� �G��C]��uB�s�������̇�_t%$
v�2����U
��"����X��
�9���q�ٰ�Gc)'&���ļ^Ϫ-��6?��1b|����"������_,�-���D���T#�x���I�G�F2x�a<�N6d�{q�7<��I�՚>I����|��R�E��?�-�{���c��UD���mJ@��j֔ ~������GKsڑӪ-�Gi�������{������ �r�A�?f?��q#��'�;	󓱎�BY13f���9	�׳�
��l��G5d&=\q���R���a�*�
��&�����I�J����������`���!3�a�)�~��+���%5s;�L��YU���/_=l�@[`��`��a_���F�t��ő�,��"P㉉�p{��J��tg��Ò�~ ,�[������T�n��rBU��>�{K Ų�
��8 ekP�
G�nI�ܟ��6Lrs����ܧ�|��$��0,mx��m7xsW�.�G ��s��Xo��lWvQلW�&�bW衛;�:�D�s^��p��|��8�D����Z��F�:"II���-�u��֟�e�-�wP.��e6��P�V%��3�ƚ�M�����,�N����aB>�����2H����2I��v��xw��0c�?��C�p_z�q&R��C</�
T��s�1���O:n.m�
7�d��|A�%齾U��w8���D�t3Ծ�n�fp�)"nI�b���=L�Bg�+�>&G��x]){	�� Jھ�V쀆�{�6j*VV�\��|��j�[�iNNk�?�y����y��+RSY�����D{b����6�m��
b���&�{�>��J0�QԻV�j5v�1�a��X�i_G.�v+y�"<\@��=`�e�	� �nD��nA�_��ʐK�g�<k��ۖo+��<Axmq�s4T�Jo�.�cZEYm\�0��,�\Y=����.3�Nmh�A�I�c����2�緝`�=�6�f��U�oH�g]a^�bG��g��?��*f>N���~ö�$0xJmHC���M%���i��w��6C� �P����Z���7�<��/��cX�V���/�7Z������$>ݽ����ۘP�H����Y��;��s�y��1����2�iƆ��H}��p����|Vr@
�E����γ`�g�7#����#gh�jěQ�$�_�����>G�A�<C�!�)����fq��Z�:Qx���[�ZV�`N�~%	�/Tf�n%
�M8��z\�r�S��y�B8�Q4�?�/C���ZS���	��i��6�5�D�#/�ܓ�8����f0����OP \�������ݩf�8Dn3f�<V��w������z0�t8asz{jz�����3jYWVĲ��Y���#��-���FkAO��$���9n�G�S�ҿ����!.�G~#/�,_O%ԁ��3��R�"�f��R�`�th�d9g;k:�r��������`�,�e����-GM�{D�����OW #;6m- O)���ߧx�m�nY/��V�i:�A��	����B`11�Z�Ů���ց¢�B��ԆT���T"'sʓ��J��+h,���q\o)����@���XN���!��P�<[�u��q�4*����)�'z�yW����ׂ�EGo�ɡ	~�Mr�b�%�8����)���TD��d�g�K���9#�X]��(0��n�[��y-Og�1�ՊlbNy_�IU�I�R5zh��:1�����ߧ��ewV8�x;(m��$�~�)�o_T4���L��<3{�����GK���8D��<�T U��{.��P�B�!0''ǰ�	��v/0���)�H\VZ�ꮽ�Rm������Y��i"�R����Qo8��X��]mʭc�?v�T�����e��m�eY�҆3���1}Z�+�aeN6�-|��.g���j�����Y�b�9۶ִ_�b�_,���S�lbݐ�M��^Y��>�Z����*'F�]�nDΚ9q���;W�� ������JH�0���=�>%u������ �)�t'o�׀�cK����o�:R����6�-��8 ���a�C+φ�J< 0V(J�ЎV^\�f���Z�-�T@�����~�c�K�ppJ�>qm���A^qx����vG����z�V[^lM�ژ�d��!�c��x�L��@�⪉��q}Y�牔dx����慯��b'��1�G[fI�Gff�&�Ih�m.��MPb7�h�_���&��ٴl���X�}!Fl�je�T�}���)Nv(�V�(2@�"��x�NZ��.*��'�3L_������\,�%FJu/���$��B�����޴�Y�-�p�;�r�/���P��bM4��0�{}�f@������k��k�y�4s&��b���VmU�Q��}���k?rr0nܒ�U��]C���m)Q5L���
v�Ўg�HMަZ�#��K��?�0b;�P�`�K�����e �s�R���ߔb��(���IK%V����1��������r��h� :�3()�\F��6|2+��C��I4\������ڮ���~� iL+�a%�,�;'������Nv��h-3��`qjd@$�'��l�@Y�:^4���l �!{9J)��I�
]B��r���&���lS<{MԌ���0�Y.fs��j��;��܋�14R�,�������/�-�������Vq��L�e�l���chr��.Q�>����H�|4�_�:�:����A����4��Q�-�M�/�J0#�L��4D1{�R�o�7�W���A�`���H;lIK򿁍����X��������u�~X���8�J�1K�\cC���3�٣�N#�ӡ�����6�Gb�ԃ�")p��Q9L������#��J�Ҫm��ȺP-x�@���k.������/�~G8���ߡ:\H���g \�T���m0H7�8���8��#䬫�����8��*����I�k5���u��r���-� v�-p��a�G[ZX�LF~�?'U����r�)w�9���5����UG��{ِbZD����,����gr�td�`bxp�-�%p��B�7؉o���*�Y���0�9�4Ʃ�t�U8�%e�o�������� tˑ:�{L�x;�?I�8���x,!O,�55>}Ms��'Ƣ�(��%��<,�{�YF�ʔky�θ�SJ<�-���o;���e_��3c4��;�G�z(��o�p��f���C��`�B��ￆ3�n�OE�H�h��T��{��.�qE���hx�Z.���GVr���}�=�Nf$z.��ػ�ڗ����9�w��֚V�}����������S��!gӼ�͞�T��Z�ꋞՁԏ�������*/㬮oOA���՞�J��0�p�k�k���f�v��D=V���d�Cu�@�	�7� �
�얦��4�S����� '���p�i��y�go%�(W���&��Ϯ�?�|���p���#����Dۡ��E񒠔�_���a,��LY�m�SV��,*G��p��~��E��+#sZ���I��lY�l�]����R���lP�C���Uǐ�<,m��1�9#,��4_�� �B!��}�e��m�����fd���Yڈs>b
V�%[��R����ķM�����s�م!��@Y6K���[��&4��x�H'ʤ��s_�E��>1$x��+��ć_����s�_�/�ʁPI����%ͭ��Ge�?��U]}��;<��G�i��I������i0�dq�w�O	�t%� Po^%Sp,��p�G}�jM��9Val�+��I�	z�dz]�=k\sC�����C�G)���5��7���$Z&u&R���0��e3�2�,��w!���@ܭ�>�!͡���P9G���~tb��Wϙ�ߣ��?Uk }ذ Z�[C�����η�`�0J���%%P�c�����OƢ����0�K�ߠHt�q��0�JTr�~k	�����+�"�3ytC��=����9s�եl�7�W���Y���8�Z���K�`�^��T�@��xYIς�E߭(�&����E��Y��Wc�m���)�i.=�	�*�݈��g6�k�{�V�x�m{e�egi����ci�+G��I�s
�?,�;5z���9\�O�3�y���Ƅ�n�q���G^m&HN���W�-��>��R��{�K�s�`�y8[�>܍�L� �Xlf�3�7Y�ڽ�jY_�"��F�zGȫ5��
6w��9`���:@���5lVz�'y	 9��6R�Q1u&��+��r��HC��*�M?�L�v��������$:�|Z���u�E"�0��S���̮��۽�ם�Ѱ��xc��:�=0>�5��<�c���x&�=��߲֏�]A���D�,.�ʃ���3��Q�T�V~'��G���D�:7�;����_�g3�[�K(�U{zކ@Ū|��"���yC��ѼX�\��g�b�������H��Y .k�a�;�ې��H^����|��� �x0d��9KЖd���+aS�D�)�*b��AR�9�a�Ϋ,[$�o�RIʃ'N�2Ep$*	��a$��h@s �iB��ߤ�J6R�ov~�8��zM�N�P>��0j 4���Ԍ/U�7�y].$�2)co��G&�kY�I��ߎ��+|D�g��	i	n��5�de��H�G\醊F� cٽ�*D���ҁȘ�񤥃��=��0��}rǔmY���A9E�+�_V��-��h�|f%��}�R���R�cR� )�12*ܓ�9���8V�P�>�> �8x��"�R�"��!<�-S��F
���$�;H���s��a VA����%\g���'��&��H�> 2~�����>�w�}.J4\C� ��n1YLyʖ;� ��VAh��]3|꧘�(�����^ �-��֍�\�I�B���=_�ɷ_4{J��I��xd-1�y�����pX��e�J�$
�)	
g\���#�6$����XYGi�ǟ�|z\���'���m��|��C͜�������<�؁�v(T4��B}i������$��������|~�a]��X�grV|�.˶�V�g�Ԫ������yO�.��RH�(Cu?��(�Yf�.q�����T�st
7q-��pg�)s����*0;�[ބ�\&y�B%悺?Z�_��%���ŷ�\�rd�=�J�π�@�����P^��nK��u1׮^S�^)?��~\�е�Y�yt�\��0��2�rP�Ӵ��LY��%�\��M�HW	l�R4c��'y���[Y�b5(����)VY������w�S��iQ�*�S���V�҃�l�����
E�"���	����K���5��L��?J~�h*s��[���u�dn�M0���GAp���`�`p���=`n�It�	��3����!E���+t�_'�S���k�Σ'$�"b��o�t'k�������9�Ecq�Q/rX��S�뜤U�VSOfZ�\��<�Eʻӵ7�&�y�*h+�Dr�U6_�L��j��U��O�H�=�������x���s5�����v'��Lё�T��Wyċ�|W���8�ѣ���X����y�X�K��v��9��p#���y�E�����?�%���C5l��Դ���&��p�Ķ��4�<@��`���Y�H��� 4��K(yK9Y��"*��[]4���6x�Q9R2�_�VD��{��+]t�*y����o�Z�s#��ߢ��w�r���Ϛ����XI��Y�Z:1���rX9�p�u�-Z}.$O�+�4}?s������I�S�W1��d�C�=m��tQ9�U���%\]ލeB!|D1�|;��$�)�Ԣ8����,��_��6Rܘ�"=��`T�C����Dȥr���jf��I�N�B4F����������b:y=i�[#���o�m���W_�`,k͔��S���8Xru� �loԖ'Vx�[��d��ڔ~�y�wFk���\�P,ȝ����ٽ�L�f9��5a�# #�e���҆ab| k������[��4��7yNؚ̡�l��H��?HJ�r/5�ͅN&W��t
Cõc�qh�t0�-�=h����2B9�����5�zNp���p��g�/�:1}�'�$nW�pO��h�g]%"�K됈��Q$�>��B�l�3i�j�|�O�;�b늰�$�*�ݵ�\`�I��QZ�����\��Ԝ'B�eS��TÒm
����ٚ�Y�[�����Y�5�B�\Vj�CN���oD�#, ��`�H��W���@F���F��V�<qnmܝn^dU��z&�
�w�xG��N_��.��x���0p��	�_&@��'--�+��Q!7X(Q���3/�_����peR�y/�f��n	�(i*���]׉���SR8�'��*��FC �D�  v�g��D�<�PT�.���^��m�Xe��Qu�3!�BrY��Xu-@t',���`�i�b�[aеv����=��$�Ϳ�x
yB6��TL��M���@�G<!E�U�����L9f)s�]�ڻJ�qm�7&��#��h�bL�|尞��m���Ս�8��{rJ�{T�1��X�����s[����-zX%����
#!Ā�����\�訌��FY������>`��HJ�"+z`~�o+�!}�]�����l:O>�$pGs��oz�q�⯉�L���p��۸�=�aa�-� ���w������}�+�4mt�	HRu��(�2�<$C��������B��h�M;xA�"ˢ�����J�T٧����u����L��{�_�]Ɋ�\�_ ���q�p6?�k`��U�
r¶�t����� ]8<M��}�#��I^l�&v��O�Hq����~(�C�|N	q�uIg,Bgh�ȁ�	�Q�v3�������R�^�x[�[�p����Q[�M�t��S�~�!�A�,��5-Դ��K^ZpY��Z����W���O�����I�r7��Z���l �7KȰ��\��\���ч��=��ב�| O��N� ��sv��x�� ��sZ��Ä�i���J��jv8��6��0�,:��צ9xT�<����*jm��g@�%�J�yh��A�s���@=x-�n�G��㞁-N-��V����rN)m v:��^�ԱV ���;L<#�AI����Ү��E� �s;!ŭW����T<�
X�ˑ�_�������X��yZ��l";�0Y�"�9��&��V�GW�)`��:X?\vxZà&}��S���F 
UA�ْ#�bQ1'/.�[��9��C�6&j��V!��tK���r�/�e*sw�+�>z��� >��N�[�*�+�6�X����D�v57�'�6����8��y�[�8Gt�,��r��&�O}n�r�9�+3��eGH��B��h@.��%��s����=�:4��$��:�bw�@��������V�ZKe��� 9<]�2��4"��Q'G ���')��a���5���q�o��xDS�F�p�x������Z�ʔy ���׉�������hw������� ����m������ch=� ���A]Jsa��.�~�n�󐍁nd`��Ơ�[2�W3Q3�JF��|��J����Z'���}bH H]k�b� �����2[V�	��V�&k��D�`׸��u6+�U�
���� �6-:VM��
*ՓY[mKmRJz���öz�Be�_�g���e�\��|�8�rr��[Em�-:mva>��k�Hb=V٠e�.
�.P�@���=�i���R Q��uG�KMV^�0��# ՚É�CK�+�ۜ�瀇T5Yz�z����U��t�J�x������'�[ZI[���h�K��o����]oM���m�/��}:̇T� �	�S.��"�r\j���\�A	���Yʓ�I��pBQVN�Uw�;x�Y�X�t�z��A�/�3�K�]a\��H�h��O�4�29#�d�� +������T,����7H߽�[+u�-�	P�P��Ǧ��6n��,�����F���˸��'A l0���IR�H2��!�kk��ۙ>���Z׶�"V�+i�g����A������{'��F�ѯ���̭��oOJ�̚e]�ط[�>��6D�՛�Us�D��:��^�j��!�8��?��I�w�U�t36�����䂉�s��a�iJA���vl��Lү����3=ܚ䳡=az�4V7�T���(�������$??��)d�V��@wi�(K�jDF�uCP�qy��;%R%)�(�K�H�%��F����?ל�ك�0����1d��s$+�a0��
9C}[���|�)�����ϻ�&�EE�/��/�Ec�}�c�|go�&"WN{�M)�0�AQ�2�i��d?$'�>�F5y*�p�	�&��v�����7N2C ��������|�^�ſ���A�s��C_,CD��Ғ���6��%_n�	&ce;�tN�R�������ݘ3U��|滈��ћY��^b����H�oX���y^�~V�S���TB��Ǡ�	f�3{�w�ץ���g�qU	���ڈz=�֎/����.�r�:`bG��3��ly����O)��o,�S0�/O�L��?�K�{J��¶GR���i�w�#���]��F&?,���B�!d W7n[۝6�p����ie���-��@��'�FZ3������~�{&���n׆��N�{�caľ	�<��$����yʯ�{i"����_�rT;?�řh����gm��E@$<"否�P@�;:���-eN#�z�� ��/ﴤص�y������hD_]����L^Ge�9EZ��4�pG@��ʘfO��⥀+Bɨ��bs{�tQog;^'�l�y5(0��-4�n��}�R��W�U.v�Y�����^�w��MUA����e���;#Ur�~�Ѽ����(q��RMȹ�����t���Y�+��*N�D�
SWV�=o5Q�w|��
rM�Of�%0���u� �C5-�x�J��t�YVU�u(E��/�W���ƆQ��͋aA�DӔ��U�̼)�Eu%]�%m����Ēb{[�f��Z��yB�6"g��H|#�'V/�����;�BmDA�/��x��aW�mDa��?-���0EϜ�nY@i<�7�	�k�R_��]T�r6�gѷn��RdN�Ap|�r�E}w�7��U�`�;xo퓜�.���@�ŔR)AB����Q���e��V��A"�X����`HPک����J>ܟl�p�T'���
����ݽh��V�u��_��-wx[d�ί1C0̘�LȠ�M^��u��1���q�	�{G��C(l�NR��G>�#k��[�a)�Zt��=�C��TYP���MCf�>)EG�Ȯe��ۙ�ɻ�������ҳo��s��{M _����M[�/MI�ڇ��c��R��P�(�h)�l�D��{������D�o8 ;��>�簹��K�{�v�D
�.NO}|�kC].��KzRS�� ��Q��]&�x�DV���`Zyb �FP����;y`�����9%aMy�$��Q�q%��v� &6Wb^Hv��7�Tu�K�~�U�ʒ��8iA�N����y ��%�և��>3��_���һV�^�K � �R�C��T��=�g�B?ӕJi�g����2�=���۵��1:Z�U'jț� M���L�B�5ۇ�=ά�n3��9NO��a퐈�@�솩���HX����BΉ"�����]�r��6�XiO��1�k���I�B6a�҄
���&�d0�슦���m+a_�e�7(�wV��Cr�nM1���~93X���	<!�(�
�A4# f�����w�h��h����xG�������-�+r�Cʌ�ͼER��2����!yl�|���f.?��|~����3H�^lf� �&����3#c�E�f�l~��πqX�<FG8�_���j���{��!���u/kl�K|��QQ��{%���S9���\'� ~ŌP������͝KJ��N?�!t>��)L�2o�J����=)Hb��,������,-����u�+�r�U�H.���8(�]��M�]�OL{�1rP!����~ޏ�)i�U�"mY�lX�{��$�3d�T�o!~˘���[f�O��ρZ���h}�~��!rj���F��HNh~0�CgZB�=6����D��2�VM
8Oj	�{�����n��&73.+s� q�qRJ�!�tfo�| P�V�6��]�yPC�Bڶ��jnxO5_A��?fP�=r�7�q��������~<ώB!��5�
�SO\]�#�Z�~vT���\�x���S1Y���&�Y�	�),0V��A�z��~���$���:�Ő�X��<�tbp�1$N8��{q�z��w�9��X��3����FV�F��/���Bow��{������TN��Q�j݈���Hp(wPF