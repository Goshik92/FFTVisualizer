��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M��*����g#φ'����T��6%.^f��8{�^v�wK�T��fAN(.�oC�Yt���Ao�>���� �h�*��9礩[s�Tj˧��Y���oG� �'!�D!�#S��E3@b����}��(��ѣԿ���:+��rYV��;��6��!�iG�{#�Rݕ_����JkK�ݽ4\�(��.*�[{��+����3J��� ���J�S��pթ�`�]JX��X(EЊ"����sZ�Бx���
�Bo\Q�t�����vw�ջW����ccσ�*^���%l���N�rd�!����Z�q0G�nRu�4Q� ���������㜕�f{$u�6v���9,(�l�Sj�[V�����&�F��=��{+��T��ca�ZR  �9�%s��E�ME�4�����Տ�ϛ]�䛝'����;��MmFM)څ�+H%��1�r��ۼ�l����<�K���35�I���wp4:c�*�׻��C��
�i84J�:츈Hq�Z��B씩�'�JD��4�K{3�g���?P���C(������� K��8��##M���Y以��5�DU��j�o�K�ِ@[��{d��otТ�q>h�s��i�e�֡��4m�����-�Ҙ��9g�`e��-�^���x�w9;{���QU������2�Y���^#�I� ���G`7�Rx`�k���]ω�o\����}��(��ɰbUޖ$��y�i���XCJe_E}��ƅ��F���Mn�d�]�E6)�^��;���X�Ǒ͖O�?u��+�
�C^~Q3&B�tA����\�ݏ\�By�hL����i��4�x�K<%[!�&�L#vZ/�6��H])k�s`R8NRL��N[��i���/p��n��JF@������o��X��d��;��G��wi"��CbK�/75��(�pĆ�N}�W����u>���k��%�ٸ�Ui6��Wy�!w��g̸��d24s��,�^v7���:�W���m��k0�E����?�'��>��!��o�N6�(��k8����"��A���0�R�Fh�|V�hfG�\U�H+�iȤ�V��~��rQQ��~W.{k���GT�.��zi�h��9J&dAFH��r�P�b
��R��tX�m� &�s8�MP��uP���Vj�/��w���<�ٍ�D�5��M�*�o�>Y�� G)퇘��>�:>��"��ۿQH#Sj?LnlC��b�u��7[��ו<K�T8p[��
����*�!�lnv�:>Â>����3)s]��#��6E1}ŵ���?]^��q�R�s_ۆ��Id���5tE/굛ĸ�w�/����]�A!?j4cJ�����2��aF	�n��dE�4a�����`P����x	z�Q��T.�W3M����G�"��$V��F�քr����M[äth���u���)�n�ϋ��a��q)3���,514r{�\������D
�6�s�>����ٻ������{�T[|��V�/����H���m��Gβ�����N�ժBL�c >"�� >�@�8��Y�z��:`te=O�lFr=�W�첀���%c��8�:�OG9ԟ�!��)er�(��g���\��l/��m�V�L�n-O	�t�]`�U���
�w/�	�,�	F�U܇i��:_��*���WO3����6�~{z�l��}+ ��W!���Lv$kF�y^D!l�ҭ��E6���:<��,r@0�귆��d��Ûڸ�Mi�[�����t�<_�����}�^�n�/�T�b���br0A��a�p�׫�z~��""5�B�\�� jB�m݊�����k�?>k�����H��*9A�tl
^���{�u����U�]������t���^ B�٥�,�N���+«-)����3�WĎA���9�cU~ߎm
L/�B�(9	�m�W'O�����p�>���tԑ��(� 1?1�Uڨ�u?�G��Nͣ�i�K��{�+�s3��w�9t����ۺ�/�ߦN]&"��K�-���ճ �e������LRm(CKK�I�A�\"X{�{Wb�`e.���9�:����ES^S�$��IZ8��P(4���e�K�ʡ���i�
�uy9*k�ph#ڵ�d}yGK��Uxyy1�m����[8�k���雦�c���&v�s�Ῥ[��[�f`��3#A�է,ҽ0��*�Z��7��6��;�r������zK���ʂP7��W��+i'�=ц1�7y�̩�ՑsZ'�N$("{�ؘ|�������S���b��~������;O^A#-�71��iϋ2.9C��c�ioJmsd�����} ����U�������|�Hf�^af^�(����E����"�&�_�2�W�5��ِ�*P���d�Z3|�O�����`R�%�D�z�}.ئ�ӈ�o�����U�"AbH��� �_,�9�^��=BB�;�^�@�en��x{�$Q�_k��`��IF28(�c�4tU)�ڄМ�L�2��x�po�O]�|�B|�:�k�O'�RU�v�Ƃ�Jqq���{\%�E��0�,���dc��ܒ��Nq�I�Z>��&���q!�B��u��4�S��bX���lK�B�����
���`�ܣ=GJ$K,O�Prh`�w`iTwlwai��lB�<��<��[���u�K�Nd,�kBdrHvN)��jh�j�aN��`Y�ы�f�g�Eݛ	|�ng�ߕ�n�i�6���`�_�q�;f�F���T�T��i�w8l�+�4.�:�w�8�v���Ƥ)�6�@����^�h���Cdw��9�T�_�>�븿v��t^���,A�a��m�0?�+���Ӭ"�����c�}҃{�A=r�LM`�&;O���qr���e�xPj{On���Ϗk���)�����i�9�U�_D���u7�kVҦC�:�����ޝ��Pq�;PEŀ��'��W�)��(�ҽ�`ѝ)S ҟ>�|*�
N�$�|�uݱ�M"��0Ӵ����t����٪�:����A���>av��&��v&`������� ���Ì����M��E+�9Y�Y��޼ϪnA�������}���|�w�B־�- cL�a�*4�\� v��L?�式�72Q�;)+}Hߔ�[C��YG�<���I�ZmN��EF$	Lv!}7vt�Ȳb���[�;�EE�����H����lp�1ʤ+֫7]�z[}�C��l�<�aW2]@[�o�Yu���H8U��Xb��h��(��U}��(��H�p�������doW��hvw��!ߝ�r�;)�7��n�B� ���71[{p��֭��i	M��(܏M�Q�@C��Z}�B͸���_ѹ7��#H�6B��H��I@[CPPV��c�\���#q���&�[A�'3�ʫ�nW�ӓ'7ƥF����"N
��Ҧ]c X�<u P2�Y�i�?�K\���ư�.�!���N�_iE0vV���]Ɣ�_�V�OcPK�O�s�a�~jE����Q�΋my\y:��k�`���:�[Ҹ��8��ǔο"�$�)�q�h��!,r�s��������m���,s�P�宜.�)D�Ӱ���$�yVT���T_"u_~�z����=�-'.�=��SUJ_	j����E�zj��7>��q�M>li��e�p��o�� a���R��C�||*��5�.��6~x|�k.��t-���$Pzc�Y�_��ŀI4pF�+,G)k<�v[� m6�Ηq�\ǣ���B2�ܩ+��O���l��(̅��0� T�&�Tݛ����]� �s�yG�K裠��a.ǘ���G���5dZ���=���?�#�MR�b�K@�*(N<�i�b��TmN�VK7,UߙK��ڤ��a�0r���|���5�<td۸�c���GU��5��������\\��Xi?��`
~��D��
xj@8�:+�ű>�W�v�>!�k��3�{Nz�i��͋�xV� �I^��P:�]C����@�*n�.���e[s]��#�7"�UK�9Q�͝c䂱��5잎h�|���:;���kT29D"�A���~�q t���$+ځBY��z҃'� �j���S��
�	 �1��BN���e=h0�!j�����TY[~���w+(�	��M9�P�|�1I�C�@x�3S��nv!���N�Q��~���W��E���P,F�`��wA�Tމ�0�+"t`��q]�DSî	X�M	�5�8�r�)&�})Ԅ9h�l�N���)*�p�Td�����`O���mdR� �M�c�NX�Rq.���[D\R�Ip�!;W�먜�(~;쎍�Y7���;��W-8� ��59�6����H@�	���W�`�Խ�S��Mk�6yo�'�^�:�����:˜ ��\Y���|��be�M����KT�^A�eB�!�DW��K�����e�ҀX�a\\y����N������|��낝f�Q�ۂ�!����Q�Ǭ��v�����]�E�cD��r����C)�����N/�`Sf�H���6��1*Y��유ǭ@����M�V%��{1�[�LF��k���ǖ?M/�ލ�E�ܸ�ߠ2�G�x��
GO޳޻v��0�Ѹ.z�@�/��q�1�
Y|F{TL�L9k@���n�j���ɐ��l�A-� �c| 3������`/U��N��1��p�)�|��i����!h���|�{�jcl�f���~�a
�F���%�]��-[8Ε�tn�ؿ���=#�Ю�	���k�?S9�����B"��� %�����QHC�|r�����sC������g��{��"��w���r�S�Q��6��9v���9��V���m�7Zt�̋�Zpr�^pN�:]�b�+Q���Hsd���P��-���/�R)�d"ʈj��UY�uq*�4G��'c]3z�J8�D�>����<��s���jX?����a�Oks�U��Ϭ�2��E����m�1�f���4�<��\:\�|\�K
F�!�����t<�N�K�L��-.��1�L��;�0lUF}r�c'����%C%�?���6O�;��0���{~�ڥ
^�ز`�;�����²6��17}�Ų�ײ7S�r��I��:��o	;v��2O,�"lO��8�*o	�LB�+c �du���r����M��nL���}�]J�t�.�
T[��D��[���2���Ժ)ٓ�\�/X��ǻ��+!1�Dl�/&b��s��7�=#���`߹Կ�9���ް�Z��,Y���D|��.�7��=�� �:a78ɪxW 2(�2�a}�甅a4���C�%�`��������e��c��$�C��2+!�ܑ��2(Ʒ�C��O�d���7И��Ca;0]��o��׸l�O(�O���g,���L-��%�vš�o;��woa��]�k�a�!�����M�{����-������Y�xK
��HM ��E���qD2:ؗpR�
/���_�p�`���J�P�.鳢�#"9 ��7Q_T�Ew��q� N
�Kt ���b�4�0R��ͤ�����į�
��qc�g��ɂg3?�����?�̛��t.�?��3㫝�3F@�]x"�t�Ć�d-��/�<���
��ש�+�<� �:���q�3�����D?��=K��4D�	��+{���ԗX���"Q(�/�=-�d@<�g������7��� �1m��8@��Tv�f-�t������[dm=�-��#��Į��ফ|��#�O�כ���+OM��w/�(�:$�1]�3�q� b=�Q�����
wCس����g�W^U��MK����J�4����2�v��6�8���qd�_�9,E��������I�	j�"gE�HA��A*��OQ��J�����*�(�w�;��%��Q9݂��[���1
��@
�8�,=�$(v����~�@Va�eS=E�o\c��ء��J����S�	H)K����>d� l�><���5��Ig_o�wR�	���� 1m!̭�$!�"�IS�����N��2��4��;��������P"������i�����|����c]�g��曺��p5��Gm�C����
��R��b7�l�e 5V�xLl��oc�sG7����כj�|F���WQ����1e�@~��4 ��S��Ak����Bb��}�@�z�7������d�N?��v���*_V�J��ژ���dk~��/6�e�s�}VdK ���C�p��Tg���9ė�́��;}E�daُ������b"�R�� ����S��`x��+��7;C��o�y���qSr�M�uƜE���4k]��5���f���?�gnG�\�B���f�Z��Ì��wFґ���T�Fק���I�$����r{<�d�g� ۢ��{���/ �����g?�碁�� r���+�	��A_��2�?8mY���UM��%�|���!�S� �c�������*`�f	��B8��P�_Ќ�R��	�~/��8������+���C��"\�����z�/�r�c�A��B���x���쀪�� ��m�yŦ��F�@x抒����x�J��Ȁ�Q*B'i�g����|�
T3TQ ɓ M�b2WEy�0˗�?����8�t5�F��[
��K��1H1'-u��	�}���hƛ[g�Uq/�y֑S�&��w�B9R��ҟ�,��`��Z�d�d�/�Ik�L-�'��-�mk���'jDl�?Yr�>^&N;�́��=���I�y�}0�ϒ��Zw��Q�N::����� Rkz4�k�eޘػ�f�5��EX#:z	�E���d�`����G�� lDc18�b�f���`�2�ѭ2���y��.�MNg����Yص���ˆ����\'z�qq���eh�m��w-�"��^v���_2]�������ͥN �(���bʋ�c��K����S��יу��j�����\��zd����>R���D��;N��	]�S��T��%��Ї��%
��r�����m�7V��G�GE��|
t4�ߒ՘��ap�Iy�d,ɦ�(Ih���S����E�D�7[l~� ���^����K������5[y��>́ �E�=���R��,�H�+k, 4��А���+�� �Q��u�o�^(��qn���wNF7��Sg�Y�Ok*�k仿�X�+(o��Y9��`��<~p?�Y�6���7�]��;�BA�1i�~�����1���U/q��K"LC(כF5�7&�7c6� h�.Ĕ��T�<�ۦ����������PP4�&Ȳ�����L8�#����B�༏�'է�A:H���]	�*�%��6*���t�������+J>~�}2X�ݨ�=-�T�Na�0�9x��� x� ����	�#���PaqM��Ͽ�6b�~r{.��'w�%�D��儧�Ɖ�� �S�\�l4��f}����k>�ǟ�W�������
��K��6�|���"z���"`}r�O��2&*D�b[ȈɑV�/�t���x`�r�� ��ը���St.ir�Ng�.��"?Uuz�R���!��H-�Ɔ8\��I�?�!�gYM<��6�vc�a`��������Jp��ܛ��4��a�!MT%�p�r@E~�|��h��s"�����<X��hz��u�R
qI�����D/��O7�zJI��g�9��;����i����R[�%ݲz�}�i�F�j5�.��n������pVYGavX_�����a�-Ȫ�yےsH���R���Y�=W!{�R���2��V�ʂ����?��ɶ!�T�|�v���Q�2��8�G~`�N�������c`τo �Y���D�찂��#�t��u�c�B��>$���5��pw�i.A8��B�{��3qF���E��$p|<P0�M�w��%j����H���s�mVd��s
�\��8��݋:6�����i*nE�����"+����$:���Vˆ�V8%QXO��|.A�a�z��^����w���u�%u�nr����EH�{,�`�k�b��tb� l�"�b���� ��w��3A<�J��M1{�8�v���X�Ps`ڝY��
.�N]*��\��7%�~*�Թ��V�p�����=2Y��_�g���C���F	B���LmM�'+�����>�;���`��o�V�4j����2l�*�U ��l)Q☸�p�|����X���e����̘���9�]���X��f���G�=��>ߞ�5�JgGA�w* ���ECy_/+�&�����S�wy�<���G޺���D���.b���,	��H��X;���;��%[E��޵7�h�M��0�w/.R�/R����M6��E3J]"�W�1�glj69k�g*���d��
I~���~c���L�^��GI�q*���'+���g���(���n.�8܀�xw1�1�x3E<��.����{�^����<�k��h�_ǆclv���Z8&��;=M��ij�Y��t$'���e��[�+y���*v�È��%{w��ͱ+�+��S<Cߢ�p*�y�	�,:�n|���b{)&HH�ˈ�K��:~�VYёR+�	=�>��m�VQFS��:� ���+EyGl���v$j�@�r���f����F6\���ԝ�/�ө�Qѝ�����[ۓW"K���&�%O�ԍ�b4���߿���H&W1���n��a5uى
���� ��A�Jh^�ߟ8�w�*�\\Xj�6}r��=1�x�6�wξn�S5۝��YA���`���u�VD��k��"2�GG%���}���3G�����<[��hQ_ �ރ$OTf"؄�4z>�v�do���%b(_&x���ː� �|�ݔ���cBvw�)rXV�H�9�S�_cs)�l�+�5�s/�7ņ;�e�����Za��F�h��b,AG�2\ؠ.�4N� +w�Y ��f-2u;�=�~u �kZۋ�P+V�	�0`����f���O �O�_��@�ߧ�~�<?���UvtƛS�//<Ge�~|J�k��E���N�=\�2V�T�'�FXv۶k���wSdԆ�ڃm�g��y����,���R�g���"J�R/�qi��w�<d��j1�ЫE��O���6m<�����0/50L�#����0��6�c,�z�1�gyDS4UE=���s�VM&�<O��v��*wlN7d�RNm��# ��K��= m(�T]b�I���9�X<�(ݾ��A6>HM��y����pB��q����Z�/i�0�=�i�k) m���A�5DW�{�ooFYw�PV�0M�N��� �u+'�otx�$�f���vq���<�C��@�Yln.�����]�'��|��_0B�JP��;�@�M�G�a�!{����)�~!����c%3�_s��4���3hr�����F
�f��%Ť4Qx�^��(Y�syrU�.&yF�-�o@�$��|����2Ö́$���s'F�UuR�1\�����v{��BV��T]h?�dG��h`���eU�oO��L�p�ޚȐ@K���X�z�2w������[k��8�ty�� ��<~�*�/�.0�n�>��B���]eQl�De�um6�R`*3]���:�6D�O�w�s7|dWZ�!�!�@�w9j*�'�.�zɳ��{ ZHZ���}⬂m^���5;�[��&v;oE%L]dj������v��Ş�U��W��G]��	�`��\����9�K�H��'P�Y��*���ݯ_!ϔ�ٯs�1~�&i��h �����Y�2�ɩ��;���@�pzm�i��f�>6L)����X��@�d	(Yn��0��H����B}�k����l���g��:���B�)Xd�GRI2�~2��	�C�����W�`A/G(���
3������M���z���;��EU�6P�Gԓpv��ٝ�P��Ǡ�����w��_"KrÂ.�@�A����UT(�!�&QN2y�d����qm~���8�wA�؅H�l��j�)5"����q�Jk�J"i�z+0,��;�ߍ[��7.�3�$;)�׬���>(�@�.�3_I��v�����^�/����y��|��9�t�
p7�1�$��p	j'3���X�-ku퐈�������z��s5�~�t���$H(P�ܦ��p���#���GXx%�\�#X��WXx��������B݊C�/W$��0�Rq�84�M5T"�����f��<x��~_Ǔ�x�*T�<�Uq�2�o4��~��x�E\|5t'1�6evFZt3�x�?�8��" ��EϮ��5< �+�A-
�OW�+����h*.����o:���ׅ�K�}���
9�A�����ʪjONϹJR��ڍ/��=�_�+|.������p!?v��v�T��sO}�_��ʵ\�JKAHɺF-�?É�V�؛���7�-~��D}��ݵȆdc	%Hf���x=���M;<�_i
������el�ׄ�/!^oe�����܃����_;����8����ޓaTIB�Æu���:E��ψ�ᅺچ�������|�AA 4Uz�/�%����Oh��XF�<������E��/dl2*�M$�(
K�G������!n^��"|ŹV�.v�&��7�&t�qp����i�`�n����q���|]��8�hբ
��C4���9��O�F�ġ'-�f�� o.�G���{�r��Չt̔�Y�XqJӨ1ϫb�s�;U�,��U>U�4��5�]uq�wyS������P��V𓜎�������O=Hc�!P��,'��Q+��B._��u\�{����741��o���k{H��v�J��wҺ�a�F�Ѭں�DĲ�̨S1�=uːҊT�FP=ɜ�/�[\�x����b�xRƼ1�kМ�I�Y%�U��I��G��� ��M󢽍�Kg�Uw���0i�	����-����ėf�73\�A���ӓ~3�ܫ�?Ge��z�3?��V||CW|�o��9R�~辽�_�'��yYb���ꍪ9���S=.��6�@5�R���*6J�ہzN��1�7i�m�I�b��,�߫N7�����	���ǏniarR�\
�vƘ���]��d ��]���R�
vD�m~<WE9K��|aqz��4} ���h᤻�@��&�1�$g��|�-��.���e�	
r����6=m�aE�2�+E���AΟR���Qc6���yIf�2�I�J/m	<#a�b׶:;����8>h�3��SL�HU}��>��q$�N���� \���}���X$�o�w����`����dr�e�\�)��=U��'2���^�2����L�$�?F~��c����+@(�� � ��Ҫ
��;0�dG��0�
4�+G�*X_�	
Yڎ�	���/x=��]R��h�n���R=�tf�h>���� �)��k:�����8��|Ɨ�ֻpW��[���6�#��+-�[�w�g�>��/&w�ipP �i�6�@��Ma�X��x���x7o� v�n�l��<��Ls=.?�j���ޘ�!5k��Ϯc5�xz!n*���)�޵��Y��Xh���a~��z%���Y��L��;�ц
X�K9��>�[Zz�n��F�do�B�,T��]�V3`�h8�z_)2ǚ���"�2��0�fW���Y��(�Q(�b�7Y.˳��"�}�Y;1$'�X��Ҕ�`�0/��2z�+��yY����"���y��F*�9����2����;�����88��8�+���)M�=r�_T�������/5e�OFo(.Զ���
���|�m<�8x��<�!S�J;� 3��:���OJgSg�7ۿ�A[��'�^��/Nso������р�"�`	��&�Ы�vkw�I1	8��7@M抶X�ƫAz�j7����˿\�6�9�8��p����w���ɒ2�a�F�B��O2Qpi|��b_��kˢ�v��n����9���R�z��	���0��^�p���X/[����ξ��:QT��] t�5��Ӳ����!薵sMi��wt�
DAݑJ&��SҠ��5ZC QU��m2��rM�MMNW�Ȟ{ƥe,h�9�9����(�m��I?�m�g<8����Ix���4@ܩU�G4�N� �{C[���c���x
4����2���S
$̙��}���р�����Hރ�gh[c��lg���) �H�'<���$����3�c��P��1QrUݨ/(�R<�1��<��pj�7��,��ԛx'&�X8� ������X���)Z��g�#���v�(�jiu�n�>�)l�|�S\���,{�I�0d�K�;ֹ����D����{7��R�pg�]��3�2v2����
:&����hC]r�s�f�Óh� ���E!���v�ލC�.`A�o�<��>�
�j�"��^�d#�;&d�����'Hg[�x��մ�G� �6�Ed0���KUպ�iQ���Bg�|'��K�\ʞo0-a�C������<ǭ��,8��T8~��Z�����)��oK� )�b6W�U"]��xlF�D��`��W1����`�#;\��V��g��y�?yP�K�բ���js�LO7�\w��O���P�T3�y&vΐ"���;�Psi֛�w�Y�e/��_�Ѐô�!ěedA�?3*R�����il�aIR-�N��p$��XW���CA����_N��Գ��r��]������n\��0~m�#�P>�Y�<3��}n hLU������h�M;�����o�W\(~#*�7cdp'��L�����yN���g=l#�����s��*M�?���f�$��Yr�#Y��D����
��pSoE͆�C�y{Y��_���	}P3�O3E��ڟL�Z@6�^��ƨ��ϟ�Mc��z�em	�@ȥ�4�19yv� �'���Py{�t�6�����{�i�Ů������-�;q08�ʖ6�beL��wjDֆ��Z��FM���+Ob.Zr6�/�&շA��<w�v�ah�����`.��IK�Ʉ���e2�&�z�u�N�߆/D �g�v�w�h�띜ęE�J��i�{Q�R&^{��]�L�����m��cV��l�&�V��
M[�;V��m��>�Z�	�]0f)���=>>�|��JyV8�IF��H6P���h���_d7������\��F���v�c����{��j���AmV�x��`W��as0hs߼dzʄ'W�����h�0"��P("ؒ����B��~����:���QI�v-߼l&�x��`r�-�^(�!ں�L(�dj"������r����i��P�g��91������(�_à'o�vQ��"��p� y(��Uӝi��j��sd�N�`��(>�/}GG��ާ��5+�-_�9�=[�<[Ea΃�Џ���a<�s��*^�SY�Ĳ�#6�P̽�;� ��nϼ�m7<қ	*l]n�^H�>/���=��V��>�8�"�-j�Wm��|�W�EJ'Lđ�H�r����'%2�O�3�s_�v�IS?�)Q4��4�������n����zC��n�"\N�]���U�Ĳ�w�>К5�N�C��~D�cZF!��W	0r�G��m9D��<��$����%`�C��j�8i.�֭�i�F���=V�i��3G�8��ئuG�������;!q����S�V�\}�o���`��*i�w@������@��_�1b�I��^i�@l�	�	�@�!"�������r�vH4ٿ.�G�2��[Y�O�r8Ώ�g�8r���M�1FN��:Ǭ�n������&�HS�FNB�����߭@���.| ��b�H�~zf6� u1�Y>;Dz&�hs�DB-</WSw��e��)
�Ҵ^Q����d�%�c�f'6er~�G��]����
6uҥ��t6!�h��$dW�.!���YYK0E����HBu5?()o����|�A�!�J��Ή.��0ǟT�bR [�PoRD.r�Fʶȸ�b'�2T D���B@����+ޱ��ِ'�2���{��"����9���x���X;%ί{ �I�_�;�9Lt� D��o�9�8}�9���<BM��>/��e�>ʣ�RZ���Vq�2Sy�!�"
#ȸA�o�
�?ltX�;b�Gvh&3VФĠ���������jx�����e�s)^'�k~��ХЈ� ���h�E��@e7Z3j��3X�A�D/��i{쑎5��>p���i(��q�N�9*�O��<M��5H�hy������:<C��3>I��7l{�Up@����T1���"�.��}���
wlePJU�|�L_�r����uq��H@�>�#��	��4����`ȆE�6��\���F(���n��X�hӫ��E���CCIo)� ��	�j2���Y:�
H�G� ���J�9SC*�ި�cw���q�I����-�Xד�5Σ�H�r�K(����tv�I�y��Cz�����v��.m��\./=�'��������3\�դ_����Z��G���`�~�/p>`~���p1
F>��f��~ÄDff���f
n+�>��ʓ�Ɔ�U��X��am��9�� XXw����R�K:\!S�B����U<�H�a�� ����i�F��Z�/�I[��r#Y��|/z��Zc�Qq�HW���騶b�k
<�{��/�J?��b���f���B{����|F6���D&�M�߽RD���?'�ٮh�4V[��9
�ߞ(	��v��{V�+l]��Qjs��0�f�m��N�kؐ����51P���1�9�q��3��ġ�f@d�!���������SBY�����k��6��|�ΩJ[P���]1�$e&��pk4D;~�?g*Ϋ�I�Pى�����_�S��/�!b��[�F_y�9,��W����G��$fD���.ʚg�y��=���=�M�f�q���+�Byvĩ�
�šC�����'5�ڦs]聫1�]�r����h�� 
��0
$˳��)[v��9������%��/�J� ^�z������w�j����t~�ᵁK�0ZZ����V� 8K���\�1�^T?������]�r��r̈́@<�!�Q$Q�~��� ��P4�����է��8U�x%/H�Ҕn�:e~t*_�;~�G���b�������M[.G��D�\�}�c�������8��Xw��1˒`ƽ�jYa60�͗�:�A=�Fh��;�5� r'���*��x����?���U-�{]"�#����������!�+3P8DΆK%�h���	S?����E^u䯝�9�j  �sK�3�>�{lSN��<OFQ�9~��'<1�*�	�Z�%�,R�����1����b�W�]�y�cHy�C��(1/r�#psY~��";�H�sʏm��1�A��L��?�E蓯�D�����r+X�M�/�h��	�h��4�M�Gv=�I�#D2��k�!�O��ұ�N9��;OT#<��ĩp!ɉ�lj��3��6�3-H;�95R�3�I���r��|㐴�ޘ�kxėL�=����k�r�����?�=;<��9����l�&Օ�����B|����;E � ��Y��S�;H)�;�f��Y#���!,ʧ��'=26�v�4�eЏ����ݍ�S~O��!�l������T�����Z�'w).>0���3�$��H-g�%D���6��góS�z�Z���}��$�*�ڭ�p��N���I��6��K�E��@%t|@���^BEU�mڜ�^���i�p/�K���u���s>�pFz�Jy�UO�+�VK����:�A#g#�w*amؽ���md�Sa��Eu����]�Ŷ)�� �}�$U����%F&�eV�h�"�	�R�*��_D�+H��.x�Z�۞,�2��P�c��8ĕ;]�2h}ti�a����N2��
�����ꊘt�e�R��;�+�O�T\�s�z2R$],cj!��������Nܠ 8��|#YxUy�u�><�e#�b/ �K�d0vʂ�!k����m�Z&��'r�\�� c��9�����Y�E�F�O�C�z ��o� H��~!Q�)�t�[��s	A0j'��ޟnpF�ӓ3#����D���6j�b�2k�'sn&t�pp��\,s�aU�Z�W�B8�`�n�4�ߠ6����R7<����X:Bn�ԡ\��!��Y�$�ݰr���x���Jw�y�M|?�~�IlZ#�@��iq��|`�J��6�>M��xU{T3��3�쐣��?��L8~���4@��%;���.eE��]� Ƽ͢&P6�U{z�e��Z�7�n���}��U�
H:�&��70��ۨ��?<�`|vg���>��c���Q�w\c�G�Ѱ��}�uy������S���zĲt�r0��q�� 1���v�Y\M�á"����r�z����Xv�i�[�E��������=N������a1ׄϳ��\�1x�-�H�T`�q��i���qpf��[�J���0V{}�ۆHN�Ȋ�  �jj?N��|� m9h\:J�L��7T���O�~mU>�m�����N<�w�#:�&� 2���P.^R>��H�SV~�F��nBh�'?�+2�@' -x��X�o%����^I�4�~�Q)�QV�f��(l(K�݉aQz�j����p�*5U's�X��[�>$?��K��K���m���`�%M]���VWBy�W9�]�Uq��[G����y:?}n�;Z��7}YrXƐb�=�'F�e>1����E:�.�8=��>K���v�>�W�pI�T��(��*��$��B�跔��.hx#�d���x�����~��W�}�&��r�|	n��B��Y��{M���j���]%L�*oĭ��F�fCK�����T7��"ݸ����p�|k�� ��s ƫ��-�0)߫x]e����MC}Q��.�0<9-���y�k���W8�=�A.N�6�����gm?�h�>�4�F�bT�K��Hؕ���M�k�M����/BS��+}���ɻy�%mT>��{����5��)[����F�;CKo��//�w��%i���{Dg�#�������t��U�9aC��!B\��r�P�����)�U&4vx�k�D���:7�:b���0��9	��i����b����ۺnU�8�*���]����u��N9k�"�k�՞�v��8*��k�L:)o\�(�a#9�I��BR-��rpuL�V�T�"�����[�Y�G6Zւ�:(Ӄ�3Y�2T��v/�`� 3���	��a^����J�L#�i!��*� �oF�V�-�9��\y���E,>,F�-�RrbO�#���~���3N����͏��I�P�ԥ���?=H�hy*s%��wJ�x�_&yj��"*s����l�hL '*���gZ�mP�Ma�ۖ?�&���.��/�]`�j�gt��=�'`�ճ�������?T��&�ǳ-���g���%���2��>W-D-w������g]��L��*�6�wE��C����`G��E�\Ja�V'���邡2�i�@�%�%æ�� ?IG��S� �������6����	���"RB���j����Źl��ؙϧ�SS�O:��}��r���7��S��c63NM/���2�n�Hu�k����G0��o�h\��V�V�Q�-jơ��\��
Y�z0j�t�~Ro� �~�����> ��6��Ҍ�$i��Y(m#�w^9˟1α�A�~qD=�/�7 k-�_�h�}��ҳ�*�\c6E�N���i7�9:��d�.	���NiT��Z�	�X*a_:м{>SV}�:<9�Z[^_�����琮�SZ�xH�\���Z ��,����玒!���eZ,����Î4�&m9e�����"F�}�E�.�ͼ���%E�#� 
]��ѩºř�Z�kMC���!�DE�r����K1G��R��JPJ���c����$�<����
�A��S�#�Wk1m��x�Dy��@�#H������q�y6m2�C6��fVL׏�I^��ݳ�N/��)�pG��A����'l�ϟ��0��X����>8�3�
�b�'�����Մ�g&����#x*�Z��!Lί�=Wd���\eਘ�.C��{��w�JԒ@\h	a��su�$@�u�0��m|+�"��	T)S��\�����9�A�F�P��҆:.����GZu}�g�ɏ"zNF�^�+ �"L�%P�G�rî��hAN��dM�bǱ�W$k��Co�"���[B-��v�Dzi?���V٪�.��BDQ~�*]�Fk���s7%�mN}b\2CzsH�q����'����h�䂿=���`�������:�ʋ�pH܂E���mo�F��4��3ІCEףwy���2焓��/G:[/\��'���z��:���x���B���w��-N�v^��6��A5�豷��6���<��6ܐ�9y.$2��w(�M�u�vM76�����w㐍x��������T����"��2�V�.���8'Ҷ6��y6B6ą+�Ń������)�w�#�US��5��G�j^��I�9�?BD�ryhv�/s���43��bɫ�}�mW<)_Q�9�\9���5��q��آV"��G�5�_hOor+��e@�h-��Tg�ɋ4	�kX�!�]��'X!ݳ~��+��3B�hr����J�mj�9CVrѻЌpDo��*l{h1�x��N^�D$�a-�&v��@�ԉ*��e�<T��ٹ�qp���f1������p[��Qh4�J��t%����0�7i>r,��'�Sd�O��HX͖��S�&�7im�%	� Jy0�[�
�^А�C��h,c�`E��G���ŭ��*�?}O{ꊾ���\7k��d]�jr9�����Z��}_�O�*`��a	��H3�Ό��h�R�~����;o8k�_}��כ+6���|�L*�����q��/�}�'����`�=��q�f���ñ��ɰBU`�#���K-3eY����F�;���l^L�Y�0�>�M�/��ImO������\�:=�U��Ҍ�!J�_��7{�+]�g7G౪+\.�_��kTac�aL������� :}H	8�V����dS֡V����/��&��$��b�-�9Ru�bcE-��cUm,�<��zA���P�H_�7���n�8b�� �}���X>Ѹ�p���,��bp������z.���[;���%4,�>�Y؎
2V�� �������-V@��sQo�h��
\�v�������ˆ�\���#uץ�T(n�/0$�W�M��_�����r-��-M��EC���CX�hT��jף�W�ք��p�.�������Fl�G-��t��r��y;���s�#�I|��v�D�Mmh`y�H�$>�م�'�>��@��~�.��R>�Hu�a��RZn��C��#�
B�]�����:yHD��߹�w�I��Q��@rk������Br�� ��|���3l�NY�@/�N�n�GzE��mB��@%5���m]�8+2��@T�j�q�F}�b��p���1+�BU��)���K��,�-�T��t���:����s�{!"�.D�>��Y���gE�Xv4�M�h��j���;�D~�M��Z_>���}��4���"��1�b��պߚ
�����40W�]}w9�u�O����P�oӪ �a�Z�4Be�h���s
�}�(�c�E�w}k��h�pD�oy�"�0u�T;��ȃb��[��*�U������nS��'�|&��R�i�A�1�
-�#&�9�CE�Z6Y����[�*W��`ⰤY���X������}�������D��K�����0S�(�tc�)����y2R$���h����5��0�ǥ�_��bV�r_o6���<F(�����R~�:ڿG�?�ݦKѾ��/e[����e3�loS���[�L������Ė$&�@:����e|� �}' ˴�p�֎O2C�$�s����z[Kh��K�p���"��:�J�lW�TT�TӚ�f������ůg�o��AN �-t�lO>q�WYI���hX��p<�g��0m�pC怒�PBV�v�����D�2�n�y3��Y�ގ{$Cb��<�O9����*u��c�x3̰�'0W0Mg&F��p���^��3
Y �<�l����wb
�Y���bN�f��qߟ:��+>�?�t_��r��^?LV}����0�q����(أ���ҋa?�y�b��k���F���BQO�y$LW.a�O`��q�>�C�i{L����g�-95�H�c�W�d��Oi���͋���Yw�
�m!ݾ['���U��Щf7I�:�j��L��A
���JcJ����T�Wz[ ��N�,N��WF����HX)V�]!� 5/���I`�{}H4��w�.���/�d�>��c_i����ZLБ�������YU�*� AW���v	����0 oS@��α��Y�׽�u4ܖ`�a�
���KF�f�Y+��lF�L�󍖗T���7�a�1�lh?����"�(� Ha�SVk���}w�P��������q3�<��,(3���N�ݶ+=TSG��{��q��Qg��67�J�Y=��O_�#�غ�J��T�R��M��� �vhP̜�:�p}u��^��>�嘅��-�#8:�x��"5��u	��d�,%�q�{Rxj��o�G���B��Yi)���zҹ&��:r����r֣�_R�$B��?A�{bm�j��]�f���'��W#Z��ܟ"z���c־IBm�4���K4�| �6�G[��w��^hܗ�P���I��\�@�Af�pC�Ri�:{9�\,���nsj�I%��|(�Q�I�ϣ�%fi�(�>�f��Jx�Z\cX!�	���x�j����w��(��J���=��e}��~����$gp���>7�k"|���a�U�)?Q�1��(e9������z�ԩX/ূ�L-B��p���<�Rv �V��D��ז�����~���v�������t"�T��Z���o��ְ���cef�K�n�mҳ�P�v�����U�?a��~��U���?-�+:�"j�mI�  6n�"��=�` ���%��@m9�e��̌�ۤ�g;1(�`�z��1f�0U.脈��;�c���X�����5#�� pN_�����G�k��1�@n�_�1:�e�D��:�7��.�A�V�^��>Ȅ�k�c���h�9�>F�>�S]��Ȫ�����>R�"&�]J��@�X�#1QO�jU��F�{�t8T��-���P0�f������B��9Q�C)ּF�d�+�.�# <�K��YDˣ�!!�A��?�����P<�;|p�
#4eP���l0��e��$��
��F����wR;6y��\S�T7ls��l��=83��v�Jj��s��t���eZ����H�(�T��!�-W���53=��m@`X��C�i�>~���_���[���e�#�E,ŭ��.r�1[{�ɣ��TBAt�@�����A�<蘪���ʏ�
���	6h"0����g~��-T/N�<�/z���k�AZ�FjH,	y�Y,A@����������C�=x�1����d�X!�ZЍ���{��#\�l��6��ں���#X�!8	|�?s�tg�ҎYs�y��4M���=�)����c�4��x��LJي�f�T�>��oM �zY��.�na`_��+;�}0�r�/�(X-.R�Hҝ�W�C���U�;Cn�8yɇ;H��
4荣y���?U�'\�)�������ɭ�~r��`�#��e3��/7=�I��TsдK^7�Q5#\��}񓼳�^ʤ�s���ª�$+��,P�T֦���r!� 1)&0�\�~�E�~/;n\چ*� d-r�g�U�=%�%����+a� AČ��'��5:��.��3��Y*�[�C�-y|���$�[9S�/�����u�|`�Cq�$�R��=�Gr�P��,j���d��\��tlW�zV��|�qt0�~;7��uV0+��)˶�������[�ۧ���B�M�]�U�5X��A�K4M�%���^\�y�~�~}����^���Eϩ~<�7.I��&�~L��@����dc@f��x�������|BrL�) �a����Ci��8O��n�����n��@�7��-:�1����( {��~O2����P^�t_�In^�#)D��kӉ�2��t|�/��QKsm �=;�^,TBI�A���f;��<�ڪ{��t�!rV��`�8+Е����Ն�es�*)��$VB�)a鲤���T���.���U� ��:G2���3.^F�>л���h����!/���OGY�&���q�^̎x+�)�_3�?7���Rr0����W_M�;�v�B��{��)Wt"�JY;��3-�����J/�V��Џ�{�Z�ީ̴1�+5j��� ��\�?����J\�r.%:�W��_�@�Y!ٖ�P����,д<���q=�_FHgP0ۗ9�׻J)�טW�<6!�+^
msO�c�!兑��U�<J����<��$��m��+nL�h"�F���� }��l@�%Gni�]�e�s��5 ��Y3��.��1�Z�e=:k���M��Z5j5�p��НI(LQ�>�'ю4�wp�j�Y�NAP��$3���jA���oƈ"�_�V���1�E���M� �M1G�q��c�<�$���R"[������+K(U�	dĞ:*��q|Y$�;�7��<�2dD�|H�7��#w�L&�]YbW�h?�H�m��K��$�%a/ĝa9f�?�m�u	�J��9�u/�������X�)�숥\�wgg���1yԆ=Z�C�tQ��\V��_E�g�?�1���q�R��������]�K��6�Kib�����:���a�U���Ѩ�tq~#x��0Q����xmr��)dǄ������>q)���%K*:k�+N��e��=�V����e�0�����Rq�6�0��._�j����	�XA,.��H���Ċ"�fIst��%��x}�B�6�8:k���u��=��P�
�zUth�
�]Y��6���F°���%�Q}� ��7�^��7:[Z.zz��ߒ|�r�jc"�X!��U�Q�m��9F�v���/ݨ�%����&ho��.���G;{�58i�\��?����!8U ��en�%� mI&i�������e����c��'5+G'\("*,��zI��Ԩ����z�kT\�4���_o9+áB/ *�(sK��ၡ�ظ�X��X)1녾�7��>�A�F��n��+�w�xN;�DF�����oo����/eا�T��Oh���$c�����{C�x�H�9����bf��!��5���n������}��	�}δlE6��#��w�`j�9�2�M[սS�&8s���W}�K�K;о�0�&�l0��O���[��폖lR��Aٮ��aW%��HN�� ,�+�P��2W��{}"2#u�4 �{�r��9�Eɩ�fը��qE�9��!7�!V�է�V�<����9��aՂP�9�Z��O!�^.��=���T�/��	J��k㡒G���O��=����B��û�V$��2��AGs1�%���[ɪ0�xk]���?m.�*� 2����+��&MPת`��	F-��mq�e���~��yri"��ˆXT�N!��E��-����O~[����}c'ܦ�������z�#A��V�-�n&!����fu�z�+�	+���x]ŇD��/!.�Z〙����P��J31��3 _Ŷ�oV�>��]�����B]ݸ��b�{a�o�}
hd9��j�,��ڭk?��/T{`�p\͒�$��CΘNePhͥq��e�ˍ����ul��`n�X�һ�Qd>�Z@3=+6˚�<�f��,A}\�{*&�c'�bf���с������T9u��Bˏ�󏯆)	S�OţE����We�%��|��O*Pd� �Xt���s�gfw�r��3�$���3�׸�o�Ԙ!�,��5�S�穗��������ౕ'c'�k��.�K��l�J�;���ǃQgz�:$��C9}����_�ʱd
́q�ߣ��dh��d8�@�����	rpϲ,����b'���	/��
�))1D!]
���ح+[:V�������B������A���"����9f1j{Wt�W g���n�n_7�2�vtVH�q��U� ����j�XǾL�V]���ԖoG�;�g��R5'\xe���W��gn��ח9as	���!D�=�4��%&d�z;dB�La���;�I����1+�F'�~a�ob�(���N�x���6@�k�S(;�w	�j5�@"��Z�x�a�&RGy���/�Ҷ�
�rN��*���%�4,���SV��Y�H<Ec,��f��m\?:��ÄT;@z�Yw�Y���@�'�X]��RZ�%jRˋm&}]�:�y���5���j�m�"����<zÂ&�+�p��Kc�8c����u���0�ցfw��Ϝyg�	ӝ7D
��1x�^:�r�+j8���<^9w�U��u���yB��gӋD�������S���mq6�U�_s�����BHG��e�����	�J�J"�5�Qa=zEŚ��)HƐ�eb�p�jN�4r��s3ke�8�V ���P::��
�L*�h�X}<-����B��u=��`G`\��}�Py�y�d`r6[�BσB��;R��ף��b��\RfFY�6�$KZ�Jur=�,�����U��K��j��1�}�a�N�/���˻��rI�r�1��Oj�=���,�;Qr�c��H_����P]�Ck�]9|�!���8L�ȑQ%zT1��*�����'�C�缲�12�!�0vV�P&D��_���J�J�a�9�)��Es�w�4�@u�P���oHfs�����9�y��j�ޛ��ys)q^c+ٯǐOe xDgq�ho�	�^�Ma�3��2�)<��;*$������فMf1�3a/���$�ބ�s�nP�Y�?z�[�]4�Y� ��}���Ê4!�&SY��#��pp�l���l{r�/@Q�������p0��k�%j�����XZ=�������2��h� 5�s��#�(��Iֵ�!���p��(�w����=�PCչb���;�x�1��hm�YD�ý�� ��7�Vj�!a6��wb��s���'�1���u����-�D7�P(��.�cZ��S��B��������C���:�d��7��-2��s��R���aj�
%y>&7*��␮�#6�2�B��U-ާ��BVH�5d�ؚ�]�X��[���I�ڐR������3^Ҍ�j��F��D��:�G*]'U�ԟo>�����K@�
��ڔ��ܢ��RfW�#�k��*3�T�vA�W�26�}ʃ���b��4.�,׾̃\k��뚧�M:�`F�<�-zg�;4g6�"Ui�P��x׾�^2���^���Z=s.7�R/{Gˢ*��2���^z�1Z��H����/��rM�͢�b���o\q>i�e���1�X�����f�P�{Mj��� h���=��2_�p�dz\qj\'(g������4x� wB\��_@���+F�żWpA���Fu���j���$�}���}��¿�5�b��=�S��X�/A�ys�T[�t$��%�\%Σ<�X`�=�k2�������m��S���P+��R�l�AP�ǌ�1�:Ȉ���K=�9�mGV_��`y����2y�ym����O�U���k[�feC
�0O�O �j�Q�i�?u�䎖6�����L\���  =�©g��)�{۶�@,�ԦRa��B$|���J��%��s�@��o��^pP[��v�-��
=kh���I�w�nj8+(�3%�}�]� �ӌ�U����F��|�=�[3y��w6��m
�J�Wo���ڻd�:�� �޳�ܮ|��{9�|���ä�&) �3������؄�R�vo�����x�����(��9q՛$,��&��>���S#@,)_,]Z����z��w���J�P�6���~�7���}�6�w���i�L��q�c��;�S��/^�cL�hdx�βQ�"F��QU~t�M�Ӗ��,�+F�YS�kb#�v�9Tm���W�% �+���C�Xl�����N^sP��!��<��[]�'�靮�����L�夝��%�:�E�i8�O��6lX;�c(`�:O������3O{%8G$�v�:ꄰ�\��;i(w}2ţ�
PC܅�_����^]G�۾]�sOJ@��ԍ~���٬��ȕ�>N@��۵U�>�����w\`���a����)K�d/4M����/��l�D���P�����k��:����7Y`G'��.�o��4`3h-��*�6��]g�C�hg��\�`M�x�(-!J!�ET�L���I+[D]P�	TQ��@%�9V���j�秊wv�AL�
��[ehx�/�o��@��&����kU'Wi�G��4.��I����T 6�V��^}�N�2f�\Bd/���[�;��CG������_��-�p��Jg�P��t0� �\
ah��! l�`q��z��8a1�8!l���{�\�o���)�x}�=���Ǉ�0|�����0'��p"/�k�|��^״]|�v��_�����@�A%��R�s���0.x�pB6+MPɛ|D�P�-���L���2u����yrU��ʶ�R,���^�=��cxO�]�T������!�aҷЦ�jc�xC�'��o�����v��-	����qV�O��:��)��t-5�DI ��&/�̊vH��4���$���`�*p��p� 74e�Ri��^�[��A�+�Q�9��ԧ.���K_�V��ڙ��o��&n=MWåwK�:6�r�lr�zȤE���(����oK�;xA'��r�� Z���-O��j�q��6y�{D�2���;�O��MfZ�%�zr8qY��B�Fo#���L8���W=C�����p�AL:W֮��O1�P5]4������o���SJ����� ad_����;��u�VoO��_��T���#�2��4:��/r�=ה[��[5Tb+�<�K!y�ix>t�, >�Dɻ�,���a�-��bR�z���*V�5|�����݇c+��g.�ð�BQ�(�����Z�Չ:�Pq.�1��yr�m�ia�