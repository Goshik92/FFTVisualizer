��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����T9 �0��\�0C���Ϥ���'ZYv�ґ��V<z?�xK���W�U����w��R�t�2���3|�1�ǆ��d�Ms/����g"��X��wT��G����d	v��d�g�B�Y0��g.����pP*7g���A��V�!�6��i68X��0-�^!�����{|�z!�S�w_�O��Q攘`��=���]x�j	�6�~���u^��J�7�;!m�<J���@	b������`�m&W�jNW!��p�\�.|uw
���%BP�H�5)�1#��QG��W�N4���r��M;�&�ʅp��"Sm5�]d�=���^�1.��-(�9�Jk�s�+gA���lwfH�ϸ'v!��*�& �ة�97��O÷*�"��u:�xU�) ��J)�����aPf�Ɇ$�zV軬X1����ƨ��
K -�i�?r'k��t����&���D�鬅_"�fV�5�}�M��ῤU��[�n[>��~��&��O>EL������I'B�B�fy@�bD��4������5%r^��Ur���|�:�)�����u'�$�80ZG��w�t�-o!��}��%�P�/���nG���9��:���6P�	 �䤫Hk�}}5�+��r)d�r�����z�mOs����W�C��&�^l�`���� s�3Ķ%zF�D�:02�׾�Z\�C����У��3��-{���Q�#DW=8R�Ѻ��M �{Jm�+-WՖ�A���B�E{�m§}P�m(�$����>�b�)!-�[TS���."��c,2[<�����bI?HC������[5bW����F����1$�+D�o�Y{�o�yrU�ɠPN0���\9ӹ�W�Y}��X;bv�b��чU����l�����+�!�H4v��祥X�S���Ѕ��y�~����=X�"�y�I�3���L�� ׊�D�h�0h��g��'Τ	!br�;���dM}���B`��7J��|T�m�5VY0C�P_�d�`Y�G�Vvs?���~ &� ��G�j��}M7��Q}�ɠ:�sA'��ww�p�&h$,����)����"�b{֕�h�)����"@FO���
ƃt��*���]���5"�%��v�#B gXei���+n?�w���T�6� �1�v�qHv4.�����d�f�H���~e�?c��
� �i��T!������7��І(��R�sA��׼�O�	�{hА�7TB�r�i�{�-I��|3��r�{���h����~Bڜ[<��=�+�;jym$l/$�REkR�,�Im��@�c��T&i]����2?�IQ�[��7C���#�KX���%�sv_��4�����{`�=�~��b�LK#z�^ߨo�
��&˵�}�a�2�:�c@i��%݇�%-�$�ߨ#}G��+�%�
�,�z% 5�����'�S�R��(�/ �Z���р0�"a��(�����~�nQ��8P�d��9�ߐ̢	���?�@Ph�q�dt��*�M*�d�rjŔ!�U"����eD'[{Q&	I�e��1ۓ1�T��� ��
+��s�Wq�F� x��HK���]�p��#�%	� �B?-KA��KU�׏)>��H�٢����%�=$�-.1�%�����2����^����0����Fܵ�?�B�eIq:��H��{N*�fc);�2�M,Ce̋�ώ�ۧ��V8)�mUm�~!8N�5��l_���V��4�6�ڵ�꺛��J�x��x���8_�ď�1w�4|a?��@�BQ�@&������4WE��G�t��5��xB!�j2�;]�m�x_���Ƶ��}i��|o�n��j�̃,���ϛ�ɏ����y�"�!� ���(���q`ʺ�n9�@V$��e�|o����|+5���bO0E*�W�Z�I1�z�f�)ÉL���λ;�
홫b��O�����j��-��Aze\�jp���Sς�R'NxUUS�ց ��HJ��6}�`S�۽nېy�g���s��jI]@��JF�v�I�r4��$>Ϩ���s��[*nP�紫�N�1�<�K�6	��F�A�^؊)P�^�[�&������[��jm��w���5A^��7;rU����U=�|E��+TX�m�{αi��X�@ �s�j�B�:,�կMn�����Ӄ�0E�F��?�{YY)�>b�?��j��"Y��ԟ�=E�jn�� �Оq0E�&Jl���oLd[��s�K��X�	b �7J[@��9��2�U���\1����i�����
�I#�aQIfW�S3hSh,�I��#'�V3�& m1E0`�Kq�J�ƺh��H%z�&��^���/Q�?5�	�/��[ ���6��4��P��s�l��{�e'79�V�d����g��T����!�^�!hܥ��*���PL_�������\`c�F\�i�� ���-޵�M��F��C܅���Ш����{*w�M}g}g�:�f�BJs*�����"�k��}��׿�nd�%w�{���3S��Rti�Jz[��w2n3Wԍ�𔃕��l͑��`����q�5*�����c������D��k��� �Y[�z[q�qBu�
?�� ���2��l[l��^�Mthsy� �?<j����L�VE�yɍ�c�;ʙh��L�+S���<;�8Ea9J��Yǩ��f���a�5���NX�=&�3���R�u����E��h�%=m�c�-�q���*��/��&F[���v�F�� �!"Za��L��>>xw��������L_,|�f�0/7��ŏ�n�PI۫�!�ۨNA?O��Bik��\{��W��GH؁�VE���d,���W'P0���7�Dg���D�0$h%4�"=|��|����Ay�G|g�s/��!=ח��|�J�O��E��kU����ة`b��)LA��NP�`M�A!����kw7ѼQ��Ɍ���M���G//���ڸ�d^��ch2:Ћb�����k��1�7B�?�yzW�#��VI;�-J�>�!����8���6Ԗ�\,v��K#�﹫�˩9UA�^�.��pa�B�娬��+�BP%�pI��_`$����!��s��p����$VIZy�]��@�f�eQ�X,��AO1.�ŭ�c8�"iq��j��͝��زQ7NB�(�
��uv�V,b��ذ��0�l�_����&�D	X�`0DY�(�43	�ׅ����m����Tm��8r��I�b���
��7����ǘ���߮���ů4_�`��A��\4(���w��i-ŉ���1����:3^��������2�7)8(�a����ע+���7��O��ƗM�?��0��W�u�p�^5;y?�B{`DF�!����Z�y"��|�Zd��\l�a�Q���aw�ȪK����]��]����)�E�p�����$����;�Q��B�>&v��5�>���V���5�Sܤ�����f�io�p����=71�(�ɾ�nU^�(O��3�|R�@]n�;���T�h~�ω���)�7�\���'ݣlù(6ް����a��w�ZK(��IZ0��*`\>�4o�@�z�d�^N��h"��$�,��M�]�_�ЀlzKF�
RZ#b��Ǳ6B׿-�І�Fy�R��lh�����������vs�@K�����Z.�沏�x[�Or�`7���a����R���>���W5�y���B8�Y�V�"M�=i�xX����M}����:�Bm��3�eM������ƫ��G���Q�.����PǸ���ˇd�����[��v1'�j����(�4
9�{����3�q��5�~�Tq�����0��B^���-?�%�oYk�H�I�	&�Z��e�b�s�2�δ�ɑ\b�d��������>_TU.����b����v,��a��bZ�^�k$�Fֵh86��yK*S/Dd$�z׬Zw�;W`i*k=7�^��=\'@��x��Z�@m���j��2�H���\;QQ�@b}��{��+� ug���3�u�7�L��Z/K[H'�DЄ�X`u�l�)�!9�D�4�U�I���2����,���W������W��=��U��i�@dꭆ�#�p��t|��Q��[s٪/��N�C�")\��ePi�#��Q�g��S�Zj��|�B�ABr>�z�\q�P��H�����%�ОK���^�A���:�4�`V��������_7��ksć[M�=&~Yŵ���$M��{D!b:�0��X�\�A0������\ʜ�;��"۞��tr������R>���5�;�������|MId�Wk��w�����&ɻ�o�hm���`}UX��Lm�\���yY��d�Z7<\v����o�q$�u���&Z�Wߤct�>3$�1�\ZB�㰌��l�����Yg���6]GJ�^��� 2�/�"�vbY�a��<0��!��e{�ӣ��bP��mO�l�-?pJ�u\TSh�ˡ�cJ���_�t(�b�h�S��!EA	Wi,2f��6��|���uaA������O���l-��~}( �`:��?J��s^��	��K����}�%��Wr;��kG��)�6�>��T�?��!�-)=T���QD0��+���W���e�lB��?�+�����,�����ɕ��U��`�oŹʞVH���e���t��~8�e�}���j5c�F�L��z�U��6ٷ�U��"P*��$�M������75�&�ة;8�M��g���Y�1h�z��6�\�d!LyW�8v���몇s�vHI����֐f��j�����D���\,�<�<��Ș �R)Y\�0�"u����!�=���Ǧ�A�B�/�
��z� ����=��-40*?���y(���s���(�����>�R+�W�-��n����m*��¾Gu04#��O/����j΂R+���!���<ip����ܽ��ݿ{�L�DUMV|��ȝ����#Z|��S�>S����i#�0{�R�}�P�Y&m~����2^�2����4s�~�W�L�{]N�<�SO�Q���Z�S�"���ދSl����e�>�`Ure�A��	��̎���>!�dQu�]q�-7���r�y�f;��͙��!��!w�W�AX��v�R�ku@�+M��{K�aqD��7Ҷ � x�(d�f0K�6Y4�ͳ1���Gк	�� ����NN<��y��^��εªp늻�,�P����x�Ge�-�"X6�����9�O��I���4��("7ˍ���I��Ky��^f��+Swx��3O�%A��,xJ���|ú5Α?@�ɱ2F��N�`���r�w
��͏�v��J��u�:���Հ\��ޗ��F���3q�HX[��l~��\!M�xz)�!��NƉw<�5 A�:��a�;m����u>��v ��B��c�Ȫ�O6dA�u����͟t��Û�+��qP�
aۗ�=l;��,��k�����^�z�r(�%�.�B(��^9q&ͽ`@61�ܾ7�6��=B�����$~N(�A��T����!f�W�c���(��诔.M"3P����G;a[��:�����ܰxM*��	�]��@Q���*�����橢8��C�3{G"�P�K׶��>C��sz�kPǤ���S�Nb9�|�Cˋ��0���F~M���;N�>��5k�n�A�z����l�I~+2�3�U��ƣV�EpOR����`ȵB�e�*�o{ǆ��}El5y ~mdK�0�l��W>�����y��ޭ.���Ӎ�B����C�Dލ0��S�����ַ6!G�ϐj�����[��8���Y!��b3�I�<���x��������:g�N�U�)�#�p�,�	Y��ڭYO����ɤ2�16t^J�=�� 8�tc�ԭ�-�w��<��s�A��ZV�^�J�&����G���k,R:qG6JV���z�(�>~�� M�~@:����j҄�` ��SL�����E5��p|�">�Է}=�	��zE///�N�?羶��x�1���*��>##$��C^�'���~�YD`��"��2��%��?���n�3"�"���^Dw�<k~�lmv���S����
'(�6Y��ʮ��KmQ��ir�ɳQL�ŏ��9�Q�q�=d흔��W�p��q� �4�'\*���r���A�:+>��g҅�����Ȍ��K[�A�[[e5(]҆7��ӵ�f��
tN��@�(G*�^�g������+���e�����H1���S���p#��:M�V�������4��G�1t�e����tZ:U)?��L=�UF;�/��].�ʝz2Q_�l
��	�"x�!�I�n�4.9����+��e���V�+�����cq= *�/�u#)ߖ���`�W$���$P��*�?�_����/!9��X����v[�
�����)���ל,��t˃6?��K;^-��:���I�U.�]�}LZ�Y�p��ܩn�}�	���r�B`�h�/sIA*���
I!�	��'�;/�_�㐟���O�G�p�4'������F��T�u$<�ߚ�fZ�cW��{C�b�bޤ��X<�k� @e���g"�X��4����Frh~��O�6��W�ՖP@�A8b�e�5u��n�á����(X�Z�j!縊�-��M]����H�=iX�d9�ive��=&�8dB�ib����dC�>ڊ`���b��Q�R!}(���l�M6�i�G���8Ղ���[o�|�%O�%'EU�����~�C>���d�h&h�id�xˋYd�����V�I�1P%��(��̜Y����_d��PD��k�?��bTZA�Nv7�����D��ʡ'�l ��HMrZ���M<]s���%k���N,O>EgT^���7�k��@x\��Hg_�ɭ�A��j8k�^ɑ��`M�ɿQ�'�=�gQ!9 ���+�� ��d�Z��ŧ=�e9����|F {��J���]��e��Lԅ߽�^�����&�ie����^A�]?^�C�4��Rqg�NmG}'�D�����Ё<}_H�4}!$��;��_��c|�i6������ Z�s.GkK��j��@_J�B$�G�|�[=ť�[���'rJA�c�s�<�ƃ�_�c�}���SL�e����MA]]��K��GW�S~�!5�2��e"�^n4n/k�{�z�X딙 T�`r��