��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܫk�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��5K�z��!��[��S}Σ{$Gx^����c��ƀPfƆ��>ţ5��I��xD�j��!��(7��� Ķ  gL�<> |:`��>!1%���Sg�M�^"D$Y�
S�N�S�C�k�܏��T���滀ގ�!-PA�t�`�Q�0������(#��g��ϐ0��"�k9��?�<��F��$�&��"֪t}���6Tə
�ٿ[������?9�&CFR�̓5�M�E/>�[٪=��x��l��\�'Ö���]q�q����`(�g�.D<�dV��϶�qLo�m����2�J�w$Ӻ��[��M%--( O����ì�As���uA�ldwP<q�|�!�y�[KB�	����̵nf�1��a�bעt���D��:��L-A_���eە�A�X����0v��)�!o��y�l���?�������Lwj��V��������.��fċ��7A�b�W
��0�o��=����s�ht�!��<��;8}��<-�$v�MpA3ShGg�T�����]����D���A~�������3e��xd�8!I�5%y��-0lvqx�Hb�k;��:m>n���i�o(���C�������"��j�P��/`ei�`|���d柬u�D����##v�*�	A<�����hܠ(1.��˼���7�l�M�����U����&��̖���+H�cZ Bl"M8�/f��m7�*�0�]|�iQZ>,Jkn|E!~sE���Z�b0�bmϟU9k½2M�cv>ɭ|��h(��,���L㝏�T���Eؙ84�o���=�� �k�G���V�o�5{u+���8Km�U��{�=8\�l֏ zJ��$3ـ�����͍#�z��C��~��V����>ᇻ��TqU6�Ю"�Q�QL�K�s|A~#�TM<N���'�7�/iv*_$�xO� PC/AZ��	���)8�w<�N;B�G��#S��9b��vl�:N5�Z��&�U����>F�ml�� �~pu���F�i5|鑨Ԡ��m�c��=:��46}lf�\M�@>�f��V↣lӻ�VP�a?��ōӞ�L���mb�-��������~�YdG�2(�&?�!@��g�5�����Z��r,���]{4�^p���=�Lx�UyJ����[�U~-�ӿqK��ޱO��� �@��M#b`�)i�����v�g����;��m�u옌
MG����`���oC���Kوc��N	,F��=��q1�[�U����ߗ������x�s�Zzt���#�ܧkX6�f{�+	L�幫�Q.���Xԑ{?a�P%��5�g�f�~3�ֿ:F�����U��~��҄<J���`m�0���	�����V�ܨ�\���ns���_6��b͞� ����k��o�<�0���!�D5�f�(��O��={�y��!`��M�4
ڄqJ�VDPЖV�BС=��A8$V&�rn0΢�n������ө�����yOz���(��=��2�}m�U!�va���"�B�l�g�%�
NF�+Q�#d��t��?,��T!�g�T���'AV����W�Õ*3�e�_6�y��Ut׊{��dm�Q������`�VⓀk��DN�}N\|�%5�>L��i��O��C�S/�7�7�!���9|J�s��jT��૵���a��u�>v0F�rOA�V`�!��^���ƽ[T��phs�ҷvt~%8P�w�>U��YLgq�����C�:s�4J���|H!¿Q�2���Kԃ#/c��(m�W Qɩ���|X��JBNi'P�@g�Ҙ}0��I�l�C-��5�� -�Ӓ��:�� ?�e)g��.�	��c��G��n��D.��ւH!�/�0��o�9ӧ�7::�{�Q��OB���/�(|Ro����wI�AJΫ��&�ZmDˋ�%�'��;2d�p<���Y�2I�Ưk���>�.�H#�rƞXY8�sz@���gaB�h�}��5�đީ�`da5�vE�<�x�Č�5Ԩnr�{."��u?�x,��R:o�w�-���كS��JS�7҆GSFy��G�{R۩B����W�W�boǋ�n<�"6�`�������|��q�n�7Vf�O�*SUWy�^P[�d�F	O�Y/rG	��r,���?S��N�.�A:�(F���6��ŀh�5/�y��*�X,����C�8M�B^ǌ���St떬��q׳���i�i%~s�)p�)�v�M�/fZ��-����G�V�� Y��ԟk*��3M��S��[�ӟt�7g��Z,�/Vߣ־�ME�j����I���� ��h�^;��5Ǆ��w׿-7����Qh*C��j�q�DLq %d�>W�.#C�ߏ��Y���Y��h������	˫�c% ����j�Ȯ��{�MF��J($}I��+LcJ����@� �g�ʷ���(���L���?�M7lFJ�I��t
����`�#�1��!V�m1�"��zs11VM <���<��VƠ,�����ƛ��v�N��R��Y�%tq<:5W���@�h������Yc�9	a���\�o�#8 �($�3�G�?� ��5\���گ�*�Lrڷy��~�m�G�n���.~7��ps[�cUs�>꾀�!�h��/����c���=��5� �s�������S����DMEha�0�ġl$�����t�f���
5l*�uf���zq�|R������Va�WBu�<�j�f�4A��I�5�J��K���"��7����?�9�}�B)k�p�BC��D�V��t��C��-��WG�t���(�[�e��l�m�J&T�����DB�m�+��ÅS�*_S5a儨�ۺgpVf�:{�E-t>����A��	�kۮ�gڈ0�<�g��;5@�