��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܫk�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������"0F��}�h'��8��<���9���-�j����,W�_/�H: 2���x���CH�^�gߎ[�zZ$D�H�=���3�r�-�7�Y��B
6����I?�����k�'aQ=$ X[Mo�o�����o~��P>��]p�]�9��D���M�y�~I�ʘA��l%�T=���溟q|��iN�NL��zH\M�I���u��L
�{��D 0�w��h�g�>%����2��*u��ПmX��)����/�̑蟕�H�����6[_ �oY&�,P~�
�c��~#�	�5���6VCA�F�_/�c�o�9JW�c#�Et&�.�Zv+^l��!����NB��>��92�L�'�/i��׿�ؼ`�n��H�L4K�oz�H��~�W�Hu�KN��;��E�	S/<}��x�
��^px]oaD�:.~��:��hQ�S�χ���Y�,���/�x��qy�yjZ�ڄ��<���'��X��
'������D	��d�b�l����K��!�uĽ�L$�e}O�z�!L�r�䌁�NB�7i$|5��b������*�]��@2��MPG"FA��Z��ƖJ��zoPw�*0.U3�k��^�4����T��%I]3�l��z9	%tm�����<S�$���从�<�}�9Ң�r�'����Jk���MN��}	B[:�b��d%!Q����3p��xD�!���zV�F�{p��s�niuψ��f��"��a��e|I����G�[}Aw���{y�H<��ͬ/�dg��y�����2ʠ�ޣ�?�]
e���̀ȴ�}���������kR�/Eb����ڂߟ�wm����ϱtx�)B#��Uş��ÌD�޿�<�$���
S~<�n�ZVؾ�F����Z�����m5�K.���w��.���9�ބl�8��+F��f��F���z�vW��T~����F��8�����.ˣ�4�0�Y���G���,^`?#�F.�2'��]vl�P���tn��3�#����i_����(�3bͳ��\�+K/��5�L�}����Gv/|h$�1�� �^�k�nq���h�-7TA����[����<k�ib8�KЬ�3�r��\5��.b�֯D7���͋3�n�/;�|:0�=�2![g;��tpOZK��=�vE������ъu�?ĤEhsC�p�z�܎�WS�n��̰߶����\8�CNg$޳�B��P�-�MT�V'�7�ےb�D������mU��0E��O� ��G��K�xe_
�u�BV�s�b5�+]̚C���-#��
a ��_$%H�
�{���V=Ƨ�=�M䙣���䆌D9�ʩՆ
�.)�w1"��zT �Ì����z"K.��
Tֵ��^IJ�\b9Y�n ;2�(\k6�I���~�H��Z5l���%)B������
cOo����hc�5��J�҈����X{��5;&�&݈i��S�K��p�>ސ�S�æ�ϵvzۗ��9Id���h�w�_�U$�W�y�Fg�ƺ��)�d�.@�P�r�W�у�KB]�/���x�����=k�ۛ�Lf�SY�XS�]���w���@d���>MBt����eM�s	ə ���y� #�l��1#�}z�'���G�_y�/XW���|�KQ���}�(��/]Cs�C<&6�g�@������cŖHbO���`M�u�L[�Yr�.�,J[1r;=r�^i\"+������%=3��ޱ�!�>J�ƻ;�x��𭘍6g���D�GQI�yI�Xjn����t��ߎ�Rwt�T�u.к���g���%�7(5�%�@�B�x�ߟ���X*No�3m譮so��N��	cF�\]5�� j��ǖ�F�Gm}|!���s��]e��ח;s�ӟ-�����0�L0N�n�a�g���j$(�1���`�c 2��� �B8��A{4��_�J�һpDӐ�=� ������I���]����SУ��IMzI�S8��'k��I7�<Dw#�v�|!�jy��j����asS4i�G���w�<P`Ȯg�|�<��(ӳ������I�R ~#�ZkH���Pr}�8�5И��d]�fP���ZG��~c�tQ�1����I���������j�J���$06��tH	zC�9[���]��+}Yr�~%��7�S�!�����M�1$x'�,Ym�\H�4ߗ��sz��Y�{�]
���5Z_�e��E<�=����z�gz��g������%��؟C��'Jf��ͻ�I�S:*����DK�����p8�p,�<�d5s���'Gˌ3����7^��DBыZ�6s_{F�&dvP;+	c�φ���`�k�Nt�H᳦
b���E��F�+����#�N����sx���6ם�	0!��uσ%o��R�b����C~ʐbS�~��\�R��$�+k8y�mw�8�|��.�ծq΁�W�z���8Q��?p�l.ì�a����ߺ�x���?ܔZ u}�����S��%Bp�Rt�aar#p�.��G�<a���Ay&.b�s"r��)��m-K��ܛۗ��4~�Z�#^�S�eM�ś����˪#���IYoB��1jF�O2D��i��6��$�i�FЂ���.�l؍���ϭK�ۋsGe���|Z�Ⱥ���?�:,�
��������������Or질���)��߼�j�x��ս�33@O�z�j��4)��:�ȓ�t߿����~�/��J׃[�S�i�0��IU������}/��{��D��%&��C`�*�c��.@��cUnK�j��:1�k�a>���~;� �l�"j�	��!W]%���WsQ�?
W;��Z �CgC�n��c��;#�r��4r���!� �	�C�qߨ*��V��W�[��O���W�sa,`��C��X������?�h1VB� ��T�ٛXU�;����SO�L[���N�}V+���^r�Z�?�s]�J�����)̵b7F K0��	����)��� w\�\Ah��(��FN�u�lM1IP�v����+u������� ���V�[)[U�@����qH"w���Q������.�/�ab�|i�F���D'�b���uC�.0!(���`���X�.%�E3ŏa	!-��,�ܮ~���H�P�s�Ps'�����[�%q1hL��@=F�#Ep���z�$��< \��P����$��Ѣ�������Y^E��;vE�`�<d�x���#+@��+v���O6 z�
�.��1"�y��?��ZW1�$Q5�\��c>�E4���i
�wR�;�e���SMkM�X��2���<�p�����`*��犲���W��L?v*7.��ܫ����Y�v6�/IUn5}V1���1h�uۉ�yV�!E��2M+�t�.�c�ԇ��(qoA9���Oa����ApC>Tb�'X��l����]��N�j�f/Oz��H=}Ÿ��dH�o54 � ��;$�!2 ,�!��h�,��������l���0 Hڞ1t/�d�JmD9:���>2;9��w���p�ȧ��V��N�HPo�$?�~���U|P]|��4]?�^�LCg>���E'!V��5�g��<�7l�����W�O����q�Y��m<N�R��^�۹�;��穯#.���$ާ�i�B��>�9��d��m5�������m����m��90JV�΅ᣅ
��@��l	�M��yhF�{2��]�q�}(���*�X�u�K��=0.ԛ�A�Q^�v��~}�
+{qA_5���y��n6��њ��1���5p7%�*%\ϻ�<�\+�R���4����q�8�&�uUX(#�t�qS�=6�I�����mЗS_�淾J[k�G�
�[z�Z���|� {�����*��]�6���촲�n=�2��Ke�8}t�$�8���?	^�m�;���d�����bfZ��sN���|��K���*N@�/�B+#?6�YF�՜�/��������!z�����O�Ђ2�|�I�*{����̥��>[1(�5�{kƛG���e���p�����o���-���x�Җ�|�Q�����`b�F��
z"��L�6��U���G���@*��0�p劊�؎��3lVqR�{�k-�*t'�MKl��bU6:5@��sʥx<��L�����?W�$c��ˋ�)���'�H�'en��<�j�9�a���$,Q�QʇU/��E�t�P�Ѧ8��(�G�i~S�lN3:�%�����e�`k/-:!$��]����as��X*��a��΁���$g�^���Yr>f�o]M��>n:�e�z}��r'��݃�rs����y�pI�VS�gh
1�Wֲ�o)c���K�L���]��b�,�9��"­�cn�J��;t^�:O~T��H�ͥ�q� �������$z��8���x��%�ħ�Д�]��f�cG&�}��U}�'(����1�>�-
���t�ʧu�-/���?���O���eP�cc"�?]��Ы�{?�����(;�߼cv�a։O�ڑU��hfb�dFhʴ�q{�UJ��WO,�&��w|t�Z���xθ�~ݛ�P��@U|cU)����y'�NE��d)̡5��8U$���`3Zfx/8�	����G�Q����P��BNo�Y���{eO�Z�lX���m�Ş�Z;�f7v�]BCU��_��	�
�8}�P�/Gc������i�p��P�QnRk�d�qz�xP���T&�]ڀ��u��ɀ����Aɨꦆ��
c���M�Ҝ�Ƅ�V6���H�?�&�6�x��͢�uFSá����E(�+�x�o�a35��:$a��]�Ų�c�5A��^�I�2Se��v_������K�=�,����ڈ+��@;�w��~/ޘT ���0���#XX�d�npv�
�%���������o�%}wX�]KK���u�7������q���_A�������t�U 2�D�48E�gt=��<K�z@���(�?0C���hV��u��X9��#����ע��g������ER	
a����z�*�<�j�����u�0>ӟUIӳ���(�|�oc'��i�z���W��[2��g���:��#>�:b�d�OW�H���7d2�XXs�bV���lA���A0k	P\9~Tj��];�q���#g��nj��
��r�a}�]S���N���ff%��>����|���,����V�+�怟��°�e͂���K��)�s�g&�DosL��(�[�����d��D(��X���ͣa>���(>�@�r��t�S�Kp�K2E�?��񋓋�`�s s�(���g!'���F�!i���*9�Q��;�����<�pk#U?{(��'� �T+�P��45��.�Ǐ���LR��J�Q �����J����ڰ&,N7�;�/��.*!����_�D����tE�l{^75G�^-}��֟�3���j��9P���b�$5�Ji.*ZdY�" _^�^�#2[
;�i��*3��J=��h�u.�||��_�:բ��v�t��%�PN�q��c���H��b!�7�l�յ?f��D��)�hx�C
 �3�&h�m}��>\�Lo?q\�Zi�ꧧc���8iVL?���Ҧ�EDح�����О y��\�U^�KM���=�$O�1�[W�r\h͌��% @���h�Ȟ\UXG����!=�c��X#Tmq��-��˅���qh�J͞య
����b�Nz�+��
I�8�����#�C2��w��x̕%����FyoxƎ���~,�\����2���W�y�uQ�"�|k ��ZU��*�:�ܑJ�	\-ׅ�v0�b���C�>F�)��R�ȺJ�}L-�Z��)��AIA¨�w_��`�����[��OWt\�9���$z�r��e9e�i��L��T}���w\��ԕ�|�F�.�7��Oջ�h6<�p�����A�g�?8C`ֈh?� �]x̥@�-�oy��v�M�
���/��j�e6��	Ǟ$t�˅���UAV�cv�stZ��P"0�qU�65�']�{\��\�O�c�mRY�~U`FӠJ�pi���e���_8��҉wrKR��g��N��z$ӹL��ṟ^��#��O�M�&��x&���8����K�� ��2:�p�h��A�K;#%���zEL�N��?�1�x��D^�r�{�/���OO��?m�a7��<n+#���W�4�����x�=���|^��.�z��=&.jxsjw�&b�/���YX����B���2�Z� ��J	���'*�$#���?ţӡ�l��P]�T��䕿e�/{p1���~��v~u��f#1�6HhJ���\�Эƿ����ȣ�Hy�v Q�K�#4u	��,4l����l�$쨝2Br�	�&u6��Z	���ݿ��0MV����,xbn'�_��ϗ:PI2N�U���
W����ۚ���g������}������^�� ;��~�s�[;�vP�5�4��S;縤fy��/1�\�@~���R8ݽ��[�;��r�tk��NP��FA�G&������^���U���$���LE�g~�{PA�ܯs]������_
mW.�;�|�-������ -쁊R[uxZC�T٦(��A�Q�@Uq�3�i~9Q�m;�`��!Mfӽ��%:�R}��0)�7���YE�54����t�����
����{����J�XE��)4y�����#��c���)X��ݮ�j ��/��i-_<��%~���X�ԘUh�S*��~�=�~L"�&�����j�qa��B�)�ɦ��#�Ӷ~%�������uUS:u�T,^��*�d���B�C ?SS��Z���Y�h�z/O��o��fgl�o�46�O!;�b,*����U}(\���ݽ/(��v�+�r'��S|�uX��/��t%x��BVX�S�/�xݲ�y9$��5M����:6���Z]��^�n���R��� p_���j���G­�͢�`�5�M�K�p�{����l��z�E�!���J����HE������^-��x�@S�ո����|~���
�̓�-�MT,�L�}�D��"�(/�e�+��{$��8˧�������wRK��ާ�6W������E[�z�J%6�r#]�c�q�6��K�kkt���{��u(J�)�{t�,T���x?!S?@���.b��~˖qE�@��������܂Ѳ�/�����b�����Y�+�
RP\�}D7��5J!e�L'"��G�Lh3{b�
0#�X�Dp�	� ,3��Ū/�������X/�c@ߒ�Ќ��n�3Uȵ�SiG��H��L @'�C��U�/�&s d�m�(�lX3��$���v��c��BS> h��iH������z�������#��� ;�����5FG+A���<ĞDB�����{jS?c�	s��+�h������:������K�������{ľ�{�,i7���硏O0�$�)�H7p���}e=��gf����[>̛f��״U���l���r�S�~"�&N���G[��_O%FSP��Iޏ��%CD��R��>+�Z��NOY~�c�f<c�m�h��}������uYU�3_4e�{"X��c�J&�T��	T',�� �n�HD�����x��^���7��#���;hZ�͒��1@�.���߆��z��r쩿�
�}g�v��B�$B����(P�n�o��
�������!%�bp��2�f(����7N�`ࠅ�n �h;Kn�-�-rH�%��i����*�\,�ʊo7�+2h�nͶexV
H�iX8���[�T������Ǩ�}�� Q��/�,����
�ۢh��#��X��g��%�����v2p+Ch�>�2|�g�:��s'��j�����?�0 c3�J?�/��?�1F¹dX����5Z<*�u_��P���F2�bT��D������NP=_�i�"��������73���4E;_��h��_�np��m�/>I:��m��3�?{,Щ�<荒�aR	��-�#��?��2DN�F�c�m�{�M�|]}Ͻ0�R��6�R!� �X����;��E�?"�,���e�#��j쉟� �Ѿ�3���_�!�BM��ls�H���������P8���Q�8��y�>��O����o�4��,�x\�BѥX�u�o"�G�o�r�A���4%R88b�ӷ����+�!4�3I����.��`�k��&A�4��Ķ�L�*85���Q4i�������*st�rǴ�6�F��b��h*��VC��ob����my^�b��,�M4M��u��&b(��N7J�&��N��ÄqHP$S����e�D�q��.%�W�TH���(��tb��ν+F �����u�3ogQ�a��#(��
U�#�أi�� ť�O�n7�g��c��Q�d@�n�JGlT��O�R)P����c����%*^�	�|;�  ��e�dM�Y�a;}�pA���L�3�Hee���L�<�.}r(�
�ܢR��l�>���+Ֆt�`s���$������8��X>���1 ����\z���R:v!�`�<E���

V��ƫH���^�����l�g!G��"�;ߠB���c��l�E�K-*���m�@B���fA����fctx�ؽZ�� �i'����,p�%�/ry���FH�P���#�9�p�2Ԕ�K��41�L����@�'IN�	3&�v�f��R�P�	��#��?����:�A�=7�����im��9.�e��3�c"�����E����ޢ�h�:��\�$?^�m�U�޻j�Rq���B���/�$�>���)��b"V1���n�r�^P`>�`~���	��0�J� #6H4!�ܮ�ۓ�ōn¢�(��tW؅?IwP�,#�$܌(��)��P $5ǍO�WB�r���u���17a���s�F�(��1��}�"*d��[�MI����K=K��K�s�`���d{1��&�H��k��.��J�nޑ� �7����_�>��5$r�u7��BZ�N�J�]��)%WBQ����k��7ԅ�5�?ß9�ȡ|$�C�Wt�,����Kk&��6�2	OK�w�U�V�,}j'J:�AvA��^�6�x#)�Q��r[�[�%��K4L�~�*�ҍ�b��:���Т�15T�3������ �ڌ��Ͷ�.�#4��9'})ꖀ�#�����@�7/�ϟQ�b��H��$@��X�k�g��X��0�D��� wYF�\u=v0�+�� ����o�c�+W�!k��-��l�MS�k���>����~��!�?��]�	Pu)�H���)�R�I�6���{@�_ۡ�����7WRL��? D��q���֯�zSx���],��Z5/4�X0a=�r�e�e��[}�"�;&���:<}�8C������K�.�Փ�4yY� �}
�%�᪃2�"34kBh�+Oﭽ��5�r�m���0�����;�+�?���Nz+�X�_Ԉ���tF��P*«:����s���fq�{��ѱƇ@�]>\ldi��K������ܲ1�rѸ�$zd~�EU�ʁ�w��bтiS��V/%�T�2�ql6�'zo��%�F�����
�o��,5�kc�_�bJ��O�mĖM*֪�hC�4dMcW�P�տO�"8T�w)��Ⱦ�̭�{��WW��gx-��96�[l*�R�GwA��oݡ��,��f>�o��λ����;<^\�Cz���3)�43�75��k���!R`B�U� *�r-��v�l#��-�[Ҥ�[��؎I$kIe�:�����{��_�\.��]��_�
9�7�p�Jl�,8�߫�V5��H�
�6e�eUYk��y\�Dk�"%�<��*�N¦'.V��P>Re�Ȃ��ƹ"����M
)"@R�M{0eK���+����Rmd!4�����b<���f�I�6��ZNl�
�{����W
l~C/J��v�&�����ƽ�	��UYoWw��='�]��"�_� ~uJ���"g�c�J;���M�Jj�{P�!q��λt������+br�U)�V6���졯k�2JZ��� ��}/�k�7:�C6ZJΩ����˭ZXHS�4]��a���{�����⯸(2�.Jq����,�+%@��B������"I�oҫ�:��W���M�,~���Q	O�T�&t�K.���mh���z�N/��n�c_��^Z|��,�}0�>��$�4
A+��(Û+�>F"0^��#�C�	do�|ݪ"��X ���H+XD� 3��^ς,b���k>�k��\�j�V�\�8C�$A�|4�m�J�;�`��.����8��V����,� �Rʈ1�s��Ľ�B��?�h��,��X�QB��X@d:��^����L+�& |%TnVO��l��y��q�����wS��Pt��醅������U"��%wC>���v�h�D���u?����CO/V������E�t�$�����^P:5���K+�hM��t��r��������Mqe�zHi5m_�x���!����
~fQ̕���,\qCxDJ���۞��Z"UYwCѸi��Q;�qh/���o1[�c]�I�C*�^��s��,.�b��2�[i����Bgu�����sHZ�E:D�L�Z�b8�h��"R�?�R�����떧:M���ҟ�����
��F��(�c-��y���v���!�l�u~T;(��U����6'��ܗ�mm2�}wH�����H�z0y����}Ϗ�|�.f`����g�ы0b���)�q��\ ��i�[��	�/�%�������J�޼\rq1��^m
$�}
��2�s��c�W�w�2`I����#j7T������5>����~7D��_�zI3�W�Y0��s~L(E ��KWOd]4�b�ĸ��c/%wC@���ی~�Z)n�%��6�`�蜭���2^kv�!����Wty{�V !��V���꥾�%.{#j��+��4d`K�w�PȜ,�����^����Zi���3q�E�0v.;L���!��Q�_+����c�����e9�i���_�pW�͟��LK�?�U����V����G�1:o���?�r�0�o�j�/�#�v�7PH�eq��GLt�
���:�y�쩺�x�P��ł��Sz+q�����d9t���3q�m�w����q�'ٝ�Z����T)C+��/�l0r�s�Z�>��#���˷�̍�����!=��Xݧ"�rӘ�ʒ�ʁ�6����˞��:�&ԃ`3*�B�<}�~k�6Ɖ��(. ���}k��T(��O�TԬ���ՕUUc�?���<�Y���T�H|Tp�c�p~�}F0R֙=փ��B���Ͱ4抱��q��YX�AR;zp���4�yB&�/S4T�D�07�m�ST�[�������_Lq�6�R���^��Ч�>����d��H�x�3W�.�~�!�