��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn�%�����݆@<���U���x�ո�y�4�z�Ջ�߁��@�~�ә83Q�f
m���M BLs�B !`	i�l���@#O,D]#GΚ���|�4�[)�qm�r���Hj�e�Ep��V �^ܰ� H���l���r��65ϥ#^��/1�ۿG^���;"��S�5��M��A\����� g�ÆČ��&_t���m�lo��T��+��X���=0�"�ԃ��Y��6�[P��~�E����y��T 5���
���Ў��q�g1�|�eX��*&N6Jr���������U��`�A�� ��w4Iq$X���)�	#�%z;�/�y�_�$�C7���T}������f�!��L���YQ�q�dy]�E���fV����nõ�����fݏ���ӼI�ܝ�'	��w��}����������Q�Rj�ac�0/p{���R=�j|g�2F���Q����m�8{q�Hº�f���_�+d溸��?~"�Mw�(��1/�����S�4�j��q���Hk,WJ\k�ߡ�z�v'�L-���R�ŧ����c�V���/���D05ƞ�蘮�|�eNjm�,V� Vc���:��BƦnΦ�r[?��������mX�����-�'Uj��R�J�#i�VĤJ@�7�~����!0}z�&;Q�E;a`\�I72�+5�dzI���;��n�tA����l�fTR�Q��1�A~���8a�f���\3P�6�JН�,��V&$����׀uAhJ/a��p����#b��G7;�k�ç��g�S`����:���-�M�\v��A224�&0a�* �Wq���>�t\���|Կ~5�$#-F�<s0�}��^������wD�͌���Ǔ�A�ʘ�ɻɢJ!7O#���)ℭc��w�"H�,�0>���Z�~�Oq1����@�>������¸�D
����$���<wA!^L�s)���{��D�#�#�h�^� ~Yz�@�w��~R5Qj�m�`5�����N��Ȍ�_G�Q��Ϫ�3U�Q�s�F��&d�_�>�����c��m�&����H�@�l�h0�W-��j�Uzpu�������GM] u2�&'�c��d�Skt��G/�S{#�Z�Id�͑r�����r�³�
.`�{�딯l��ΩJ?���\��X�QF��Z�� �F��?J%��#r�`j�^5�B��:^���9 e��$�w6�����C��s���}��8�bV�@!m��CJD{RU@F��ї0q�b����wқ>[�}�*�'���2���+��}0��(�-�������-�+�}��ZxCc��ڰk݌,�&"����ࡡ#h�]*�� 8�#3���>ޖ��o�#M]u9��S�
�r:� ��&#{��Y�a�1�ZB�X�#B�$����>7Խp�i�B+�����l+{�h�pg����d�z3`�;'���q�C�e>��CLr�el�r�`ޝ�
��3�8�����>��[�kU����o�.j��fR�w�����]��a��B�/�S�?w�ζx��O׊��C#j'8���X)�N!I?�C��E��t��Doc��`�|*�e���))
ġ)�M����ɚ�E�['	|P  `��
�G.��u�tE��`X�+̇|܉���S�)�'<������h��QPtۯ����%$�	�����c����K����u�;�"w�N��Aĵ�=Rݤ�5⸭�W�K�nT��� �޴��s�0彃�T~�L|���Ԃ�O�)c����!�D��tȾC����&˵�3��!z��<�>�C{�6�H����ʛ�_�J�h��)ږ�A�%�[S���h�jz-�]�o���<&�ջq8�Z��KX�ZҀ������6�.LE!z�'���� �b8ߊi�#���9�M<|ѷ�5��i�1��S�q��������GL��,WT���!�o����`�حi��q�&�E�D��/��e�V�#�;%FùgX�!��Hj��k��ЁO�f�	#n��:N��D�}Pe�Q]�9{l:Z�&v�W���d1�P���I�r���h��dtO��4�֐
�w/��Az�-��}��/k);�J.�bO�Y�ŪPj�z�r%����0+yHJmp��rM�rTL��|�!ڛõ,�ǭ���y�,�\u��-����d����'q!�vz�ct ���tO����I�v��_Ʒ%&���SD�U����h����c�+�4���D�7_l�>��ãtV�S*4�̿5Q�"�ދ��{wV����~�ܸk:ND��:E�2T�}�aJdߣ��+
�F��C�EP�u�4T��{�H}4e��vC��b#u�h�Lq�uj)A�w��bi�k���Ĳ��|Bq͸Яǖ���Cd�A�1:0�@B�����0����si���XP1A�D��l-{a6�r7��1�<�u�	�k���3��*���q/)c���AшI)�RB%L	�U���δ�j'�M
�9(��<q��+�Ah�J+TtRt,*!�MM���w�����`+Z]��BkU�����J�\FU�|���Z���)V�;��*������C��a�A�ໍ.r�j�L'0��`�U���;�S�9Ό_��sĮ���s21��Ūi
���n.�K/��L'����C~�� x��r�* �g����❏�V�E���N�1�C,L���(>��ll�M������1R��y��l��;�OD���HM �����C����<�QJBCZ�j�'�	F�W�X��@Z�L��Q��a��KGY4���u'��R�ΤLb"��X�1��'�&���D"��-;�:�i��wf�	=�=��&hfW<�dO��遏�����lMwǏ�ƪ ��D}J4ɢ&����\��f��u�����k,{��L|�r�T_�Ϟ�k�9,��	Ƈtxf9��:���� ������o��gķ�I�(ƛ�<��Y�� �U�� �]�B8A�jT�HvN�9�tb1OO��*�c'cm;���N.���9�`�c��m��vM_0-؄ID����e�URO���;tN��N��M�a+�%��q`�CB�D�e_*��4��`�����w�B�.:V���$R*�T�
�L�n�v$TA��7t�}?�UV�]�/5r�/U7-?Q��*'au�!��R9�*xE9��ᛕA�IB�c� �%�uB��HQ�qK�z7pù�L_K���M�oU�u�s�?��yv6�-AE�+�C�O4JP�Xp�M9����pV�;�t�����������Q�z������)5PA���r]���d>L�u���@�Ⱦ��7���6X擞lx�S
~[ܢ��k&;M��F�L��!���m+�#n�����c J��G�Z/B���ڈ�j������cc�e��Qb�@u���Y�ՓJ��
�~��U�\�'+Q@��W�]چ��:�?�-���v4
۲��~�1v0g�o�5f�C�!��m'�r`����zjl�h��}|���z^Z����^�,���`�lG�pg�������5[$	�J�
��q��$��)�+���r��#n�N :�j�>�5v��7ne���)Zd�T��@ў��E%^�:}��=g��m@��+��(��"����Q�(���n��nuF+'�tL�B�r���5y
�ܜg�S��B4�c��9ʏ�qr��5'˵���X�\r�S��6��h!�b�`}��C��F���1梞M�!��
�XD� `�P�����J��%7hW���3��'�,?gJ^ ��?\����h������@��1�+��:�AO]��ɔ�Vc���
�a��"t�ӵ����Ci�~Kg��~��y}7�Ɓb8����E��X!��x~��	I����J�Ӏe�B7��5�<�&0��Ɖ�c���p�؅S���77x�%U�/:��3[��$}�li7�W
L��7Q؇�i����!��ֹ��o��Q5+���yVߢ����q�=
�j�)SZ'����Ȃ�R~je֖��g����h�{��T�Y���HHqu��X�VJW�.9��y�4o'�0�e���nP+��j�i��u�4-����>L��.XuץɁ�]�	2H��?3	A��b��9��	���Gqx��,H�6���N��^��5v/�#�W� <a��y����BH��&��	%�#z�W�hŠ�������z.�\���I��W�d�[(v~e|o�%�2���(�Q��+y���2 `���	��ڔ>� Yhz��.:�Wm���6gߓe5��G�e�������a�S�]�C�%d�\+�� ��z�to`�ܛ��?n��3@�Ɠ�{�G#+�b��l���	��� �\�0.K^�#L���Z���}�@�+)-JÜ���	똜�Dj���/<��&:[��ˣB�K*�0��$���ڽ��&D��agR�v ���`]�#�<�ݧYC�����\���m��Ӳ�o.{9�!$J�����ug1#Ԝ+:cHl�����Z��`���r�#�Ӣ�HwN;|_�\�kŧ��1�Xy�jN�}�W5��d�z��v��yNe�+�Y ��k:m��dM���kn�o9������"7�>bk���	N��$z����\�08�AW�~6���u����ߒ�1;f-CKu;
WNk�۩���K�J�K2��Q���0i��E#a����	�������d2n-؍m>#2=�X*XV��M>{��"A�����0t3IW��)�;]�_�o W�(`[�o*��5���Ј��fb�X�Fo�d���w�?�rn:��>!ar��4�~����K�qGJ�����;#!�bm�ɛF~ވ�<���ە��"�Z��*�5,�/�-�b�h�:�u9�:*�S��۶v(� ����0d}l�lW��%�(�����6�ri�n��K!�a���p\7$X�� ���>���i8����#�C��x��c�u�Y&��������}̓�W�x�ah
c�S\�pL�,��@H�����е!덙N/#�64kE����jV{(e��@А���M����ݸ2c�?S�=����ͼ7@��L��s1�1<|Dw�H.�ݸ�'��C�A�Z��;a���=OFN�\Eb�,����=H�l���"F��/������P��M�����tl����p�M ��⋩�A�6*�Y^^�i*�:S�<��T�}ww�8�Wd)�Pn�-�nƸ�A� ���:;�*�n�T�������r��ك~�Ur��Y@}6�+�>��bx�����k�a�q����o,�"�]�����s�
%Q�H��F����雡3��G��o�돓T�����8
�8Y��cB��c=4��m4�I͑��o"��mx���K����/W9��/����*Z����O�ߑOw;�Fó{�c�ZkʆGY"���ͣ׆x�O�%*o$j����;Ԝ_D�3��J|enV?��l�X݋�-z��0۳�a�/�-Z�qx�K���whY3agn���=ı�i�������N.E �8�µ�٬(5S��z�o"߃*y�$��h]����ǥZ�C�F�=�u����7�w���ϱ�3����le[XB0���p��'3���R��?�WM��=̼�c�a�����Z��Q /ݜal)�_oQ�VR��σ���P������4�y�K.y�\(���K�&W�p���X�C�4�X=�ba�bz���f�v��#s0\#��7�5"�q��3����.f%��������Q�n��G�!w�q�NGuL+��#�`��a�B�RE�������#;	�	��oQ�J��B�DHN��^�To�J�̬��ԇ����6i�p�z�Y�)3����@\j׋���3��A<k���c�=�d�;E�'�]��~��Z���jǑ�|�@���t[�^�����Ǹ��ayBһj%�O���P��ԩ_�j|2��Z��>i�؉w���Wš���b�f��v0T�IǚNxk9
(-.�����=��g���eږ�\�4:��N�^�A���θ���n��>1��9�|�_i[MQ�> �b��%,�8q����!ti���oD���!�Ĕ����6��N^�D��Q2����6#�iq<���nk�)�]�{V�m*"�DCQ7=24���~w�'#��,a�y�{%�M� L��A��H��v�A�/���)�U���̜�	`��%�G�$N��'�������uk��kJt�$��8��X���׽�n�
*f�����jN>�ȗp�����F�_ᢡ|>鮗ѹ*��$ps2�������ף��8hcO�_NU$��{7t{y���z�p3.�?�<Im����ˋ�J)�������_���T�'�	���PF�z��WK�C'-2Ά}9�8�W1��RT|"Q��D���0�/oF-�Use��}�{-S׃�ɼ��4�x��"tR��2甭0a�����u�<9��Њ�}ߗ����Rc-�U��P)�!�.%�vp� �ڣa�
�rmyʛ�����I���J��^�;���n��l{-�؏e�d�wz����pI�K0���vc}�̶7�S#v,�*���h*�r�u��l�2��Ô��Q0���`fg�I��P����6�k�)h�޼���T!��RS����l�����I����F�L�_6���:��R�<R�!1��W5Ql�"p�dh�����X�|�:���8���I�̶�%�� "�+m6�*�+����-8oe��{F�3�L����IX_�;6���Pa/�̐A��*���A�1�A�(/����m+��!��/j��xە$��!���62�(e����� ċ����6�(:�^�����M��k�ɮ��ٲ�Q�$��M%�F�؛)��/�}2�4���l���Wi��
��1�著��f�nШ|d��{,VW�'�*�`9_����*L7��/C~���3�6n�@�O�mև�)���f���!YR����v�W�˖��[��9���r�:zgC_I��$OQ��r�I�_��o)�$&y��JN+'`��k�����L~�r�!AR���f�f�k�΅8-�?�,{�������)PL$��������Ԓ�K`Ry�cD萝��&��3�|WB��Y�C��_Z�kM�̩֏��c����jv��܊Z�A����e^���.����=�z���,V̈́�
�V�qy�?��B��BX�$%G�I��Ae���_��ӗ�	2�h�\�3�x���m��~�
9iAi;8%��dg�8�>+�Uc���+�I	��!�`���D4"ٯ��Y|x�;z�I��L�ˉ�e)�D�R�S��@�zg�����LK��-;r{�JU���w�4@7s,�q���z�Q.#�Up����D�}"�c��J0� -TA��/�L���k�1�{+�������K�5�gvu��^܆���ە�.+7Pe�	!G���d�ȩI٢���µ�q�w��|����~���\�z�:(�ڂw8o%��Z��'g<;n^eQ%1�0��>ky���D�<"�xl���$����)2(�s���q�C�(�Y:���oayg薕Z��l�;Iig
�����α��N+	{����G���	�n���/w w�\�iN�W~�?{�~�ЏHBZ�z�0�'܀Q`և������abq!�x;z
�(w���H�)�_��x���t-ϛ6��Ej�%�Q�*����ė�� ka����%�=w|�,��X���!�tom���.mMBq��!6	�&���Bd�ݬ��8����Tq�%���Yr����p�ˣ�%���K�|��6k`��n���L�Ʒ�GhH�]���l$���.}�bt�w���G	P�t��Wa��穊R�\���x�[/�;+��A�48�*�����$��De���6(��|�z��)�Tz
�0#6b(�0�w�g���|������p����/7%$x�� ��ÿ�1����<��9rǎ�9!s1q��[	�A ���������1Uq�k�,���Ŀ��3<�ٞ6�.Q�l2�|n�{��mcX\�b8�^T&K�\z�~E?�I�ι";�)Z,�x�ݠC�����b��ZF�[�AZ0�pU�Pyҳ yW�?�r�(�GWR��La��h���y��*b�r2�>t�!n����W�cVႯ'�6_�R,��?ǫ���<SW�Ox�T"�Y�X�z:��ɿ�� _ l~�s7�{&�m� B��|�;���<��z�W��~�9�kN�)�n�ON�N�������vB7�,�e�V����tq�ǻ.<�W�,�Dw����5%�������B��$�:�d�7��3$�&�졐SS��o�ͪ�.��Z��ͤ�Vm�̩�pV���	m!>wΝɚPCq.S;g�n����� �L���$��kf�E��>Z܀� t1>�BP�^=0�D=i�!ۈfKdT�q��-%����+���Wl*���tam�/04�q�u��<�_ܹ��,@3<N2�^�]��x�Ć�č����PG�b���ڼL��O�p�>�2�T���4Ւυ���~�41 �����"5���y]`�]����N>b*���L��\�i8�o��~��k($ޥ�5���Z���PT��������3d|��;K!vW�Z�7����8���,�L�]�0��PvOg ��	��������/���P��+"�&�'��\ȣ����50��R��#��"4RF:���չ��@t��V_H��sd^S��x�S1ޘx��C7��D#%��cj����隫m�ľ�)�[B�)%���T�v:H������HZʥ�W��6O~x��aOs�q�Eqp��A�|n�;λ��Lɳ��	��MI�� ���v����b4���1[E4L�
`�{*ũ��Nߴ,�~\`q]eMIEl�{8��Ԭ�\��?�P/(D{1��;+Ȑ=5C��Z�P�Tj����0���jN֠� !t�M�d��4c�DE���z�%�JIEW�~��a���w�Z�0TițO䔃�E��2z�� p9�k�����Ufa+5bM��xBR��.���@�W�LR������c�v}�īc�e��yTD&^�cc��.������\�Z�;�*��O�"?�6�i�UE��Cen���Lh�3:�:��l�yD
��t۩[�@�u���0�(`���y��VJs�̴�m'$n�$�&�6�G�f�� 3񥂰��~8�}oo�hj��\����㢠=e&c�JTڌ���]7�߲3-����m6[��I�/�,����v2 �G����_ռ��r,"�1S׶�6'��\W�2���w3a2G��P�@T��\j��c+�b'd�,�O���"����Z�W�R�t�𖇏���σ늲c�N�{l�����u w\�;��]��j�����[�b{�Bw���w���VF�aSpV}P_�%�{��A���7]��HRokG"�Xc��}ʋ��ԩv�g��=��I�uG�T�f�����;�W;��I~/vW��)zZ=����P2�W��`�7�����T鍘`�k�p+k�/���5�&U���4�m�W.��
��%� ����;o=!��� ��P�J������r���m�����,���z&��g���㖳A�#��E���מ�!DэF$��ar���:�	�häx��>������"O��Tϡ���wJ�W-KeA�-f��8\����*�=]�^�k���I���
��o�z�v.��������bz�Z`?kx���ħ����Lmݴ�����}�c��.��)�(\��IJ��;�P:4�]"l��и]���_�� ���I|���S�~:�H���]�Z7��4[d�Q�q���O7�8�.��2o��F"?��n��L��D	ѹr�:p<d�"��d�xS��:����Z4��y�_��`'���װ1P�c�Ź	x��}T~��CP������g�]%�92@��ߐ�����_�Y�OS���.em�Z�ϱ�b�q\b^�`Sb����Uj��RY$�?.�
q%T��e{j����7��'�Q&r��e~SEq�k
ذ����M��X�z�u ���7�"=�8�����r0��TM��=~�RT�c��.t���5:�
��"�i@)K��х}�D���v�e��$�Q�VoX�a�̧�X�)ӂ���X@V��V�Be�D~��F�n�
'h�/\�'�>uv�d"��2��|�iS3��"5�9�� |11����&Oh>냮u�����N���������тtSS(@C����P4wrJ1��j��hwڱ�"���p\U��7q�:?���$�����ԫ���Ғ��^�)ts�ڒ�v�맲�?+{�~,��C������c���$�������7V/@�!���1��@Ϳ(%�7&���3�tT2���@�ۺ%e��Z{�&��'\��aV�Z���������	��#�xw}Q�B��![)�"�<?���N�Oo�J��ee-��T����n,����[�O�o�
��[�#���&��q,�+��z�x���&Q�:9�5��(b5��,�bs<Ѝ�A�3��Y�l�߯_�	aܠN����x{h#����5��-�Lx	�I��ri�_�ุ]%n]U�GX����6�[�ۃc�o�/pa/'�!�Ks�9r񷘕T����g���\9J�� ��qfӞ���,t�X�ǡK1j�+u�ḓ���V��uQa����G
+�{(͞�Dx��_��������p9����F�dyռ{3�o��� ���Gu���w�/�������,yF��i���D��\,?kV��E�[�I���rT�SƲ���6\Q;�����|>��Ԍ�>o�r>��{8��8�
�K�I�LH���*�S�w����7~V^?W�s��ɸ5_�AM�wO6����,@�)�����)"|C��|GmQe��\���ėPl�}�,�u�Eju�e� ��\�����Y7ρ����_S���đ+�8��)-����J�;�V�^r��"ms���C��K',̰����9lM�Ub�Ǻ���<��*��yp?�ba�b���?���ǃ+D`u��b�#�^�'+�2��g���Zi��"�mGω��v�o���RBF�i�lڹ!C�G
Z��6��>͊|c����{=�U���Q�ɜT��-9�uIX�"�� ތpN����m��|��Z'�Dox2E��z&n�;�P:ؖ���^wE���l1�_���	�
�18R@R���Uɫ�.Q�>�/��{�M*��D�QD}�SQiM�,���^P@�J��������|�)�!	��D&��鐨������Ȉ�#��d��Pc�z�׈�`�{Bw3��Y�<���E�z��X�U��D.=�����	��7�	�&
-�=[��� �n��h0�uϣ�h�ISZ�B� �<��病�]ϋ/�Lp]k�k�C	��Z!��in�*��,c�6�����ҳ,-L����V6FH��i��ԅr#�H˝�{$ٗP���L��\�8�Y�%&���<�o����hi`b_~iX���bZ�#�@3�s;gN$���S dPU쳥�~X�+��d��OQdދ8$�#�����(~�"پ�l��`(l~bd-�jAa`f'�-.�N�5��;.=���S@����]5��rHN#i�|�NWh^�V����7ƛ��6�%�r�%,T8f���y_��B�g�n˪]8��i�Z�#�F[�.y0BuT�\���$%0�׳4�Wk��	�59_�#��u�o��}e���Ѣ�?Wؑ�}])]�!��B��mhV����A�]WR������m���u9a��a���^��͠��Ɨ	d<{f9|&�>�~k9���t�H��ȝ�/�x�oO>��&�E�&������1���5�8ٟ�=2,�OE6��Z��)�;9u�= QZ�IQO�:RQ��-c���{�C��7����\�ʵj,I)�-�{�_������+򥩦7m_+����r�*3�eN0Y��׶?��v������g�-T�4��9�����/�>��HŰ��E9�y�f�z�h���9��2v��� ���O��>�ިD:�,IfƧ�$�����@1[L�h���M`��>>H����T��?'�'[�M�i�"��ռ���l�1�2�Y�
\V������+�n��x+����)�o�B�-��z���bJu0�29����K<\���.X�X`�/���I��/h?i��&����h/cⰬ�b=���t��j�G�ŚX�G�O8QwGy若B3������Z2xz��]�������(c8tb�,���0���؝�=��@��Ȏ���	��Q~{�u����]N���]�F�h�Ct�D|!�yj��F�U����j�۷�9f0�hNNŚ�hj�ǋ[Q�և���M���/�m#EpR�6�1n�r_86G�:����? �qD�i6�8�����؞�;;�����F�o	9>��?E�}8bGX��j�/��4��pO�@�  |���įXg��7���&�N'��P����C>Oj����B���h��ь��o��W}[�%{g����F�i���P=iY�kg���'J�4F֨_7riՖ��WB�Q�@�th��yh8��{](S^����=6a=*���."e�������5���,H:W0ܽ��݌���[$�ТY����*�|�hyF�JP�uq7�Ts�)g��to4�HlT�7�;`����T�y�d�2E}2F���[�E:����1 ��{�ڎ��;:���A�3�ߖ� ӚE�l�iqչ�����󓠵vԿ��!�'�%� �4� Cw���((y����,� �����qO�MY��@&�~-�@0϶7�:	h)�/6y���8"�u�&�SL�iT ����xx����vgh�!H�������M��O4h�6�E�Y燨�׋!��'�,P�
%u8�B��t��%-�q�N�N�Ke���!2��;��+ 24��B��2�����P���5d�ʤa��~h!B+tm�)�iz!�	g� Q�B �l�'Q��-�[�o��	gh��v��њ��0�nf���誣1����N�F@Y�����!|^��b�,lR�5!���GV�"�~e�2��K?s�o{�ҳ�S�v�N�絆&f�Ξ��+6�;M��Zu���W��#T��=i�->����y���t�'�K��xaL�7fH�Z5&-�A��Lne���m����7����C[E ,�VEд6�c���67K1�+tl��?�`��-���N>	��$�8kk�!ל�����3&ѡ���g15b�60 �d4�)��8M���E>8�#�ރ�4�1��JtmKگN6?�A܀�9�����iZ�(�D;"��3DZ
�GkZ���q��{������J:��A����v*x��^��9�j>]�@�R��+�9��5�v6�V�΁��`��3a��51i>�$��/bn�5n���M��/���z����I�Rb�A<b��I߹�-�;<�ؿP?+p�d���k�X��:�x33����_�WV�_��|�e�~ۛǤ���څ(L�	���~�G|E��tx-��\��l�� ��w�#cIê ��6�!hOTr=4٠HY_6����oIE���hi�����C�����]��>���&I��:7�f��'�P�vi�py|��N�7e��#��/�,�S���`
P��?�C��FŅa�Y��PNb��ұ�1�,&��]�ڭF6�xut*#r�@$��f�6'ɵkO�����&���7Y�;�Y���ĩۊ�s��	K]l��|�-W�{Sҵ	��*9���ɚ��1A_˳�Kw���p�1�j�6��Z���N�;�O0�q��A婉uV��í-�� Er�|ײ�k��D+ٚ'7KD�&b?�
��x?��V�7H�L���������U����m�'��SO��%�Nh��h�[ė�'_��RS����t��o��)[���o|�`�m�g#r����r�i��]hKSJ��I�hZ��N���b�!p�ܵ-X�U�J�3��,UīF��́������;�%S����b��9��r�5�.��d������׀S9��	M���瘚[�nG����h���Cz���Z$��̖����E�>������
Qno"8 �v#��h	'��o���`s7�)6*s�>�.�R:�$3a�[����V�|K�ዞ���LGe��ÉDZ��}��Ô��3NCK�g��,���y�	�$'�	M&U�o&+���wꊟ��A������� ���/����X����+�v����98��dFd�*Vs��$�>r\�K�9EW^JH��vvk��R��A�w�"[�	7a�C���1�RIgi�v5ǎfD��(�OZ|�[���7�ONx�-���q�_ҝ�Uv�n�ߘ��H�j�\�x##T��9y���������*�/�`CJ~�q`��|���O���ĕ��
���|��|���8��߲Q5��s|2(�\R�5�~Iҡ}��Bt�B���W�k�zW� )��g;ʲ�<�
gz���rf��x3�a�/�h-�[��+���;��f^Z�D�~���F/�������?u�6��O�������!s�*1<ܯ`��&<�,�G�MZ,�����_,��;��￞���1��.%��$]�x�[p�Ӷ�!�_͊��~lť��&�"'���� ~5���4�/I�F��L~:1*�1nY��bn./��S �Y��Yb�T�y����:�a�Q⡊�q�W���=�Ui����� ]����B�p��)�y���ˎ���g���HAB�ܴ�Kz��J1��b�H2ʵ�M�(���/����l��clg�q�!�o�!�ζ�ˍi�����^Z1:���=��1�e������*���GSP:�������u��%��ҨUX~��`��\�]RKb����( �RH���W�yW ��E��Kƕ�0�ٲNp�{��ж��A���~ ���-Z�%is�o��[R��5��l5mt�C"?˟5Ey�����ݐ9��� `ʱ^�Z�l4z@r
}(ge��UO�4n����7�!���!T��&�h�36�����<*�l�b���,4�9����(���f��D["�lW���=9��|F=$������.��z�9�H��$���T�ƞ��5�"V��y���.Ҁ��V��*煤tB�HG��='区T���M��&� vTX#o❌�gN+���ړJ���t�F^�h��Jy�w|>ǌ��>��#(U;'�	�wg�C���9�{��u9�JQ�%��Ơr��0�_�������(��)��x���j^8Mk ��(��R*�Ix��M[�/�9� F?S��IG$RK߃��I �c|z�xn����&{d�o�ot��=YA����1D{=�b�t�*ͻ�,,k�Q$�-r�������a',�P�:���W��/�اcaLwЖ�i���t��?;H��5mx��B�/z���1�d��;�Mt���unB칎ӊ{�'B����t ���^�c 3m^{��Gf���"��)�AiA2D�g8HJ'����{��}�΄�]V^�=����N�2L�݌n���ԻҺ�y���i�%k!�Ѥx��b��.3��(�Xv� �|DF��pkOD���E���.�R~��a{��J��]�� X\xc����L���,Y���vO�j�xJ�Xl5�ð�_��xO�<D�%?H0�m���c���@�U��X�T4*����,�998�J�hN�>�p�����_o2V(��V�OM`F�~ �h=MrU �G�y�a]����k�0>B���a��1��[;�pB6I9�������������uh��b=��Aoz٭�l���V�'�ų��`�\s���-��N�q�nim���QF�W~��İj�#^��l��I;^�=����B�Q׆)�1I�@� �r�:Zˇk�"|�9�✼E�q�*)�s�EB(�C�ȱ�L̚��hN�
���M|z��g�$D�x�V��$���S�=˦b�%��;�6�	��?m��"ٜ��ǘ�.in�]�ٙ�,�p������Ɍ��`%��}Q]��ҥ3�/��ū���v�泘#(��,8����5��y�t�[����mA���"��_��?5��6��5ԯ+���OE�m��x��5&��JF1���,[�z?�}lR�J�غ}Q�����M[�1�1�j����<ʣ���<��LY��y.D���d]�}Y3>���?p��_cL�
(Z�Ρօb%�<�.�����;}�� �M�}��rͶ*���8�%I���K�P����\����~�8{����뻂ajb��W�����k�P�κz�	k~m��L
��h4X��b��~�H�=��vfI��U�_}��V��M����,K\�Ԡ�O�YR@��y;����EQ�[@��������a��������-�o��+]ӵd��H7}��`
�[S�-`/e���\iR<bnDs��I��,;���y]����U.1�����ep(
����6>a�Aֶ��3��ʟ�y[���o�t3�"�x{j��{M��c�Œ��;ƛ����*X���-]��e�z�t�U�Y'ҏ��i|D�P��0�x b�ߣ�[�fƇ�$"kG��N�a;;�X�#����TN��2���#K|�=Z$��K����.�������˪����)��j�Ovg? ���g.�H����7^jTbo�#�������g��^��t���ӇQ��|��R� ���,��C�� -���l|��&���ߗ�ޅ�Tߒ�ږ�6�a�gf���z���z'>�����A7{^�vrr����;�cLvN��Ѓ�/R�O����My�s=4�on{�c �:��(s7��I�/��H�t�6*�����Ǉ� �Ȗ��ѽ9�U�)�����i��7������G �x�"�*ک̝�f󮤛y�%�u���t3�V,5ߎ������X���N�Qz���e��n2���M^��/Z�z�:@X���u'8�R�tNg�[$��& �.(yNDӉ������'M�� ��o~� ;Æ�'2)��eayB�R��������01�H�^/��\NQ�N�X>�sz)Y����Zp�[�#_H2i��G�IR������*��@F+�kX�ob iRϚx$�]!ȇ/s��	Y���+��]ּT�ߍI���xv�w��h�r�a^��������� ��z����)j���^H(���`w$�;���#��<�s����7M������j���y��O�kf�j��00�<J� ���H�cF\��M���2�qʋҗ�K0"�P.�>����cY����M̈� �9�[8C�xj=I2���ΛIr<m�Oh��*�� ��\Kg�8T?����� /�V&�h.�#�VT�}hjřW�+ض�1�4q����;.�at���˱oNq>�2D;}���[�5�$��X��������&�ݴ�Z�$��\����xf�g=��k!��,�e�s#�ą���,i ���SZl~����~?��%n����r�� ��Y�u��j%�Pm���*��Ԧ��&�����ZҺ��5h@Y����Ca�*L_{}����s��be�}�����yv녧	����\���uyp�U}w+h�,�;��0H2��M-�}�O���k���·|���h�ߥ	�v�40�<q���yY%� ��6u[�E��]��m�@A%���UK�o8�Qk2�P$�'4���I�G�7��I�7����x:"���l��6�t9d�%[���-u��A�!����9F�u�bj�����`�����jg�!���O?~ơ~K��mR��R�2B��l���UF�����9���sx9�&8{�#_MB�S
@7ă�S��Z$8���/Jw�z��_���뛌�j��Y>xA8����7�!�M����	d��. ��U�IV~I3wf�>�1@a:7j��ĺ}�:�xU����&-je�s��šc1�F������Ԯ13J31���7HRz��zȬL�W�����#���C�UP���u`f~ġ�,�A7,�[+>vw�`w�i��D͘����;��[ʬ�/"Lw�V�>ӂ���
v��,�E�I����+(��&��`��e0�e�"�-�.A��;��-�ůҕBI\�,�)"H��� "�~hɬ���D���m��"�ho��>�z���-�Z�}�>���gF����M��P����,�_�°�$�\�Ŷ�O�D�֡Ɋ(�.����^|N�}u#?v ��2l��n����=@�Wc+Y~��LSK6�rӔ�TGj��[�4MI�mQ�Y�店A��=Tl�xE��bbD?8AYG�'wO33�W~ܿ�k��j]x4��Psyy} G�Ҟ�G�]c�ڲ'<	����pa���<6��W3LnU�$Y����-FǬ�g2v����$���1�:��8	T���а�,[v���XK���-;ʟ���G��^��H�������A�/��1%Cȑ KN-����b
�m/����Δ��eͨ8�&�C��:D�L!+U~2lt��?���o���P��r�l|���tț��T�-t�2���"$�S�P@����e��t���Y �x��ZƦ��B��6E|�kf6�<僸��QX����n����آ�όv��U�7l7E`���~��-?�'�ʸ��u`]bmK����𴯷�lW�a�]0V�]�<{yO��(� �_xtb���!�+�+8��XӰV��A�x_G�9K^��F�����.��-�B>�4�� ��e�vi��fSgA�=��������~��3�0���[�#��@̀{�2�iw�0�Eݿ� Qж�s{�D��|�8�(�F"�N	���/���?���/\��Xۺ�� �+�*�����l?��$B��OiӅ�Ƽ�X�ԁy�Y��.lQ�Kg�N�Pj��Y#�W�ʼ���f?CKԯ��gX��lʆ(��B��<�iR�ԙ�S����C��������ݱHv r!_�5�
�ڬ�����r��֫��zp3*L����߾q���"�3��7�K�d�Ӥ��3~�dc�H0�{�i+�
�}5~����#Y/l"��m�`.�JFư�.���,ծ�%6�:���}A�c�!�Ք�n����9�.�5^I#ZHB���¶������ x>U�*�`�($3'<��PR���B �}���~	����^����{��&�)�)���6�@��M�{�xK���/�ʘm�]g�*LDe�?v��q��֠5�(�w���c�����i%s{+d[>����Ҋ�!~)E�袛 �a�V�����N;�(߭�KJ/A�r���k)���?�H�-+�Y`|�\��:�ܬ{:�F6��~U���+���	��W�}�~9m��,u4e��L[[P�,�_^j���e�L�����4��r�P-C��v���'1� 6Zj�D{L}Δ_�uxC�J�Og(Z��W:����v�]���*>^�+\�¨`j!v'��X�#gy�ٌJ3�I�qa��D���2�PW	�;5Ʃ��x�?0V�nQ��;9�+�6�nN_B�3Ґ�'MČ�ʜ~\�Ww'�猴�n�����E9�L2	�Z�-Q�}�;�$���\j'@�k �k�Di�Ũ@5���+!f"�f���L)0�PA�f$(a]etQ.��h+$�7YG*�z�<���@xk N��w����G�(C fl���Z�y�&������8n����$�뙑�	���Ϡ�dt`��x��(.��KT���8�w�^��K���thDXWk4�M�� �)h +�p��錐E���Ȋ��&c�:7��su��M--�H�po�fa�2����m�L�<�����X�U��) ��ѓ?�w�!�����gie�	��"�e��?����Sl�]�f��"��Ne�8�*����<J�Li�w�%���O!0f�6^/sSK(�-�)|%5	�,q���B��m�a.zm�Z��P浲g����g6��(�q��������B��1{l�hc�u�p�����݋uH'�N~UC'-�f7Z��XӤ�\��y"32G�k��V&d��� ��b��J�[�@4�r�����aZa�L��"�"���T���W�Y�p��N+���g�?vC:��]�ඪ��I��A˩ȳ"�1H~Kx�6'u���ݗ�G��!7��a��3rgf��{ܡ�?�~�1^�C�D�)����D�>a��MX�}�䷩,���Th�3����Ye���H��V���S/�:i9�T�*/�;���id�[��)�~�>玞�Vў^*��j���q���I=�!�4�(}N�(��D\��vO@���C ��]\�-,�@�N��cz�(F�+�Un����}B��Y]�D^�UJ��x�ުP��  h��i:=�Bߍҵ���ch/�A���zh��F:�=�o��(1�$� %�Y��qd��&w�+=C]7'g��Y�͛˻���I1ɳ�ë�Xn��''�N8��3i���e%F,��I�B�p�b��Z��.�C����ͦ�:uan0i��S���c���M�]Xm���(��m���p4(	"�#,3*Qk	�P;��f�=1�T1��!c'[�og���|}��h3�/��h�-�����(7��eTG�����8��?�F�����+��5_}/!'��`�����:�n��2=�E�B�=Z #B�A��+2g(Ic/F��;e6U7�
%�����|S��yg�6ūy��t��R1�/�N3=�+-$1��W����ѱ�n��?�75��g3rA(�����	;��%�P6r#�?F�$vP�u'�w:�!��Ig���K�\"`/�<}93K-�/鞬�l�����$Q�oʵ���w1;��+=�##٬���������q���?��p�k�i�����a���d���.l�9�32<�䤓�&�: z���HV㭻�����Up��橖|v���~��m���l~�?'����Dxuf�T�w�9XF���o��:�r���s�_�N�`!�{�V8���@���Lq��q�]"���7��y�k���A����k�uN�^�$
"�	���0�����i���� =��t��~��2��X��W�5J $��l%������c�p�)xE��HHu���v����l����Qa�G��Ge1����R�_�d�{-��6��]TdA�dRĎ���|��ĵ�qcJ'���v��ȧM_ro�)-:Qr&T��KN�Dȷ).#���F�� 4��֊�-jO�N���=�}Y���,��*S�C �BZ��l~)3��/�v�M����\wX�t�ZFK+���z\���!�J*�����|R��G֞5CKAt�t�5��+�b�'[\�-A���d@b��x(Ԕ{���cH��Ԭ�:݋�$b�Wܒ����/W�9�"����fV?�V��K�lVG'3I��35^��8�MR����Z�5��ʍ��~�ߌ:vk,ċ��h�6�=J�N? =�I�p��<B2�vb�jJ�<�Ϫ���OVQ����c]%mM�gw)ʂ���$���/�R
^�|O�o�i���$�_�~>�/��_N�1bp	��Χ1̙}�P4_o�ԫ��!䊜-�|5���r�;�e��m3ь犗ՏnA����;��X��+�\��HQ�$�ӱ̉����O�'p�D������(%)��&��xF~n�<E^mnt�Q��`����r�x�x�D�	���$Z{ƄԔ�4%��8aǠ8ns�ej3n	 ��f)�'m�����F���Ѐfs�+l]���c�R7�t�Z�';`�.���~�^���IXͷ1���]Ω/1�m�] ��8���!z'~-�Q�#���RR�������}!�������zJ���I� �3M�Pp�@K)��Ħ��G�N[��襵r�����l,����a#��{�����X�����ro�	�K�����-�u�������Գ:GpM����流1�6>�����_�A���rIT 7I�`�鉶esf
���xn%�� 2G�K9�,^�#�����"����T�C�V3t!���8*��V���z,AQ�V��.?[���4~���[�WnS��qTx�O���H�My���Q?�$+��\�����vQ�p�D�~�?����G[�&����L���Ǜ���&�틯�{b^��K$7e,��-��R�7Yx~���ئ	4����f[e�9	��9�b�<��\e� a�&E�X���7�E��������B [%���PL�+;��i���PX�}�1�w42w�&�[��k�zXGqG�.0���k=W2Δ:T��\�����骍�K���ء7��Pk`ij�2��pБ���&3���E4�����7_���q`$<}JbK�u6���Ɣ~X��TG��
�
�hںW�t����<�'��c֡�wT(��ѕ�ZIR���dSy�Z�^����f�3)�H7�K���f��V�,삥�����y2R�١�~XgY��X}�t���*h�:��ބY#������+�ݧ��26����@sy�w��:o��Q���N�����.���E9�����lk�*����0��W.KO[ ���{ќcaJ^�@O���J�����D�#�^�l����ԝ_7�'��O�]����D���j����qjd���{�;XS��f�aF��Bqy&��I߈),�U[��6��enD���/T�����6�(-�27�&�g��$��\�f�S��x�	��1I��:�_ �1Ku�p���MwD�\	A��n@�%�H�	�FH��@���-����M�He���W~�� ��<3;�eA_��m� ��9@2��� :�)n��'}A{�DRdHY�V9�?K(�(�m��{q��XX�(��f���g���"W��":�5��`_���;���S��s|�0_�c
����L0e�/�-M�Hm�7�Pj��4���<�~�Aىt�!<�1��$BW�ή>�=��2\�3x��O���*��3ȪW��$�|��ɹ?�ڪ���v�͵�'/�, [�	���i��<~�f����$���VRS��T/��~G�R�_�5W|^b�-�Ej�+^�	�>�8�}$?��t��֣/0��|��y��-7+� ����U��
��wGG�Y�����i�*#�&Ω���_q�~�� �����5��}�M�b���֔Mh+4�;*��ϓ�����@!��L��%��f՝��U@�_'"�t̆3>��L/?v�)yS�QFn�!��ODXx�����M�D(��9	��M]��o��r�lV�oa����kq�t������d���|HZ��0��V�����`#�?�J�ʶp���Ĺ�ԉF����-J���+a����b���u�v��jͿB����\/f�۵XZR�a���?h�atm��p%q�G�E23��ZB�&����Kɩ./�\�C�e,���G�h|ꮸ��a8��1�H:D���1���续���v{/
�BY�`zl2���e�!	A�͸慰/g�!0.��>�J�V۽��_��?�Q�:-���IW�As(�;m���ٍ-�@�/���%Z�+䫝��{�"(3>]�6;M�Ʊmˤ�^��Мdz���x<���ޖ�\d5�hI��su%=�~U���N<o��xXc��T{��'d2=n<�	�(��$��!醊+M��=P�{��R�w�.���E��?¼�8��Yz����i����Īc���&��>�l��L9�v� ֹ���Uu3/=t)�S�����e�g,C���L�-B�����4�aXc;��@��@� ��QMǔ�+�A6��Z{G��j`|�v@��K�A�w����#����3�Q��������3l3,E`��Z�(T�˴|��vM����X4�}g��W?U��O��x�uA�S�S	S��B�8�k����G:����|��G�^�/�3�v��.�5�;a��~d)��%�A6������$h鼜[F룾Q��6�?F�2�_Q���PC�:�y�������KT�C�5x�W���3m���4r:�v����)Iز�
�����R�o��[�\��pS؅ys�;�F���<U
S܀y<���e�FWQQh��
k3Q���F<Nj�o�\b]�'��㲑A3�;��/:u�=q�*0_��Ĺ�/}��}��ߪpw��'x�H��͉E� ��2O�P7�=]����(v����^F]P��9�I�n��v���J=h��RQ��,����^��5]<��	M��}�QW��#N��x�[�S~���U�*��,5�#�{��#�IBa�cGeAϢ�P� ��w5ַS�=}7�|��-׿�!�v�G����F�MNb+r�ȵE�|�b�E��o��(��jaSq��P|��iV��^H�g�đ�+�D��zNh_	g��-B�ү<9l �G̦O[v���MX�!Y=��z3rpm��hR���{(-/84c
���aW����y�p���͊���^O:�g�iW����z��%�#?��:�6܀���;;b~�-��N�g��Ż�ks���+됽~�2l���Y�d���_�$�}�D��p����!���*g �N	l�S{|ʚ�D�Yc7!��8 1�p�>����z�v��_�E����j���)c!�d�+�	�㝷q�0<��	���N��<ޏm�B�zL~w�ogǊUߩ7x ���!�?�7H�Dz�^Α�R@��1j��RMn(M\'�wvؓK�`ԗ8�F�V��rp���-3>\��[	���/%I���~�SN&��(<4~),Qs+��W��/���/���$ڸ��<�%^xE�%��$�XX����t�/N��S��䳷��BgW����9
QN�]j����K�ٸ�޽M�:�:w�yw�������]2�MG�����W��^HtlS�O��N<��BG��?9�AA:����0翺��^ˊLo�j�@��A��t����:͙Y^H�@���dP~��Oxp����5���C�����QI�N�]�r�4�VP�X�mb$]&z������v���xÒ,�X�Z`���>?Q��)�C7(�Fz�������e��._�����~���f���фob�dv�tcL��x8��3Ͷ�R?JR�l�D\�|;��Jy����ҏq������?A+j�\-�dǰ�E7�3?�+�����9	MS�ש<�J q݊���R��Q�B�ɋ
S�����.��=��|cY�m-��.6�� *� ����;�lk�¬��̺튤L~
����M���w,q��Om�ָ:�S!e" eT}��*���^$�3qx���M��k'd�n�HҴ7��teG�6���J��}���=`����F����(�x��2j��.կ�w����6�i���h�O#�Bf� hd-����q"�GK������tI4��]�Iɯ`��L�a1��}xV�6���Km=p�.w��G�LS<���y1<�j�Z� �w7��	f�J�F�è=��h-�f(�(7k�mW@9Z�	S����n6��~�y}�wO�9�I�%O(T� �`���"�ʞ��8����;F���%R����I�M;<B�iCɾ����;�&I�bE�Oݍ��T\ �;�D�a����6$�-��pM	HM�x ����7"9�H��s��Q�ef"�EHR�-x��A���ko��M#u���G�G"
�g���qR M%�*�&�O���#k�\k�u1��U��׍v�gU���ZL+��\6���B�P�֖�.�f��y�-S��>4�?4��6 ��C���wfN��{� ���^8�% d"�L��&̅r[���|�R�$��C���]�#��$L�4]���d�y!��ʨ���:'s���9�9�y�0�m�p��a��_z�a���R��[.BX)]�=�g�Y�r���>q:��'�AN������Z��.������R}z�4�ҍ-��7��{��rjN���N�L���55���HL���%u��-���I�!�h7Oh Y�&b���1���Oy,XY���sGb��>Y���/��S����Q�@���"��r� �g%�Ѳ�3�T�i����	���H<�;�*�t��0��^�B�P����U�=��W��f��ޛvm�/�m�������4+�E�q������xIyĝXϗ�U�E��{�=�
��D��&�w}��q���������.#�)S���!��v# %��BQ�̺��������`n�)�d.�l+�&�K��MV�t6C};%PUH�ء��5�%l&Q4�8�e8ڏ�uGp%/g�Z�������n�Ǣ�u�gS�cLӠ�$�5��z9p���k��,�ir��Nw��8�yIw'���ڛP�	�~�%n"31:a�!wb�V�Vxq�BJ(���ԍ��m��KC�wB�7��ۻ�y�[y�*��]���� Ў�G]w
g�Q���61CC�1s���Z>wKN�d�Կ��}���s��!:�T�ߖ�r&�/��u��V����.��z�w�g+Ⱥ��,�??L��$+t���7w�%M��v��4r�zuu�j�K?n��~[�E�Oer�����cnd�p����\T�����vpް��Y�S�x6�?��x�;��X�����By��t���ѕ��ӴGϪ.�*-�����R�)r��f��=ԀK�Պ�3P�N�����,��"�/�6�rW������7��5��;��2�$�>%7Wc�s�Y�e  JX��B�G�h��zNG�(�,"Ⱦ3'e���@�������������[u�b��O�!��-6���[F�g�h�$�2�,[���9�Q;�`��L���c�s���6�^6h�w�u�Á.�l�E`�- ���s�]R��J�4�}F����oh���x�nQ,g����N��a{�e)�o����뛰M�ӟ��1��G��d�(��7���"�y�/�Di��]�Jk��h,��t���-a��`��u�_H��߮����.�+�~��X�t㊤�����r�J�+���H�b��e3��9ϏB>���#��k��NiG�u(NcSSj��B⠄����ds��S�r���-��
�S��q+(�7����l���@�y�i#&BHN�8�8�<ݞ���U���h���:7��PswݚN����E�����	5�v=��mqBx��M:�6x@ծi�Ft*����`8��;�h�E 9s|l�Z�({'vL�!��Sx�2�
(t����}���O�\�)���V_��=�']�dy3�����
f��i��tc����(ܗ��������B�Yܹ׭ڊ#�
��R]Eo�[N�e�Y݄�+��ʇ+�V��2�??���>��*2�p��!r9_I�>�^q=�2����}��b��
���ìn񼮛D��1�����eڻ��"A��"��D�w��l�;��Vs@�̠�#�žQ��Ko�&CC杋�zt�RE�������>� ��D6��ѐS�j��+*�C,w������?�]2_u0�=��T�Ҫl+n��A���c'��b��F�Ej�8����3��@Aٷ��Vx�c(Y	O�;�1\�"Z!O��:b���� �,�������a� ���6CO�vR*��N����;>�h{�Q`�&_S�^�YНL�2�^ Z�k9�s��a&naA]��}Ka�u�0��w`�V,t�w����PW�^�feX���[��ep��7�P'�+|�6�Qע����¼=��n�^�!�F]���^ZG����t��@�)fQvu��s�HF[p `v�k"3\��Rq�0ɀ!�O�8��8�룑���v��s�_'a6��h�X�W����X?(���A�\�P�٥�ES�ſE��-�Ê�N��C]8�4�qpIj�3�&T�6����*���Vi�J��&�k��*��&w���?�Xm@�C/n�ޟ�aM��dX�^��<$.pE��g�;��I���$J�l�h�M�$e�	K�(�-:�; �!���.U����V����?+�J�;H�=�����D���`P��xVZ�zg�h��}z��su�g�q�Jv�����? �Ӧ�AV��Y��!���Dc؃1
����D"i�`�[���
�z�����D.Wh�f����<>3�Z��{��?o��<�'��=��˟�y�QF�� w��ͯ��Bƀ�@�75����1�c8T?����DBu�1�����2P��;頴�G,:�f�S�jH��ͦF�Z r�o��9�5i��<���A�	�5@��^4�i��~&�*�)�ck,㾝��R6�t�ɝ7kqY���E
zhP�u3НСDȁpiP�LCQ�
w%{�z���1��oB���r)/>{~%u9�2	�t���8P`Tc�ќ�2�r@�;��G�1@�J�Q�Y!�ک�pw�H'@(�8Sڢxr�/�}��M���Ex���{=	M�z ��>��8��^�QG�Y���!p��̷�]z�1�(�lʱ�_�ֱ�A�ቨUНW��q/��x;:��LM9�����6؈$�2-���R��$��k���K����~�S/M!��&�_ k��}D�8��PJЧ����8�3[*<� rl\�#�I�Kޱ���pƑ�������tk� �X����9�3�}��l�C��'n��&�����[�EaC��� �Y���2�)��!������H.��������sp�H+w����C*̏�cIH�X:� ]˧�HB�aI��މJU��]�ͫ����ʊM��ԛ"�Jk�O1����n͒�Ur��W�{nbnm�ĸ/-����d�V���(4O;���M�ْ0����do �_����7���3$]��~��FArB��j����'ĵ1&C
"rY��j����
s�QL�h�WS��$&�ZBx�q�$ʩ��c��%i?MKC�sF`B��:`"�\��z�g�$.�.��*��}!�����/�{[T��2�I�˟�X��ʍ�+�S���y0$��G攭�+�IL�ou�m���M�ț$�D�}�:�ں���75S�
m��������d����zv"�'x�~>�tp�U�ފ�zap-�GQ���lYf�]���1}�a�J�'zUg�JҬq���-����r��.���c(���)>�ZR�#�,x�2�y����V%��l!\�D��xhU��E�.��:��dg�ƒ��ǝ�W?��ɘ"��rMW�V�5"��D�-=��lS���� t�8��U�n}i\��(�V�_ta]c��ZF9I��#�ԟ���#cԴԐC�n�,n�� �,�w����|�|�k�b��O��d;Ak��ͅ-e����퇬iGDS�Cޮ��^��"p�mc��K�P��\`��;�[�	����2��B{��b�̀�,0��JL�bcB��]��I��d�$�2�#8>e�h�%���:�ˠq�p��b�y����X.WI�%�� *�Y�;����Iw�da�a`S&eiq�>p��E�y@E����U��}�	!�W-9aZx%��#�EO���B(]4�S|&I��h(szy�&H��@P4���yd�]��屭�V������@��]uɋ�m�����I7/���`��A��b��7���3jв�)3��JUdL����^��d����Q&&͵��0��\�b�J+�bp��Bӓ0����H��z���\�J� ���}y��6�.z-�	�,���9�C�*$�U���ߥ�4e38�h*j��:uԸA_׬�S���*�]�[��,8��!�w�U_@	L5@vY!��f9J��ߧ���(�o��R�u�/eNh�I�%��;���V������CT ���O��Qt�ɚ(QZH��f ����T�&u/Y�g�Z��A�p܀�����f$��QZ#�k� �Zq�KT\��bM�l�k�j��g�Oϸ/�"��C [B�i�o��%M�?Xn%)�+ÕfT�:�\���~�:R6n�qY�r�����Dn�k��D���Buv���U\{<:��֟V(�c�.'������������Y��ر�N��a�1_���zcE�0[�-����b�t�tb)��ArS�B#���]�`�cG�X���TH��,�W��f#w�͚΋��D/v��G��Ai�[KMH�1�K�/BH�\_����U�F8����#�k]4��[$��ɘ�T���fш2c���74����Oq)j��c�#>#��6Gh�D&�{���_� ������ǰ��7j	>u�o���]o�cά7	ԡqߡ;�
��'�b�;��+R��k�xoQ�B(���u�JH�e��iS��2�x��
��>��W
�A*�`�N0Sъn�r§_Oa��N��a�T���//��j����/v������®�L怸�6�N��;�,O��Z�|0����Iy������eR�wf���۸ +Љ	�~���uj�#�������u��l@��&�Ki_MY�T����
���p��Weɉ�Ux��616����!D�K�8�W�*۫R ���Z����#Pػ��$N���  �6Y��J��,P�$'/h�R$3��@��Rl���#�L��#`��3�?:ӐP�#�4���{�eA�o�?�_�Уe�����?�����Aj��P��$����y�sn�'C��E/�!��X߾I@_�'�pЍ8O���&�8����*�� %�0����ԓ"��ţ��#^
��撽�6}nc�z�DmwF��^7)�v�l���d������nK���Rb�ՃI��Gs�c5����3�+���*���x�'���O��
D�q�I?�1�m?޵�w��Q�j�S2���=H(�~��֕�w�(��)�)x�����|�����x3�,�G>�% �(��QCmP�{ � �ͯ��GN6ۧ�˓΃�{)��؎��G���4O�g{~rs;Mi�hY}^��t��<T&#�������>�7u,]���NZuY>@��VJKы��?��C
�V[�`�d��0���}�k�ifte�GM��_H^� U.�E����Ⱥ]�{�E"JT���t��G�r�[ض��c��X��P"���hV9�/�7 e���P���?� 9��yHkme�����R�k{0�1q#qh�/���b|�S)��L{U����V�۵�kU~���BS���N6h_�����ߠ�z�ֈ�<�=�s�n�6R�UY���J�-J�jgD=`�X��A��=�~������m��a�D�M���3�Z��8�G��mO���L�����/�'�=�!�c1gc\�Ybζ�Ԑ�r|�*����&"�5ݟ�g�r�v���	_��;�e'U�m�����s<��Ҩj|�3$4X}��mķ)�v�q���Q����S��u����r*��;r�� 3Ş�Z��<%�h�Ĝ�ބ �:5�j�%.˦PX�ED74r������椎�o_�Ů������=]�C��"꾄<WC!�6"����\�MQ�w/��_+q�nw�z�oe0X����U;g�p�1��T��1�:�4������Jru�=����]��7���~�J=���ۚ��z���l��d�jc����F"<V��C3��~i��Z�w�'B>�_t�Q��U�6����������@��IW�����F�^��-��l��d��|G�1�HH|�_0wT����T��s���Hyh3��۱���"�>St�"�Z����-��CP�XF<��G�|�9U[=�� ��Pc0��k�B�
!��$�7�`9�f� �]=b��Y���E�"p|�N�Ҫ���a�!�9����-a����z�9��˶��T�� �Ѕj�t�Q�c��G�Q�O��ep��l�>ys�މ��6�n]H�؀�̧��{ŕa���.��O����`E{[=�xg�w�<%����+�:Q�2v
0��^��#��=�c�UYʂ�e�f/A�mr�5:�	��*	�~R�v �.x�. ��2�ǡY���݁��pԜcC�)�!E���+�P��>�
���'i�Ӏ���+r��qzB�Km�Br��w/t�[a^?��SD]Z� �H������g�t����B*��SU�h�k(���<m,�$O�:+�	��?S%P��ԋ-p����*:=��H�x� � �ʡ�.�c�`;%���(����5=����T8�u���s��E����d_�u����]����(66Ƶ��M��ѹ�K��~&�`���.X<r �,��nX���`0�|��r&�3p�s�	[���	 n�����r�K���όڲ�Nh����g��̖��|�!����-��T���2�c����1��zS	R�b���J�|���׳+�D1�����Oe�����Z�7n��"ߎ&U���hܮ��k*ڦ��xVD��>E�A�ӫ�9���ō�P���!��юؾV��Z
��+M��c�w^1���KT��K d�$0�P�s��\�k������a]s��ZD���Ϣ:�O�6p���G
VDO;D���H���BU�0��3� �[(�K�g��;���f��Wo����v�[?m檩�9�'g��]s�#�/F�t�&�ZV8��3]<G�����J�/k��JC�V%Rq��|��m�=ٯ��(�+�<�m��WЉـ����|�p����Oj��n�0c��zޤ�މ[�Ք�S�e�7�%��0�4�.�n�F&-91��"9��_��Kw����P|��T2����B�W��z���w��C���Z���eH���ʔH_�I�*�0U��3�wC����J���В4���y�������U�hN{�E�����jᤜt����[Lβ���@�}����G�ѡiƃ�Ȭ���_��*�tdf��*�R���?��u:�٩ �����CV��+m��[���Dd�~ ����3v�ۣ\B��5���*��mΠ��}���}�:S$����1Ĉ�hg�ߤ��t��V�ً��� ���^I�=K��q�i�āua<A ��f��fC��q��g1Ùqy�XcI��kfӬgΟ4f�����o~7�;XB
2�}F���n��TJ�f5�mUȚ�E,�0.��YIf"?C� ����y�b�>H=���P�X�]u�^8ϒ�ï�cf)��r�s����0�_n%�7�V�F*3��O#�z���b��3'yS"C����"��Rv�z��h��^���#�s�
����{�Xh�Ԝ	�	�=9U�w<���g�����b�]IN��r�.I�-7�g`ʂN�௩�ˠ�����Q��Ȍ9���%�����[,X�BXEуfzX���	<�1���~�Z�\�A��5DR��|�\nW�L�J����3Un%�!E��i��2Cmϡ���y������������	��TpN�y�QP`]����뜃�#��\���i��J��'�~�؇�TK@DB���fI�c�U,Պ��l� xҚ����d��YOP��;����*c�&�9�k�2JD��YfVL
~���7����#����W%o��QEL� �D�]�Q G�1���� $�+�R��+�kK�COCO�|��Ǽ"��/��z�0�!Z!+��G'��L���T�xz���<���O#[����������JJ)a� m<�,�����B�`y\� �pA4�/�{T���$����qn�-������M�; `�\-~5ޘVܢ���#"�%*�f'��
�%���?�Ϫ����j��j��*��՟�z�8�<���5��lh=(�rqع�>f)�K��\��<Ly��Z c�C&J�W`�o/�1V?�b�O�h��xY�0� ��@S�5-��
���oҗ��]CSX���+������_�?�·�bq�"̧�v��?���-��?����~�{���oڿ��w�m���d������ Q��z�߃�%��=�=�I�pgu&�(�vVW���T�@��^���PyEu�#� Y~P����'��E�
�`���r����6��I��KE8�����qp�n���+���x�A��D�ң�!�o8j�B������'V6̆�<���Oe�ƅC���?�K���_i�&b�&����B�r����R`��W &�G�錀�����-iX��3�2�8��� e��˴d��llq��TUƜսc7����O�O�%#i��q��+p�߇��c�#����ƥ���_9e��K����,<v�V����.>��l�랰$_�eF����Nu}�5k�y���E"���9��G;�6l���W��k���@�m7krlU��C���Ҕ����������6�R�q} <K��Z��efz��}a�fTK
�c�vXW��ν,$7%�Z�$ݲ�2� [�t�130�;z��t�H��ӵ� rv��ð=^}G��^U�`�Qu� ��E��p���ˮ�h����#�Ȼ�pŋ����9�iͿ9R�����d�9=�c7�g�$�M��1n��qC{��1*�v�r�E���=s���%�䰰������t�'\��ɀ�L��г�����<-�H�o�5i���o�`�9���I¯�z�`�iəUh�0�
?�����E+Τe�U3
�&�]��)G��*O�#&���ݕ��@ju/�S{�H�����@ATS���zG�M�N�l��s�������r����7�S��Q���S�Rv[nU?��~mV�Nv��'�����Tm`��ic�*�Xr�n%l��w����@[\G����ACY�{��Z�/����Cf=.ďT2�j�̐O��� ���3�?ƨ��I"��+X�lڎBZ��bVoϤ�i����d9Y���^l:n�����Ng��Ka�����)��{����}_��e�������~����$�w��.#wӘ:��=f(of�guJ��@8�����(�@@	��)D L9���U���`)������!���	�G�މ ���/�2w�jqīl;����v�ܐ���L|�v��0k��J��y	��vA���H�����op8���Yύ�kwl��WmЃ��������׶�ɩC�Ɏ�6@-��][ �=X<o�ÑI1������ʘ�r���(3na���6�8[Q�G�r?�g�d5h�q�@ʒht�F�rq�۠a������U�ۊ �d\~��F���Ω4��oL�'B�����쐚`[�a�b�ĺt�s�2�앂�ä�C�JŚ�ۓ�#��B��Zw�Rg�LE��`5p,b���c������J�����@�Y1�[�S.�����|�)��lȀ�m��)Er���T��@�r��)yjoK�۳��7�%���$n̓�5�'z���v�y(��-�N�1y�O�mC�gp-8ds\~]YE����.��`�x���ݵ�ВZ}6�b ����AV>��~��՚ٙɤ���/�*���KQk��ԃ�P�;�ww���]�A�_�~�	"�x&��|�Q��^�d^��\0��s�d*d�˱x��T;��%���iw�ұ �J�˄�Õ�0Hl���=Im��W���2�aM��c���%���I�N��_J�sC�@�S)�k��-	�����/<ͷC�4�'��A��Is�6qہA������Yi	MY쨐Sl+��W�>u|�-�,Q�'<Dw/�d����WtB���{Y"?fy|�ܵY'R D��	�k��-s�q�_�摟ui�L��1���k�!��o��"_�cG�2��]��ar���(����+[-�⠅��1K���h>覌'	nD������4ni�:�+�����1I�������AGk�G��؇=I�	ވ1��� =Yh�^noRƄ+�P`ֆc�;����!㬍�!̇	��z�6��������6��_����13{�z� p_�dV��%�T�I.��ӊJ�u3�п��]t-7Pt�WZI�F��w����k��t���"ϻ��q�)�\ը�k��4�m���/`��5z��z� %��+��3U|�e�X`�������,wg:uM��K�xf�����n�7����Bi#��Q7�("5�R<�N������QTOSQ�nw�a���� ��%7�Y>]Y�����?��	�3�[<�� <��{��|���]�zA�t���;v
Q��s��������	q8�!�~u��M���@N��ܚ(����e0��g��.���X�f�G_I.����O�&!��:>nOz��>�a���T��G��<b9~�xJcS6;\Sug~RA�!)��)��X�G��x�(V����9.՜Xx?AR�@�n�۸M9�����E���������j����C��Ξ�=:+�{g��7i�۲�D������&���J�h��<�ߖ�3�/��c�Bj��ZW��+tg
�|�)T���0�J��:�8�6�W���݅`<����<t^�Dp�`+�\h������,����վ����.��7��*�����J���8P�b��Ÿ+��R�C�M�	;��`a�H�h��n�dH�{��_̷���n����dx 8���Y�9u����>9���k�4��R.�X1�T���w�w������`S�F�2h���~��|!aZ5�L};�+�cM�4pka½��~��:�,'
��8���v��Um!�@+��R���aΕ��C(B��-���?����I���Mv)�ݯE3����9�涿���6��f�|0EG��*A���x$i�I�zMQ��������:��Q��ϟ(,z���z��.r��R��H�v�q@0 �A�ʌ��NQ@�� �Y$?����^�9�l�Ly�șk)�>8��T,��yv`�H?>��Hx��k�ĩe��[�5��:d{=-�C�a�UZ�~Ю�H_5�B�x���!ww�#~����U�Y��9�ݟWS��@[J"'��~#�?�Q��ʋdtM�w��s l�V��cY6Hɗ�jgbgqX[���#��7��0�<Z2P��l, T��ig�B�()G���C& rD�㟅.� ��ܖ�&�{�ͩ�r4�I$�5욹�fcw�2�e�x�Q'�P,�r)��Z浰�)����|�m#_�V�2m�֫��g��47��G�\�^����Ɵ��6�(��/`�s�Q���]D/֭��{��f�$��-����s��
��`[;���/���������z�+��@�_�B�U�N���n[cI�ZBe�g�Ӝ���Y�0�O����� ��Ѵ�����; fJ���&��v�s�fP?�oɉU�� ��6%(r�U��A�@<�؍A�f��ä���PHu��$�dc/?g<�)7g/��
���B�}>ܴ)h=@f!�(=�3�����d���>��(�L��e�{U�O������)��K��be�aL��4;�x�+0�ɸ�&~���SwU[֧p�8c+7|�x>7G^n�>r߬�*�h-�P��w"�c�-�]��
�{��R�+3�5�a�.5G�oK��e� Q׀[�X���3��_��~B4��?�I���!�N?|%�b�똪��M���u6E�฽���<��Vb��k�n'"�z�Z�NK���Fi=��-�WD��6s\���Y&��ʤ��	~?	Sc9�V���o��m��d8�^�s�hFT�;x�
g!����TL�(��.Q^,��d�^l �$/s�����F��]��?F���Ћ'�O�̡�޿�?.~"���71�!Ri��25M�Qbx�~�?z�ĭ�'�O������</��%z :��
C/��>NvC/.���P_\c���:��k2���͓��-Y�z��AW�D�����G6�E��Vc�M����̏>�$��R�ے=��h9��:��̒�*�d �Ri����Ap��[�Y`�'JI���-.�1,xh�Z_9��>}�؜0�Ev�*�c�W!kt�9��.U	3*4Dߥ�'�c��f��(Ļ��z��ya0�z�����]�����֡/���V�Jd#`(��zv��Ɋ���ݱ�eũ^ښ9*�Hz0�����o9ۭ'�H�T��C��(��j��V5��i�;���k7���m���������u��񕊷�$\��r9�")�z���q^�Չ�(cRT��ݛ��V�1>��z{d@��?�"��%H*+H�/0QHS��5��>
Kil���ޥ6X��LC0�����U�==����Q��]�b��*_�L�Ҧ�*D��~VX�εzIb ������ϒ笘��ϸ|dY؏Zݠ4	�>?�ZS���YLO@?��f8>*~0^o����^ﾯ���?1p���g�9N\��L)�h|�.�v�6��e�6X�y]����IcО�9����
�l��l[ǩ���R�YO��O�U4���E����6�*5����v%���/��"m���i��R�Y��)�Ր��-U��5�ɏlg6xVQ�p�J�Ժ�IC��h�9�B=�E���w�;~�-��D��7�p��~��.c�@61m~��p�I��n�7s"K� �g��q��-җ�j��s��Z�aC�W�2� �/Xg�-!�d�ᤏk�H+�x�Ӂh��^�1�H�C�E�������ڂ�:0r��Y�1�1m�`�sY��Htm^<ޮ��vF�[�н�J���y�[Ӧ�g�S	n��}u$��"�Q��s��86�yS-mf'+�`���!�>�g|���s�}��0�H�j�r��*!�ݮ�[��U������D]�g�b�Mp� "���f=��S�	K�l�a�����ڀ�su�J������YX\���21�.Z���D;޲������ŌŢ���?�En����e�@� I��,Q1�rx %���%mLV1��jjy=-���?3#�
k"
+�}u�(dA������0te���a�X[;�v�u��y��@Y��a��D���i`V�7�v��Y��	�1��;u��|n���)�0!2��c��J����W�tLd�a�#=D�GjP����M�������e�S�cz�$4��J	G����O��Wҥ�*���w�7�����f䁦A�=羴e�Sl71�@#	19�_�����Y;,�_�������nB��NP�(���ao�@	2b�f���b����z�Z�2�[��T��_��GOy�A1�`/{�cQ�S���^�0^XN�TϨ�(�qU��g�0&����`�.o�������&;{�Rf(#�B��BR��T7BgH��%pHy���������S�<ʀ�I	d�@��m>�ca�5���� i�sF���?���ti�����m��}
[��O���r�$��-SV�^g�>]���y�c��sC��ބ �*��˟G��:�f&��-q	����\�j�����Rߝ�S۵W�ĬA+e�&������ۉ#���;L,�t��T�**�rJ) ���}�o+W�]�1|5��C��)�� qP�iXʫ���<R��!8��n�2G#�-l�x�T~K1�@��::�f�V����uh+�)�����6�S��t������&5d.�I�w#;^��cr��՘���S���"g\��$D���-�!�;��� �B�g��f���ؿ�e�5�<3�������O鲈^�����V�1�&��U��_��=��[�H	�!��o�wvF��"���5%��s?��m%�\�c�9��z|���^�8R��,Td�l��~C2)~}꣞d�����]���	��zh[�RJqܭ:!�|�tb9W�D�A�����]/�3����N�A_G�.���h��BFR俀^a*��=���/%���"ʹ��m�vo/�T9������5#�Τ���/����Q���/��ZX���vN��z,��X�<���	�Ec1�w��o� 5O�9�ӠU6�:�čY�*~�:фf��c_�~��6y�|f3�V~�j�x
GĳT�z��,�5Մ3ڸF��˨9�L�H���?���պg���(�<~��8P2�p�2z>������A���lc~�� �b�������!��'�F�׏�h �=~�/���tXܚA�G�N,���%��dR��D���� %U���U�[-Ç#NJ�NO�o-��H��o��.|<�U���h`G]Ӛ/K�p�48���U�~v�!0�N��$��G��`>��P�K��a�Y�e�^''�okA�=�D�~qg�8��1g�;"rY
�LE<��
�]h��>P�cm3G�K�(Q����=���#"��[�\��Z�p|��Ϊ������]Kv�����_�c��m����`|4�� �W�S��%��o+g|�_dr�p�~�)��!������P4ŕ&�W���v��܎���ɛ�L�Q�gQ,3QS�\qb�p�l�j��Csy�`�@@,<��*'G��]n��>h�y�����LS݅���5��K�y����^)��	�K��;��雊�L.��{��������� �=�Y?C��L�w�֡��+Cb�Q��gJ���3���? P�hx�?}�Sq�B!�5l� �@/B�+��M���m���9R� ����a�լ� �d�Q"��*�c0�� �Ǆ�����j����o�\�^�h�ߨ���1Kwg�����m��;�b�����������H9�!��o4ds!d�ye-�BGl�$����Լ�I̭�G|�FL�'��`��gQ�w��n���Я)�6�����`�FWd
	7P�!���0-&-�N�Bp�W�I)�<�ۼ�C���`ks�����]���K�A�u�|�<
#���[N�i|��cQO�K�{@�`�j~�l��Ր{�ʧ�2ӣ.�����Ԅlo˻�f�T��N5� ��͠���� ��U�"T��d��O	����~������n�P���~R_s��*������_-�O��9q69�
^�Rz��M�};fJ�����W~-`�nXY_��0�Ӹ�F�~��!^�:m:q��Y�����-Sx^%2���|�����˸���$Z�l{,7�	�\����
�k�!;R�D*]��T���Q}�F�^���ENC�y��aJ嫳��˂���UnwG��Gƨ��E".��"��C����^^g��&e/GՀ2W=��wB,�T(��]���m��&�.=8����ic�N����D	ԛ�Hhtu���S��,ā�[�3��&�8��
��
lY��H˾+g'����M46�T�=m�7�噘@Op�hM����C�.M�^�����J�好7Q��\ोwϕ/����C���
����_`�Tɜf�0�lQ�nQ�����)ZѺR�+��
 ���}y<j�KL���ɗ��'�?ft�/�!׌�7y#��!��L�:���%-}!��"�����T�޹ڍ��O����<3�*����PE��;ۯH$�� ����"D��K�����6�pf����x �"B_���U��nV���y�`�u��_�[�L� �F��~k�U�T@]�8��+=��=3w-�<CbxwY8���	�S]z5'����+{!|����O��qB�,�����7��c�-�Xk�V3���RM�_�fPK����2H =%qnN��Epi��-:(b Ϊ�����7x9���T	������}S�����l��<��Ɋ�J(� �*� �<z=��5�)۸�"e9V��\;�m��L��`�v"����_�sK�th�����r��z=��"�]�����J�k]D�z	��[�� W]G`��yF��ia�*N�7����[��-v��~��VW�tP4��o"���6�4]��`7"��+d{�kOҔ�H�t�RĎм�4�>t����	��VhmCO楆�S",td�&o���5����Qa�Kt§(g��F��K<Z֫�+y�b�$��J�ia�o�Y"|�*w7�����!�Cu��k�{�#-����IB($�FX_�|��r�rm�:R���]ppA$_���Z�V���/U���ƈ��;*��T���0�䬏��V�-W�T�c���#/����&	���'�F?�"�����d��=�76��0aɩ�WIat��qS��Fg%��̟���IC�J��i��Zԟ��ч��UԴ�G��W��9�.�J�A_�7E<����T7�y���(c�?��e1�^��:)��z�ɾ���G�v.���A5ʛ�	,x��g���_	)$�K,&�i@2�xA�g��n�{&�㌥�8Js&�
�
�?�X�j�� s��J	)�
�8K���E؋sJ�T)�6'�����uみ�#E9���fV����YdO����"��c���QG3?���%�EZ����q�	�\�/��F�K����~T�������`�034@����$B0�S|N���֫�><N���0v�F��j��XW��Nj��9��a^�r7��~γe�)f�.N�Y9��㿼=��`R���(�����UH)��^|o���w��T=��3�j��eC�O�����O�AN�q�U�Ƨ��z�Q13�g��������>c�-e���>��n�)�o�S�5B�߮w�y���(]�Ǫ']H����<�A���zw��.�~7b�
Ff����l�eN�n�%ے�K�X!�5�	�g����u}�&��>���CAr���?\�_�Vs�5P�!{�:a �R�Kjy ��9e��Q�Z��*�ېO��� �"���;�05k�Q���e}O��������Q`6�۳���2�I�ԬM格h���%�CrW��ޟ�'��uZ$���أ�y�?
I��� ���O�ܶ7NwnY��55�G:�����v�'���zy�L�lȦ�os�H�$�{YB���v��d��n�'+ޚ���,M
���:<�L��Ѝ�2b��Q�/�~�0�i~E��g����=.�Ĝy8;�,��^^�"�@\G�k?�C	��*Ȗ�#5���c�$9�aDG���kVR�֮g=$����υ,���Ӛ�����^�yn:��	�����<����cW�Y�~�Q�B4��G�����V=���(%r��v^�ԪG� S�T:#�Lr;W�Y��7��nt���q�ޘ��/=�N��)y�h������1�z�:Y�|Ge�^�fÎ���K���K�߽��|��+)��5Jy�46f�=�W��1��L��A��#o����?�C��Ic��6Cy��\��{he��,�:�R�Ջ�G�=��	M�N��Q�xq�<5�>�eJR�*��^�o��5G�ms���r�C.r��@n�� H�k��-j�w��bv�;)iK�Uu��`n�B���L�uF)4��p@�'<�t���xe��.��>|�f�l�'�5��>�m�I�6fm�ڸ��
i}�Gx�/߉�w��|߽vc���|�:�/^<�3�
��\���҈y�Jg����Hh�SN;��R%~A��UBV�$"ɨ�:��/�����_��&�-@Vy]��\����8bdCI�c�n��&}Sm������'�;F�dj��ynh���^2	 }0��y/?�@�B�%�qή8J��@h�CZ5P�+./9�����mm2'c9�"� se
a��䲸�pD6@��s�Hv�L�"� k*1�E�=b��.��7z���Fs:��O��L�woS">
ϸe��75`��)���5:Foo�f���ׄ��,"�+Q�q
nj�l���l�ж��T:�'�wm�y�9T/	PZ�"�,&�WN7��X*�O�c���g�X�d�m]�D	7W�b��t�S2&q�sP�4Y}�,Ty�TL_5�n_ X@���=���H<�Gcb�:���>1�<)*�x"�K�������U�%S6I��������VX�w��y�
dc�(��ދ��!Wm��[��\l�V�Fə��^Cji�.lr}��K���H/��<$IS����d� A˒[��7%�`����#���Z��r�C��ݮ��?���D��Yñ'��)T+	|�z8ͩ���3{/;2e��:��d�^K�_v�Ɉ�k��RJ�F�W�ճ2R{�@;�藀t�>��r�I*UFu?u��;���d�P�{B/�nH  �g�#��R&���t2�3�.���sj�)V�����[��&b�8J���jomb��> �px���b3�.'�+v�;�'7�����gˍ��S�f��4v��h aJ5�Ax�:���)�Uk?���>��&��yr��M�t��io,�����1�����(u+w�V�Q��ΰ�ɔݪ��茶��M����`sc�E�Qϴ{�o2���e���~��M�I���.��V$�-(��G�{P[�8�쑮���^a�x���Ͻq��eNW���X���t�Z/c�V��>���|�o��&����7�F;���B_Y���|/+��jb�d@�s���}�l���iq����UGɚZY���k�M�p�H��q��-إz��T�sa7�����)!a�Eg�	��u�=:��^�"��, Oi:�n��J��M��<L�[�%|�P��%���ap��[�30/�ig�Q7�y��mWv��ݣ؟��+��s4"*
��!�%�ʬ=@�r�@��^n�5��uv��n��q����@?9uǪ��BFe�Hݦ���yo ��s���:*̒O�'�~�>a�p�53�z2UuI��N���t�5���p���E�CibY�Qk�;��� 
�h���6���ͱ��@�')���q�i�;$������l�gr��<�oO��ra��@�>>i:h�T��:t��N֛�s��z%��9��P���gPT ����� b������ g�ã͍Re�s3�Hg$v�.�KM��l�B �m/����s7m;"�X]w�9�$���(��r�@L����{��*�h�GC�\I�Y�P�`�������+�?>ZD����5�����?6n��Ђ=�	p�k�hA����dU��;�-�0�MX�Qu�ѷ/(�"P3�&u��chY�eu�hR�$�6~���-YPQA���tXEλ{��)��8�.m�])���:ؐd̻y�f?�$m��^g7�G��oeQ|�)���t�>&��<�t�^Z��XApc�����������cO��I���c�w���;@O+��!���fM�c��5��6����>俔���#�>V�<�,kGwȱ��񦄾9�Wd�����>7�
 �o� �f�_$k�`��o�	�����U^�
��<�(JC$�2��A��!:~.ph�@���"ƣd9�`[B��ICݧ0�hP�N��(fzʝby/x$L��*nK����>c���c�Kμ�a�Ŝ4ߪ}�d��tLc�V�y��p��bY�{eh�FX���;�v��N�q=��D��?��EC1/BͲ�f�"�-�[�^��y��S4�e�¤m߃�m���wsKiV�������3}����rImF=b��H�>l�������b#*f�����u�����	T��&�]�)tC~9Մ+��S��*'�6�%h�Y��e��/��oZ���Z�G��"�ҥ�IK��x���_�v�'��}_,��B���d��L[m�`�x�8��d
�8�~d��$=a�.���t�D&"�f?�|!�? ����YW~Ќ��n�I[(9aq˗O`��ƷG<~.H��|S#�c�Ƿ,�}��nÆ^h�8]j0�Ip�?s��D�?T�����a+Ȫ��!��&�-h�ˊR���S�l
&'��m�&�����$
螁o������S>o�襘,-`G~��അ����ⱺ���Y��_�ي\3���D�����@�L[��i�ʝ���@��<�sy�e��R�^�r5�n}AbG*�\��q)���U��y�v=:R��5�K8��#��E�s�Gk�s�����hWR��x�Jx�������4| G�ަ�����M{z*`�j�(j:�Oz�<y�#�47���l��㓱GoI }�����=�k�d[�l8T�[�S¯ObI#-��6�}�⮥Ֆ����a���)�[O��ǭ�;����v���3�o�hǩ�n/��[�F��|��������� ]�d��AI���7Q�axc"���O��{T�hV���M$l��ߠ1�]k��Pb���y�w������&�^��=��.<���˄� 2���ʠ'3s/�q�G/V&	-}�S^n��(�w���{34��0��	v�F���lIE8Ĥ��X���_Á��=�Z�BW8����R�ٿa���@k�Y
��F�r�����
9R��:%���0�l`��_J��$���m<19����MQ">Vɭ'�k,�znK���k"�1�ez�p�I�4UF	F���{|i��Η��E#Lr�Q3=q`���G�`ڋ�ɲ8?����*��OE�y8�{�L����@
W����;�0�t�o�4c��$yّ�{f��Ԅ���%A}��%�F[�Z�#s�X?���k�Y�,�J�Š���G���/}�O�[���=��١����'�g�VH��N\�ɍ�^�\#@��`��/eMђ��f������,��/ �(Λ
i$Ҝ�����
�������ٕ�R.��M�`����es�S�ׄ��������Dho�
0L�#�
��`0p�.S��tw��Ј"}b;Z8&e.Y���ڂ�]i�\r��GGߒ����Ke�WbG-��8x�#YV�GnfGs�NG�0c?�I���P���!H������4��ω(^�$ߵk~� W�A�R
iBu�O�QJG���� Ѥ7E�p�0�^�����K�P�����5��3ڟ1-N&�v�@^��s�X4�0�OB��k�F��O���w4�J��Og��$Ne�k8��2IX0*�IΧ51��#�A�؜4�b���@Zdȃ-)���N��Z�ѷtӾU�Jd-���[)�6Ǉ[�E<�a�
p�G(���6|��D�<�v�o`�
(a�+0,D��4�B���~��/� �{�و���{�����E��i��E�^7��)_�hV&�o�O4+���v�}��a�G�˖dOhh���K��
��<�V3%�<�}��D�ISq��b��rKS�#���^�{H�-2�"��Jyi!�C�	���שg�g@��)���/^'�<`8!�/��AQ��55�Mt1�p�m\�k8~?"�����[�D<9�;��mU@����*"W�:_�1�\p�������hj�-��7Lʡ��բ�������F;;;_4���DxD�P҆h���7�/ާ[4�Q�� ��3���Zh����ϣ�����1V)3$W� ��g7:�,�O"��P(G�C�G������)ηŧ����~1UE\*B�De�7�f�w�t��g��ZW��O������p�d�["���5�����V��Ǜ�����[nƑ*��˼9},��H'����D6(��(Z���CX�9u|�i,����E㬯W]r���9�����������,�(� a�xe�0hZ>5�JT����;Lۨ[5m���bm�����A�4\.�D�-핤b֡B�!�<�Qz�z��t�I�w]>x.Z��*�t���?����66`�`U�Y�2�F�a�������'m)g��j-��(L�%��R�ɲ h}��w�'��	�/����^�J���l+��0:�q�SNS�_,���e�<s�� G��w�5��
��c^Z��0��I�d���
g.*���_pc�@}VK���z�J$�����AD����e��. ���;ł�MH�O�I���<�T�m�i�n�>-KKs
k�FG�̽'W'�yօ��޿7�?A�i�]m^[zpR���h��.ݪ>�a�ˮ�n�$�ưv��g��HY<���������A����d�N8�
2s")�!�|��)���`�z2���R��y �sht���w��b1n���߯F�\��ް��s7\�� �����$��*�ֆZ�뜁wCh9A��8�\؝�M��\�1��\,3 rD�:s���G�t�Z�����$���/C�z����<N�� @N��_@��cF<D/VJr,!�C�#�c�^�����= (�2!z�)��������z%.{?#Bo�5P$�j,-�E��M>b�]�F[���#lS��e���^ﻫ��5�VYz�q"�`�k \t�5�y�Yy�s�����V�,���\������N9\?�*H�)bZ���A�F�?.�����2�G<��ʸ��/AP�W��&WHb�Bq}�A�yl+����]�J��E�s��-��G�}��܆�u�[�tcw�b�����7�B�@>��gP��{6`k;��ː��{�B��n(1!oU�"or��a����|3�
���WvtU{~�� NHi���C`��z�M���.�ގ.�r��S6t؆a^{���z5�1yg����5N_}�2���쪜�D{G�J��`��W�ܯ�>��k�S�;��ֳaC���	H�9k�v��d�/�#@�i#m˻���
�`���U��ӂ�h'5�����H1Ә��L�u7�o����0H�ܹ��S����=�
_�\�mɏ�	G!X�o�������:P��Ǽi��2)炑L�l[�Ld�Enf�R#�x�u��پm�Z�S6GӺT/+���+��%���r���.�5�ag�la�=�yV��S1�z���M��e���^�|[�p`"
��E��0��k�RVp�������mHCW����Iŉ	A�S�WMv�@�^��/�yB��(��K��<|�:.P�H�tdTpS���=�/ ���t��Q�V~���I)��J�q�����-Y*m��E�2�<�#vif��)Vd�0N3��|"�� �����ڹ4����aɐ��V"��.3`��ײ�0]>��N�B`��*���o�)�b���o�q%i'g��QSmu����i��8�R{��]�Y���-���5w%���U	Ǯ9H������IAM��y͆u ���+ـ�I�rf]�v�4�a`��	OK�:;7}k�Rl}��=�*u��T��y���~�3��Q����H��T��ѩ���r�E��fQh�sQ���ڊ(%�U�3l�JL1&E׈�At�U2ȾH��3'�~�d��^�=�=�1-�E��:pH�vcį�']ܙ�g�����9vK���@vP�|�w�]��T�;��d����M���;��D378�k�R�B��?����4��N�s(�e�N<{q����0l�t�ВҠ�a��q��L��4��S8�W^�׃-�},$���5SUPZ,��\�� �Z��B�)+�E�����A얚��R��B�и����"]��>��{Q
�gx�\��a�m����u0��W8�����zd�2�?�F%��m\���.��Yg�G��Ɓ`O��܋ﮆ:紵�o�V��0W�+�?aoI��,��L�6��3b����/0���ݐ2�7K{\_� V�;pv���*��N=Rd�|�D�䜖Z�D�~�ǘ��&�C��y�2i-�-HE�6;�K���]nͩVY�-�f�
�s�!  �EM�Ab��🦗�QX�X2f�θ�N��n��-f����[j)_������j�P����n�~/7�6��x喦 V�'��a�oc ���������=��B�`��϶���
�R&�]�,��ʝ�������' �����E^QӻR�wW�S��i�6�.����2�?k��r<��0���gy�'�|�p�:qఠ[A,NX�s���#S��"��� �؍Ic�2��c�����(�j��0��M��,�P���i�W�A��Y����P&@��g�X��Fv{=w}�e��É���A�̄ݑ��o5�ի�lK*[�[��&ŐPC�
T��������� ��UwL�>�8',��0S����z��R���A�ς
t֞0��8�H�l�;��}s�Xzy�G�)�!�!�x=�Pr`�b���oF�ȓ�Yb�'��._�蒧�O�̘��Epfג�r�hhkY>t�Ȏ2lcyִ���~���Q�^f��<N�\-!?nvY�*>�Aп|��t+�3>9�����U�W�U�{�ń��w�<.dM����|�GI�:?|����@� +�ￗV����M#�+y�-����B���%��
z_!���LLz�t1#�D��v�j+ K��đp�[ߣ�E�%옮�('5�O��8�Tg��+ji���{�҄V�Г՗���d�6�'�:����f���x�я����k���M�FmSy~�K ���jZ9D��(sR�N�N��*�2�p1:�n���x��V
"Yv����8�W���=��s+y#j*KX�R{����s��x���7�ڱ�E�#��R�=�|�0������s����T�Q̭uL�l�v�=��`��ܐ�8m�q骳E�֨�o��ղa���Y\я��.;���^gG�u��zR��2��¼��pzC�T���R���3!�Q�GT��B���rK��D���պ��-ʃ�[�����C�S��R���S�^�\�/Qo2��SZ�<��x�*��9����y?\ˁ�4(PPmq<��8
����4����Z@\ˌvx�qḱ��UW��w?�|둒\��<'�%���8RV���q�w�����;��$�_T��N�W8��Ö�,6�N�Q����S2��d�*+�+�-����C�!xq�`�#�"G'h�~
:��p�R#ؗq;�F���S_Md���<���� l~���T2��c5�e�k ���zn���U���@�|�Z�Qz$8�X	����Ng�+>���Iyˆg��u,.F6�ީ�B5�,=�Q����5�l��+�B1$�zգ�c��~�u�Bke_O������Ƙ� b��E��X7�Y�w��̠IJ���c���huu�	�i����<�
�;�v�-�F�i�n����z�QO��v�2c�F#Y�:�.b�Ǩ�a�\��3]��M�Ѐ�	�^/Re�?$wQ�[_�IIC�_�G�*�K��U���',�X�3wJn� �Q�Hʹ�}�m���f�5���N{Ud�_o�R`��	b��E���������`�ֆ����}�t�I��K�a��ZAQ�.ɛ�����v��zM�1�{�ij�x��,Y^��Jk=��zp��6��+#;�5�e�/.^�;����]*���O���5J5ֱb6{65�F�Ѽr���M�J�z-��<�W����7dAN��E��Yt�r|Ck$^2�z����	�^<��1tWbE}:���~AP�����y*��"�I� .�S�J�?=O+�[����� �oG3���_fn�a�mx�#!_�A8�WÈ˱�瀠���ovU�!|�, >�)&��XE�pNN�ɒ���mй�+�i&mSr��ӽ��ERsd6׫فQB��?�|�)+"�Z�,I��7Ȓh!��+>$�>�h�rZ[ҏ����-�^l��ڱ��.(H度����2����F�oI���V7�J���%�F��u������t��@+�XzVOM���7�n�%�� ��p.ږO�,��	�����}��D�ȶ���~%_0��f���T����s
ee�h�]hk�L{L2�>6�[�]d�7ZqX;�0l�\E������H�MhL���G�	ԗ���-Ώt���/��p�4�h3k�k�k�u�H���N�i"5'�A������>]�|�c��w(�P�LI�� jX[��|�cxnU�M�J�f�'?h�r�+��9i���{Ձ�`�?�Ў�j:5�xp���{u�,����Y'���G����(��m�#(K#��S-a��\�MC�P���z�n!s���m���p�X��p�#�Yb�bE[���G�8?�Hp�Ӈ=�܍]����kTEG����ʁ�̼Q%[�Z���4q��jMD��'��������x#,�p�
�Sc���$C�m#�K�������g��E��ٿF���}D4Y�:�=Q\`��+@GƏ�����|� �#�"���>�4�s#P}�9�9�ñ��G��m�,#�$����T>e�R:$��SsiT 6�J!���[�3[1��L�~䭸�Ŵq���d�߱�����eU.C?���ϯ��In�%=(pUj������!�(.Q�)2\몡�^��~^�s���J'^�G:�u@�V}����c����ٳX����Ĉ/�[��P���B�o� ·�׍��7�؎ Kı�		�zBJ�-��*�ݽu���M��1�O��pY�
����v�!��H����M�-ړSZ5� <@h��w�C�ftS��}�ᅛ���S�lx�K��w�E��a?���@�A��Q����6׈;G�&i��'v+(�u+�bˁz��7�s���?x��EԬ�{�^pX}��c!�W��R�_6Z�W�J��xO�a b�"�ҧӯ6;�91��E%��!'��VSVG34z��A���i��ܹ��&ч[�"����9P���!g˵ ^֏�l� &,�qt���i�K���I1���$xA�&��&�|tq�np�#X�}jl+
ul�� ��)o^߷:�'uԵI \�M&Z�l�{�y��G6�>r�ݒ#��A�����G�)��n��~�ya�UmL��Sÿ$(❓p�ňQi����k>��Vm�I&��z��4 �	����H��I���ة��@	'.p�eh�x�'�W8jW�����О� ��i�7ۧ0�!U��h�u�bec�2���?�!��*8پ�.��^Р�r���?�PH��ќ;�B��#:�U~ *�_M4f��1J�u�ґ~����G�7�#$��?�u8$V����L^'^%���� &��^#�[mH �'�j�am3�'-wud�,<nA�.2-�Y�£V� ^�A�@'#���ߣ3��@�xz�	4��PZ+ߔ�L�_�����-?I\,��
�5QF$}� &fg�+S�߯CW�Vo��|�^Iq�4!�Vf;@�6���� ����mn( *����<��������R)���X[9�����,�3��;�f��1�B�P�/"��/��U�����D'�X��z�_RBQ«�����Ʌ�$+W̗��4��Q�$��{;Ba�D�"[G����T�/վU�я�������$p��D�p������{Q�>��|o��H���^gB�P��_��R3��K����0}p���k˻�.���T��Ⲍm��׮�8�'�%�4� ޺�/2^w�֬yqĮ��j,C���M!F}�Bݿ���3_Sz������%#��Wt�Y(�:T7��F�%N����}!�h̓C
�����^۲�)�68H���x�>��Wv��	�.�����I����i.k��/�{�7�2�<:�!h*(�<g����U�a4�Nu{�b�{�֓�~I�6u�R�*�����ʁ�Xyv �a8��(��b^Y�g����/	��@�+�.�`?���kgq�WTw�+[B�;�Cf�| j�u"��j���^oO�wV�2�p"�
rkB��Me	���$�da7.�q�i���d��y��-�c�j#�T8��N|[cv�G(w^Z�`�N�+Q*#�_As���]0��ڀ�o�d%Rh��4h�)V}��q�E˙�WxCa��r܁N����m��H������\�s�f�ʔ�#X��j�A��iG��#����)m��-�i�YO!wK�����{*k#8��#<#X���ʖ�����Ƣ/;���з����S.��ZL����V�B7�D��ϓnD�b���厮�z����<#qm�tX?�����V7#蓪��P���o����Ste�sA`�RK���(��k偵)ՖVa�`�����$�|�k]��:�o��W�r��f�t���Z�x��s�w�Y;}0pzޏY�~��A"���V���4$^���eF Gڤe���ps�0����%k��{n.�qĕ+�fm-��j�C�O��Q5�.�k���{��Z��sSG|��P����Z=�m��&�W��$� �uhY���3Q�B���P@㝫>ne��x���N��/�+N��d��=h_T�]��ɦ�af���K����6u�f�w�Xs2\��w;Tg)^�+�2Ũ�{6�.�e}~�Q�+�M��� }5��U�X��q�7 x����f���Qo��GFD��_�����'��4Y���Lo�����a1
�`f+G��z���I��Pd��	���e}�N앃
"Zm��c���V#s7:�fXIk��������\�-�ɚ�80����'������l<o��A�<n�y�l�Q�y��Ofk�wt�H_��
7l�Z��:#���!L��@d�ӣVt�����ކ!�u��shKNͲ��\Ԛ,e�SN��Q���)9=5�f�*�h�^�0�7ģ7aD}0JÕZ.=1zlWAb4��ԅ�E��X���p�$����)!R��Ax��W����D �ьQ˶��,�8�#�~��@S�'��}�G�o��Q����w}m���B�49fۋ],��4���o�m��w�y�@T�G��A�ET�\=�P[�A2��{I���`��٘����x�Qfԓ\�{�}�����f2eCض�J �#�4U0(.��N�Qq�ﳱ��\ �d�'�h2�_���H����38��+R7Kf$W���*�OI���S_���$�ov3#�&Ӛ�r��B!�J�k*�����D�ϩy��ҀK5���A�h�Sj�������;��m�L��5����Xz�C��S8���m�W�
2}���z�)�t�=%c MHő��g�N��6qu���x���3�)uo�!7���-�o���[���cX\I��sM�tf��↟R�'꿛�V����zJ_Ż�o�T0���k��H%-�ϩl�VP=��nX7�fz���e��Ikr���������o����M:ʑ�����h߲�����L������D����uN�k��r��$�)&)�2,�I�<E�S�j F�q�l�Y����<t���~�!��X�O;]�ҋ��p$�����@s�Q�F���EP�lt�(� Hf�?ѣ�VR^���g8�>���;��C���>�7���i�ON�O|Qi0�s%��}k̪��S�gE�XVjV6��x��(8��^���G`h���H�v������10��S D�ɩ�^¶�!B�-��t%�,Nx|p	2/�^)E>��&0�X���E�����w��g�\N'��n�H�f�)AwH�	Z�#8<,��D��$�l�A`��8Q�����=ߑ�MyǫŘ�����l3E� ��6�<�=��p��Э�@2:�K��0�f�&�3="��p �}6�gK���n��2Z�:�U؟ۛ�����T֪E!���oP�Jg mi�u�U�^WM-��/�HB�AgfH�{
���|���21�b��B73�ǡ"���G/���0	���y�㵠�6uv�`�r��R0�ׅ[o�V��ĈWd�ye*� �aJ���!C�t�1�, �\�5k޳�E�R�ѼU>���Ӳr�le��c���O���C�e����I�^�t^�b��)fD�Ʊՙ6$�9^�g���{%��$̯�y^^��~ ],$� |�#�<�<��/gh1���>�*�ғ6ɰX�v]/����%͹�;���EZ��'��~!}�i�{v�P���G���"b�2�~�)A��^�W%�cR>@T ]�x��q%���6?æڛ��lx���(0E����慓�{{��v����(�sf���$�Xn$*5N���� �1�=wu��ѓ��?hc��c�ցc����`n:V��)9���:<nVx��xeik��3{N�����D�#��C.lM�zc�E���YFtB]�N�"�88kl��Ю���KA'^SO�<��:�$P�0gb��{� (�P#%�j{���c����q�r��>?*�����awӌ`ם~}յ��1�5�'/�^(��Hq�)w���mp�px�R���19��@�MEj���eɠ��y 7�>��zO�׈'���`k�C����jL����h��ɩd�v�w����V���0�^T�J?Gg�c"����dG!
>�N-Lq?�+�hk����ہ�Ȱ���X'�\�4.Վ^�Kgkt:��:�&c5�7>�IF�3]FJ��L�?�����bL��<"�b�GdM0�.�Ya�685��E�q�Tߍ�c��F�׏�\�$�{��p?�z�*S�7�%�:����=�T7��Ia����Ǣ ��+œ����=Zy��v�k�Ē�x�?�a����z!���+�+T|Y��l������!�SӐ�۵`�w]�21.�L�
���i��-).�˽��ƹ�8���!�%5'I�vyHs�>��ۺ�E�`��5�Ƀ��g�����..���I�m�k[��'$���L�a���F`Hhrܛ���@�o�+��n��0�$�
8�����T9m>.O]����"�v$�ʢ^����VO��w��6uI�ٻ��Ѵ>Hp�2d��*�x|T��$;��s�J���"�ɺ�p���f�e9\S�k^&��_0��
i7L¿4��\=ݰ�^��#m����-c9(�pma�م���('|��6�ԁ͕�Q��F ��E���UΟ�;G���W?R��S�P�u�n�iXç1�FS�Q~�e�rRg	&:Wf��'�6�.�ɪS�C��C��pd=�tmГ�V&,������M�Xt7��4w�+�,�V���n����'��x�x%_ g}��Vo�`���-2��ۛI�
����S?.��^
���\�(*ϬX8��vMԐ.ϡ�sS�����\�l���BR����������_#���#�1Z�W�ny𗟒��-�'�y����/uZW���m�hx5�����_�4��_��š���6}������f�f"3�įN�yvH�B���'4A=�l;��h��9�/�mL�W �8��gV�3�z,E��Y3��y��:�^�	-�c$�b��?HڿRD Ŧc���ֲ�:4�>����:����w����>$��ILt�?������y?\L�,���
���X�T��=�2L��v���CΧ��ͣ�ܙΏQ�Fٙ�H�n��<����|Rn�`�^�?�����&Nu2�N���!����1_,�m�k/߶�Y�%Xș�����.���>dp��$�	�T��f	�bw\�K5k� ��֍��Xj�E���A/��TFW�o����^�)⳨/���Q�)P;z��UX����ۂ����q��^���Xϴ�Z��D�#2�Z�Z�y��\�~���\;�A�l;!�%�������ڜ�e�j��)j�����e��/:~@��,A�#{q�W��v֟�E<c(=� � ]���hr��12�sH�A�	�ف�P�ڡ�T�	�[������"p�-и���6(����rPbF�&)�G���C4f���=�p ;v�*��q��Z9s�O�"����q���Y]G�%��c4���p���U�n<@g�� �e<�C�y�@ 83���?�Eer�
o5&,�?F�N��&�=�n����/9	������5c�M��g�f������y�|c[��QN�̭���EkZ1ڻ�A�@i��N�u���߂����`�N��?�mXt��Va�9K*d��b��d./���{�g�����5X4y���=k��1���[15����M��G�5GG�_�}bʜB�<���ڃ�eƴ�̘d������s�$m:k,G�}S�ە�IT��t������:Q+�s8���W�^��
О) �+���ld�J[�؝u6�Rx��}1v���Zb��ڼ����WB���b�mN��c��������ʥZ�L�
V1,�n��O6u5�r�og!��а�m��d�rH�;�bľ]��Zd� �>I�~o^��2z�L�l�af��V��p!�s�@ݨ&�?��J.{&w�Y�Ms�;�Lo�3i@�k�;Ԏ�3����e'pZV[|vk,!��5�T��z�)���F��d��~��J��mA�e�I�G|G��I|�ącB;�7��� xDﬔ��l̎n]���B2*��&Ξ�����`�{��#���D�vD��ɳ�匀[GN�q��^�]X�����F,��LL�T+����:�	F��0�PT-�X�X?4�"�/�=��;�쟉P�����?ncs��4�0cUT�~P����"�lc%%l������!����
��E�L�e��=�G����,bP���I��+��R+�o����O��UJ ȕ��ZVr q������Y,�P"����8jTc��osi���5���x�C>�yD$��u�o�0�zy��D����й$�t#���,�V���E�C]}�&����8G^.�^w"��g�p����t���7LPD�A�>��Ht�ڦ�Cޤ�/_�X�~���[�@����:�_����&0�s���(3�4Ό4"�JL�����(�1��YިX�hdo���v-�"}�r�M�uݳ������N���9��8ZhR!2����gyCC�N�Vi�,�db6�8�2^`9(X]�]���I�!�ך.�FDU֖����Q�n"}��s����o����A��;^�egN��?�=y�iD�0�^�"�.�{4&��!�@���z�qW�	�����,?w �Z�3/^��xkZx�m���ac��)TY���}D&�7$�M�U�Q-�2��H��|mv�{�C�t��F�L��6��zБa�~�o��P����lx�O�>xSzcR��r_z�e.���}�>�c��LFt��| #�@�]j��:�?,!�	kީ�����h��C'L�pT��=�ߏ��
[���.ұK���ֻ{4�sD���|Y#OQ�� �qE��H:
�$0V��!iCd�/���j��n�҅6(%�9���Z��w0jc�����ŊE&WF��M�h��+#�V9�}.j�'h �d��P�M-o����>+����{���?�璧��b��L�8�lù�wDW�A�!0�å��g��Agh� 2��d%�~��~)sqox� k<A.���o��M�����Q��_omg��F��~^Wp��B�a�:]��7�@�[�knGSכ��6�� �Q�rT(��bwZ��\��m��f7=�i��E�u�
tܐ�I�u������/�I(dY����/ſ��}���ꞻ�~џ|pM��K�D� �
��.l���zlsU> �������M��� �	�	c�J9�G GkH��| �$c"�9����kL��ky.���qϩ>����K���-�&G��$0ꙙ+Y�s7g}�i5z�̉�JA������:��\�����Y6`E1��ʣ�j�L��Jp�c�X�J1;�O.�5���2`Ђ�k Qt��Hz*y���J����=f����2��Qg��r�`W�Х]jW��^�,7ŹqX�p6���!������!3��d�\>�y>&��-�xVP�r2Zx���i���A=����!��mwS�ꖸ��ʑ;�/Hk��MF@��\�B�ۻږ������ir�z�Y�[�lw;A���.F�`/�����!}V!�x���(��&[qm�0�RxV��Tѩ5�N6/����"a�����H�.'��_+%y�+����1��=��"�˫�B$n�V����E�6<	�ۉ�V�L)����3�F�6�y��pR��N��=Q������g�)K�hO�!'� �K��o1h0��F.�ǉ���ׅ�����]�R�}٤b�B`i��Q���I�3\�[�0D���Z*/31/�р6��q`�t�B�o�7���'���1uI��6Ǆ����w��ta�P���@�����fj@�JzEZ�:3{2F��]�庡;���#�b�!H��^��nn�/�$��b�������Ax��#��#��D�=煘������^�b�;,#�=U��k7��V��ZuEs�R_-/����bfoR��F8��F�>�d+���;@�S��ɠ%)M�����������U�֋.�jnRj@N�1ִ�c�<��Z�c�M�Pt�2��b�g�����S�|�7�V�E+U�`j��0�5yю�j39���ܥ79���>�U&7G9�!���m���7r3dt��MA�d��G�`>��,���Y��-��I��j	.F`��Z_��<J���E啠����	TSeW\g&�c|�\�(U�Ch�E��ma�j�8�J���J�[2��`	[&���vyTR���(��?��-�A��Ld���~��* Mu� �t��!z�o��HPp��]j�� _K�ې�zhQGbbN'o}�A�D�JS�q�怓 �3T����%�Ă�'�^U�g.�G��gʉ�mG�4YJ�GI��㱈�$z��X�?��u@W�_ዶ�9}O;��)�a����ѡ>$Λ�O^�؋I~*�'>wm��9y�}�	��dD��(�+k��Tz	�fR�̐)�WP�{}w�t�Әu���G�/W3��
?M!���|N���}a��������)�=�����C�Ȕ&��F�(rR+�����\p2�&	�������8[�7���f&=����a���4�Fg���%V���l���Lf+r`�>�d�u����+C���n@A%S�`&LQxJ��d��ӽ`���!�Y��z���(�] �_IUq?���{xu�xd�Z:%]̆�©�&tPe��@�օ���?���,3��C�zY��I5�M��a��`��	�Q��\̈́��ĳ�Q�g�J�W��P=��j����n�]��ՓWv���}u�)g��C��Jf�n��-YIe��`���0��yK5����
nH����4��*�g�� �����a&ߙ���<�X!Ŀ�a9vW)���0�U8K#ǡ���?���m�9��qN��=���E��|MlF�s�Bc~qFa�#@f-�L�-0@��$I�qD.�B�������T��-��-CHioH���ɔ{�����
�S��g{V�
����Nbma���fqMx�Uc@�<C��Y�&��q�2o�F	���	Ђ�����G/Dt0h~��u!Vv6o �K����{��^Z2��+��#�@�mrFl���G4�G��:��ّ����C�R*OI-A"#��^C�6�"���9���HX&�S/���݆oZْ�I�!bSJ�A�2�=2���;�r���=�yj�	5���$,v���oP�[H�V.�A���Ոs�� �p��V��aW��
�y��we��q�_r��ʍLVjĥm%%������d����{X"(���d24vt��F���i4���Z>dV��͚e��0�0�K�;�P7TZ�&�#E�׉���bdA��N��_z��&��ֿ�M�a�%g4�g?�����[��>�G�|tÙ�\���&f+�!q�aK�CQT�)O���m�L�u���s][^�Qص`�k�O�j%�Fpњ^����߆���umQU']�#���!�����Pm��޸%n{6xN�����RS܆8���h��� �'|�\���ƀe�'��V�d>_c�?8��Ah���"z�Iɔ�@a�+�߁�N]����> ���>\ݷ���]����+ 1U( !���\����k�� )��,�`f퇡�[���}\*_:�u]�@QHٛ-0�:f���l�c�d�H����'���}GɈ��z�
�G�r�1�x�-�h#���Ci�[''`��w���̊i� �=��R�1��p�o�*9���;T�uP:� ���rv��W�$�+3:�
Z�y5 oX����Lם-���"᭫�&
��Ug�Hw�S:����`��(���I�4L��7Jm;�I���@>�{к��� �:-d*nX}�_�%��J֌NJ^W�y[�#�ˏ��m�~��[a`K|e?�,�߱D�IU�`J��w�&F��8��� �Qr��}�������3�S��߸N�-�!�9��;����/��,���#�Q�#��%_��3�7��j��7KW�#11M���&H'<���#9_�!#i�&� 'B��NaP޾�o�ң�ra��V������
�
$N�4Q��yT��a9Oj��������w���QJ�߮�<g��έ͕���^-oY�x�{o3<�C��e|�d
j@;��rѱx�OK�o�w�".n�G� ђ3E��.�f��@���:Q�.�$�I�΋�r���@O��*���	��<?L�JuY:��qf�|l����,�,sy����i��:A�Y$��c3���\;�n6����b��xP~�q��d�N�j�����T�v�=ߴiwkB
�d��)�Pz�Đ����;S�~c"��duJ��1f�]��A�{�%��*�k^2��������2�Y%��B�wܭ�,SOu�0�g�@�}"P��CHa	t�)�.x�ٲj�@����L�(S��K����ގ�SK3-�c�c�wE.�'���p��u���5I	\����M��Xqp�[��Xv���}k��l�@�88���WU�3B1������ i�����U[o� �azК�~� ��H��� �5K�-�/���+�XF�I� &�Z��7gR�H��+���Ot_5]�Il���ځ�u�6�kL-%ݢ��E��+�d��9�O�{����V�m4Z��;^X���mqjR��'�z���s�.���:/K��=�Y��8��h���<bG_o*'N�-����_-sqe]@�b�bG�?k�S���Μ�T;��e�'=�`��9�Lh]�;�[�o�5S���@?Aip��ӭ�;��O	DXTܚ��P,_����ͦpL��U�K�q��_ ����@D�t9 �ѹ]�^u���
2��&�Zq�@l�#c�ML��-�S�n��y-����mg���0���1?���"��Q���� �A��R�������z��xj~ ��U  ^8����
����#+�(��d�HH���(+6~ԑ�l�:�T"�s�G�M�O����H8-���č=������%�k;|���ޮ���	[��a�/��B	�,LpQ�7�b�aVkQ�r�2���C?cK	ʎlr�V�ŎT���\P�(Ũ��poz�ATgo_�����L!PC�2pW���������x���0=h���~�@G�;�[?��⊮�Cq���/��u�%UzϜ���6��z�.3X3|�N�	��x��o�_�\�.��#�P��pG-U��h�(<0�o}�v��×Pc0v$��;�������\��M��a�oGN@�ѓ+̛n�U�K��Jns�Zj~��K�y��WK��R��M5�;���	-N��}�<���K*�,��(�����M`��8ۀ���7�{�>�p41-�2�WN��Q"�c�f9�5�h��!`�3%����,�`a�(����g[�sț���k��b<���xS���:�Bv�ϭ:�|�̥��*^j+�Ǯ�d���Ff۪��a�!Y���-��y�����@�}u��U�!�Զq\�.RR17��Q�!���T�8�:�@��Ш��-*`=Ӳ�����H�!Ź�pG�u�	�F�z�qX�l�]=4�q.2zSg<�K�q�P1�[�^D~
�>o���gl޶�����q��K/ ���s��;�#) 0�����M1�c�m�.B���g��Y(��Q?�e�@��,�ǻ��:��,[��N����gPG��n0�Y3�|��t�4$�x7��_��I��0���1"= u_a����H�?��Ӂ��"�./��>X�_���_�sb�#�O�2�7���W7O�9�'8_#:�O�;a���yĮT��$��N~��4�@@���7�ﹱu����ń�~o�ap���Ҳf�G�ƙ(@̌���Ƅ����Ln0O���Z{hk����;"ݰ8	?�77U�	�����������穭�����ܑ����I�i��
�Z!�'�j�mɲ�j��1H!핊�;p�hdص������� �`h%BU�(�[{��,K��+1R��T��MA�=�2���X<P�^Hi����5�O����d��&�	�#{
��w}5��l�W����[���qv�#7��.�e3���&����"���'�T�erx(������K�6��ބ��%2}�ȔY6�r�d�wm=�:羮��%uM��+���+��h	�Ϊ5���tے�� l��i8�"[�v�����FeL$����|c�����U�����x��S�eȯ�p0���Z�C�>u����j�#��Ĵ����v�(�d���X�T�KKAy@��h]E���M��0��!*�Db�μ�·�#�f�^�z�X�� �,ƠS�!z��~�����"��O�~�L�c�yu"ۨ�Gh=Mz���1�m�]ϊ�|���;�>�N(�Գ��\-�4 �NY�^,r8TW*�A)ÿ�f�
�K���9���951��Mnxͣ��XKjQc%;�������Q�aeU�F�.�V�uϋ��y��+�$�[9�(�8&�f8����b���,���8"���W�*u;:�
pF�q	�8]��Q 0��A�u��
��?�9-�H�]�>~|��ܔ �<Ib`نɭ�FrB"��C�n��[��ªЊ�k �I��*=�(~�B?��a�o"in����9��2o�J\�dtXbAe�>���Q�u���B�C��^4W63#��1`�i��� ��W�@ava��3�kB=�+���Bb/|c6ņ8��{׼oH(��]�z���L��	�3�����oc���j��?���l��-U�hn�Q�r>E�jc0�)�[4w'�iE�\p�T�����uŧc�:�R`'�4�
�������Oc�������awa��j��sox>'+�[lܪ���2D�[���23~6cY7ǯ��j	E�"�"-盏��,��2&�0��!�ֳ���([��M6P��h��hx�ҍ �>�Ns*Xw7E�)���L�6�>�L����Qt��p���	H�G��т��0w�TD��'*l,{�פ���o
��B��B���ٶkD#⦦`�E��e�G,t����ʛ��V�K<)>]�S��<9��Y���k��?�А�u#䰳�&���<�F5�f9�#f����Qq��d�'�O�(g�d-�٦Cw��0P�k���)�t��OQ)�=��~HZ�c �t
D�O5������X�L�r.�:�|U������6�e��i9��ˍ�
aLI[g1纝�l_�H�`6�l�J@�d;
@$a�]}��]�`���>f��YP�Hl�D�d�֪�vE����:T� ������p/�)���ƹ�Jp�y�]vL�:#
���K\N��{���(��iGk�� ��D��-�XS��*�PF����@�1ά2�F-� ���\'��^Ͳ��	��!C�iE#����r�t1怮�T�@�W*�!�dy��`��|�ygL�X�k�����$i�:���U��5?ט�<Z����l\���,0����g? �^CW*�_{�A�A6��~ӱ��7D�[��u�S�I��{f����M_e`8�>x�_P��@�,au���ѐvL~|JW��d������X�|��U�_��e p_e�y�km�U�C Kϳ���R��¨rxp8�S�r�c[�ɋ�?�Qq:���d)�=��G!iQ�����`��#G��}���{oLpWUmije�_6�}�{؄�/4�#�4�m�HJ��Z��N�q����Fٜ��OC?�-���V� �7Rm��;���	��%[��Dr<줚������maS������z�n�q��Y�֝�)c�v��Au��u1��Ţ��z֒�(NB���V�9�H����z�l�������u�r9���n�IZ�#Ҟt  �E�*GSb[5�+���Y�mgƀ���n�t�GӬ9^�3���I����5d�\�%���oޚ����P�B�9���~��Y�r���i ����uѶ��?�,.����/�$$�Ww-U�����eY�`f��j4����]Y�C�ڤ.-���Ӵ�v�W�#�3�s�܍��9����iQ��2|�0��;�S"I���Z�!)Ъ)��]�HT׉��a���'��/��p���|���A��C�Oc�CM�����>���"o;�r����(`v�2���	��2Myu��F����]����r4�N29�i&�KX"��a����3�g���i�n��2�'f#'��q��z�S�!%mH���]��%�^����=�A�Se�mj�b�3^�K(� ���w� ���B��6����z|�������=�S�+E�� XT$؝�5B�+�=ٚZ5�Q-d�|��_��B�>�����i4Ή'2���`��W'īr{��Y��3S�[v��@�e�+�w`�ºj��$��ɰ��q.�J��K�g�3hH��ǜx��J4q�p��}%��f��B�RD/�k�7O+��z"�1�?���4��.d��-�.� a���_�0W/M�e����sվr�
I�Z;��N1p_ỹ��l���}xB���eic���:E* �����|w��0�swsR^Ct	�U�L���a:1Xز������Μ粤[�m��V�'<R�?
�Gh-v�E"�FZ�t�%q���Zz�aE\�u�d72!�k��<���L�*m�Vʔ�˓����UV0�^�l��$��.�&���6[Efij�p��ULgv�kr�[�.�:��=��^��H>?�V�B���@;N���G�znf�	z��^�e�0��O%��궪(��Zr}��_��c���D_�_����^���wn4�0=�KD(ZH�GV�
��B���W>�˃v���vh��z4�*�ubv�����V��p��g)Z����.7n���q�n����	�G�Ui�͎�5L���ϝ�_�i�>2(ξ��{j� 1rJ:d�Ȍ�$R~B`�޽�;�]4ZZ!}Y��Á]6�q�e���f)��z�# $OrZک�%1��F4rS_��	ۅ��r��i�ܻ��IS����5קp��54ߺ�5g��	8���~`E�4�옵��<�C_I�xm5�q���;����Q%�����5�H}�}�͍�3�Sf���\�*4sʿde�&��*�;��_�B����v0�x ���]yU^�~@|xa�����<ی���i��N/R���r��B����=p�S l쀅�t�)�ivb�+��nxV�g C��g~3Ap�W�z�-[�sO�d�G3"��(���J=S�W��ن��r��fD9w��.�3S�X1�����)��!�A[�A�mCK�X �!	�R� GI ���Dl����VI�<��D�38��( �l�^o�.�Ǵ���`0�:�(D��镁տ��*�@~�C0�g��_�daL�A��,JH�"�����,��)�~𳑛ʜa���Z"��{������Q�Y�wvv��W�k{�aj�=Y��w1�ۄ����]w���]LW3�8T0�ɡf{��fo#;T�� tj�-{�D�?��*���dfI�k���ơ��������qշ�ˋa�Lo.�\]O�9�ߒ��Q��|D^!�c�0�|�OPU����o��-�	n�� $�{�g�-�e_V��^�{�T���_"��x�l�����0��LA�p�/�,�݂����m���G��8;}�6�;j��0�\�� q�u�7�u�a'r�ZV�񙊴�B���8��Y+�6��E�ghq�Ҟ��A��K~Z����:[:5�5��>�����U�@E�(!��i\.zܨQ�D�K5^pq�,�PΏD]�Z�@٠rv66��Z����UB���:Sp�����AV(�n�o�oy ev�=t=R�A��?8����'��<�Ry������ �z�b��xxƀ�&�̳��e�vʹ$�(X3Q�����/��: �i����<4F��<���3J��4o�^*�g�h��{�n=�wQ�b�>��K�'���!f͡)�� �����H�*�r�t��F�Pbz�!����sENč���ݙ{�baa�V�@`p�
n��aXG�LĚ�""K��;̗�xo��Cn�Ch��j�q�@H�/1��[����w!c�O<�\�;R̝�V�+I/Q{[T@3���Z����~������g%qQ���KԸ$~�~*e�ʦ/p�U��*o�d��)�/�*�_	�o2*��Ƅ媀Wg{��e˺���u����m2)X��ɻ)�7F�}�y�hK�cX�[�����P�u/kn&)��c�.��P��+�Z��f��+39	Ժ��f��Գ�h���P�]�����Uk�,���3��F9�	Ș��an-�O
�o1f|���QZ<�o�]�d�����KZ�vT#����-%�����Z8��%T��z<f�+,�x��o����?+�΁�z���0�#�7j/��W�~=e)Z��4�!̼�mE?z�B��G�uE�S|������jUq�����'{~C���YF�kb��ʆ1���<�!G�G�b4��*��(J�1����	���ݒ>o�Zd���E�l�dm9� u@�Q|.5��n�	;�cJ��R{�
���Ȧ��zv�[����xP�SM�9A�O�'(�
�_��IP������.:}/���swn�=�Fސ���8���У�T���<,��a�kg��rX�����0�v&(�����3i�{�i�-�X�K��1�, �r�b��-�2��ڷj$���G,�Aw<�5l�T� ��]FP
��2I�x�C�05tԴLQ�^|+RgzJCB����W]������B��4�\�.�!�u�ܔ�$�t�κLտ�'��˺CwyL(�l����nci:1l�B�`��m�&%B�s���sC�$��,j{����WH��*dM�}q̖͝�~f!���>w�/r�NVCs�	�9=�ć�����i�4��Mdє����A7�
����B GSq������`��(�7�����G��D�~��Y�S#�4T�@���I/J��N�{.��L���x^�O�c��D7J��N��!�O@q�)���#��	8����9���=�(�*1SrQ�"��4Y�V��Ȣ��Ϟ�
��������d�aa���T�p�+6 ���W�+2p�Rɛe�&���w�A�U`�%l�D ���o�KO?��9y���B�Ϝ�xu\�Z�W�5�i,w8��ݰҞ�P[Ӕ�-Ѓ�01�M{�M�f
��bYg�O��1A����ު;h�WA�	�=�]��\�gUU�P��~Z*~w����Z�@��zS	�H})��Nub
4��t����ڰXP��1��-zF*��A.�P��!���9���L)2U��'g\��_w�#B��m�g1࡜�m�ޭ���{,]���>�ꭰK��!ի��qX�Fe\$s1���2HnƏ���^)�ES ���'ظ N�qxx.X��z=��D͑�F���M�fl�j�I	?]�zU�,�V���{���w��G*��Ta������S1@)\}A�dQS"8bQ��WO�N�n��xOa�@�V7���Yk���d�{��B������O���!!�2�F	=�o��e�a2jļ.ߴ�>��`�u&�w������ �ƐfA��)u�R�#�q�E�Tv�8�T׌�USq������3쿛;�M3��_5p���~����:Z�x
���`NM��2�V�E�B9C��������1�����q�F�پ6&��9���H(�������3����݌J��3GD�1
��} �6xf�Z��5s����Df�q����iT��V��]��?P��7��������UW����Iq�b<3�j��\zF��)���ܤ� ���w��f��	���$:��l-2s�Q�j��zy�Io!����Qx��i����M��=���ӟ�{��Sj"Zb�Q;�-e�qXVm����kT���q�DD`��֯[�ˈ�Ǣw5��8�m Cb�g<"s��/�0M��xl�p�I��Js�L['>��'�D��>��`|���Lvgk���[�fJt�1_<��ߔ=�l�E\3(��6���#�;r�B �@�Eɷ��;��VM�(�5���B��a�jڵ��V]}'��񌱧[voB1(��U�B�����}��8�Ui3�Wʅ�&L�-*z�G>R���u>�I�4j�۲vTeC�D8�$���1��0])�l$��b��7��J�	�>Nele��br7M����-��e�v%J��;6��q�I�6F����h�p4��Ϳ�ꝲ��ţҟ�6�.n|O���
�v��I���Tp<��Tde�
�9B�ߢ������E9p"��7������dp��~� u��o,Z.P��5y��qm�b�J�C�pf��I�ӧ3��.y��b���+\��8�����F��]���]6�����u��t/��i={m��!���b{�}��,P���B�N�0�),c�Wtj:7b�~4��Z�z�S��{��?`W�Mh�N{3oc{��V�I$c�_a�߆�K�`�l��J$��D4�o<�]	h�%�m��=�>F��*���|�y��s�g�D��ꑦ`j���3�4��H,�� c���)�#�	!��h�LQ�ϐ>(� �׌�d2l�k/8����*-g��4|���Q����.�M^�ظ;[�~2����|�T;iq(����a'4p�	��l3�M5;T-��Pa�;ⷖ3«4u�8F�&ZA$/R�s�;!�DC�����4nA'}�?��E��z�s��Kt[�v<�/�[���;��¤w��$7��A�?����
Q*}�e���Љ��ѯ?��Z>h�e_ީ��)��#V�X�کc[��)���	�Ȟ���ѽ4pn�,�6/gU�e����)��|dh�yMO��m�
�g❩�����6�X2J��)]�ZF0����g	qڰ����]Y��t��FT]�]��>��.�� ���A����h��E����Ǩ�kub� �������ٶ�L7AƎ��n�e5������ϭ�$q�eT��('`�����ص6��ӳ�_�4����wG�#{���l��Y��@�Nwզ��҈�@xA'a�|Q�DV���X���v�����j+��D�����kR�>�d��[�'���?M�O���j��P��S�,Nq#d�d�f��U�;��L>G�0\����dy0����v�Tķ����-R;(w��.��vF�#�tpm?�ڇ���צ2�lp3v,X��)�W���� 
ɵq��	� ��H쳞U-��7��תī��oT�D��������cO-��4���E��29՗�{�8^8 �J��~j�!�â��'s�{ [�i4�g�!���]��{ ��JI�䯹�Z�}�~���_��)�nR
i\�g�2%�IJ�������I�;��g���=s�8o~�b��Ǳ�c��:�*@�o�̵:�B�l�	�Sk5��Fgm���3�Q�J��������nC�ŏٯU��N��L�BtEI����S��Ɵ�K/ܨ���m�X��R5��x"�:���fS7�8���lhН��L�:l<�W�j�dR7����ָņ&g��"��)�|BsQ��@�$Ns�W���>g�����AK����;�:<�V��q��1S�z�a~V��v?Iz�<s�VC�NG��Jj�ԗ�f\�V��-z���e=GXiW�2IlrU�b�Г��QE-�	�j�ʌ[����ld�Ǟ/�-,�W"�o,[H���*����A�r@���B~����;����/��+?v��0gw��d�kb癏I�E�`R�FZ���O��,Ә�/�%�ؑR!θ�N��0����J��͗�x{�Kٙ����2�N���J�چ�0��Q_�p\��Gt�3l�����q�Lo��T4\���#^"Q_cr�x����`t���U�m��v�@̀�s�г	��<f,V�.�]��R<P�p�rs�1��������!�8!��.��d��X��ču>E��T&1�hC�sk�G�e¦":��2
��.(Q��"2���	��D���^�q���Po��ھĵq����~�����&��c�J�,	Ъ���֯ATU%\5�t$���h˾?��~Ӣ1�+��7LLU7�;��&��p1Y�Fх�K��M�w	���:�΂ES��(�B�y�x����H�$���y�v��y�b'��"yT�߭���`�d5g��"3�p�B[]f:�{k�15�]�2e�a��E!���E�|ntP�U$.Xv��N�;�����9H��*��~�,-�x�Ԉ�Ax��^/Z�������k7� ��E�Tp�@ 2��74�]��K�{�+����Ֆ�*!,z]��􉎅���ō�aiIH��������F�ՠ8%�X<�飭�h8�J��[�����5��x��r���
t�f�����9b����X&���!|ȕ����wn ��V���-���\�"��wshGk�L�#x�7�~�4��k;^<;��L��<����G��p vͳdSod��Z�	U��"9���P�ᏭO5�ys\k���T�h�5�௢����ȫ�ʋ~�+��R���9�B���������5qr��Ns�����sT����@ªx/;N,���kog,
74�Դ�Z���:0}.<�BJ`�`�C�O�/6\Z[�Xb��h��׽R�]��Y�ժܪ
b�E,���i� �[�d���wb8r��0���݉�&Y�z:�+9VB��o��I��+�6ۛ3��M��r�/���i��x�3�� ���gKg�_j���R�K2�W���� CYM�����:�XD ����:��b4Ż펒��S�
�����%��F��؄c�6'���<�N�r�L��7ߢNҖY��*��'	��s:pX\����J��4١ʚ��U�.{uvR�F�[+S���=S��`]l����z�(�oލvF_�t�o��ܛɆ� 2A�r7<���3�@-��'ܟ����Y��;��,H_L��g��ܱ���έ9�y��2�;^'���T0���O���鬻��D�x�B1,�fD��7����2� m���ښXpbɸ~�qU6�����_~��X�
`�%�Qj��6h��[��DX:�)Km�k8�>��.�y�*M� ��r�M�!.N��Ǫ�b)�v�K��4
�!�����l#�\*�դN�
����ԭfB�W�wk1���#��2 ���� L]�IUf����-c�f
��׫k>�>LG¥\����h�'��~F�2��k\L��L��<E�^E���uUi�γ�ন�H��śdάJ/����U��a7�qo�c��b�$<��a�)����8<����e'���\�<n�m�N��k
�����@~y!J{�;Q|,��\���>Z=d�R�\)��/��Nn�I7��mĂ��yK���RCX�o�ʼӟ.P�=��N��R���vt)u~����~;�ч=Z����j$)���n���J���0�|�@���$=��� S�������B�����+�_, _(w��w�R���xoq��ʕZ=��.��ǔx�3�b6u���_ay�7��7�B�Xͤ~&���"���qyT�&b���U��Z��օx%?�"�u��u*X3���� `�V�4��)2�R��[(�V��f�	��`9�t�V8<ڸ(B%�<h������v��-5��^&��4�?�=��x�I���bSE���
g��8H�s���C0����7�D�	B/��lxRg!v��U�W�?ў�
�m�omꌱ��)y���K������m��
��6�dRR���c���i]��߮�e+]\S���(���g^`��������?����Yw[�
�|��]���jga��úm�Iv�M�hk��Q�!�D`n]s�?_Ϟ2��'�,�&Y?�(�|6|�HlޘL��r�0tU��)�
����>���z\I�>������[b�i$.��*�������Pt������5��^�=�d�i�~qt�����<�W���Wf��}�=r%
J��.5�)e,@w�E4�Kp�=��Bm�Өٞ6�_�$c`3�赫�;c��.4ݑ������ORxW��ɨ\ȏM��b�M�1�Cʶ���~y8G��H�%?����ۭr�X��+����j#��������H����S��酟H����p�\�n�ݨ��V_��OW� �d�8�B �}��~��5ٖt��
��ko����G���d���J�2ro��8��S�. Kj��2;�bv���L#�-��Q�I=�(Fv�Z�E��/cmXߚ�}Zy�]k$�^z���خ(U����q�݄�(Fϋ�&d=m>ܙ7�:@]��H���c���wU/ʁ/���8��W1���K^������,����>A� ��Ǚ,���~�`M��ȱ���ֽ��S¾p��V/j0S?k����r�9uޑ(A8���J�ӛ_Q������	���?{�`b��ڔj}��r��j,ҟ	6�O��"�y�| �\	�lE�wU%D��I0w������ƔY�n�Q��=��
l����V�\�#c����(K��T-u
�u`U��~��۹΅�%��@`���aJ��[Q�wO{�+��a,z'T�ª(J��3�L �S~h����doU
Z������f�1h��olƺ>��)���%��a�rY���:<�Hy�a�V�Ѫ��	5��dS��)#�`K���A�D/R�m2���t]cqo12+������uD��Z��i��s�F+�A"{���4V.
\�� �Nh?��VVzJ�*��T�m�r� ~�]�����g�f�PgH}D6e�TG>���}��a:'Ӻt{��S��kr,���Po�%�< ^�~��,���
]���>>G�U���S���v��6�;�Gᜅ��t2���	�j�^Z"Sy/�� <�k���eɵ�9�����c	�@�ɏ_\E����\�{���裺�jmwE�_q���X|�t*��2�sy��L�(��d�Ljܺ;��{#Ʀ�,@�;�Q|�sa�t�5ƗF0��
`��c��VA�iZ��R-i(�7V�\�L�[�x�ݠ#�ȵ���0���j���>�Ӆ���n ]y�)�U_%�#�t�B쟵+�3�� \�R�(��
h/�|�a��e�Н|�쁱�g�.�aܪbIA7�[a/��2�Kh���oE�L��	�H�IMgl�L�����?hr,O���� ��g\�
ގ����b�KPߍ�;`u����T/�_����8�.�Ҭy���&Dπ�.#:P�s���/`KZ�k�^��7���dY�y�# <�͡���hH�Xo&LZ����:��t��?�.���>�eV�T8P���/�e���uR.4A� '�-Ki�z���P@#n�q`D�:�gv�m����*��B.� V�k��C���Jo���s`7�� �A�L�x�?H��6���t�0 ='�w,��KXM�����2C�DK,�~�q��j�
�^�F�Sx�Ig�N�>12r��٠\��oޱBc����jg���.Rzj��ddu����c#@,�	e�[k#d��}Yo�W%��s�p(��0��X��)��W4 ���a�W[�+Q�+e��<��Ӷr�[ϑ!�ӵ�>-�^�Ü�ȁ�n�
F�,��QXJ�������@��T1`�n��-[y���8���C�<��P�n�Q�o-:��&"�K�g��0J��]����uc(�R�暠ͣ}�҈�`m�53�#J G�B��xu��X�K#(Z��^��ax��w,�k���%D���*�F'�~�5�Ɯ�m�@��W V�"K[�=T潕$F����6U���f�8<��hї \[w�=��d��&��[��D�j���+�~��[�r���ƙ����N�l�T��:��g��k?L�9*W>r�?��7��N�J�d���W�?ո�E�{Avq��zGwv,�p�.��K�L}�rT˄kx�|����6����Z��������!�Uv�]ҷ�1�E(8ˁ�z�R�/�����h���`@W�>�;- �2w���w����ۼ�t�9|5�}�y�D���d�;SW�kgd�R�e��� �a�۔ՙ����[����4�{9�4�E�[VSc	ä�����m��L�g�M�v�nϦN,�M�'�r������6����C6#�7	aI,�y=Nҋ��������MM(N"���R�D�ģ�rc�����ۆ��R7bI���[�Xqdq}��>�i�~�<bP�Y�$�s��"��V��HoC�Y䞸6)3�w�OC��p.�KDN�Tx��
K:� qX�FH��������(#���E�Y�_��E�W�����<��-UFmX�#U��D���ۜ,.2}Op�=�6�q� �x���5%��r%	.�k��lyJ�ݺ�œ��fK�Z��7���d�ƦZE���[+���zM���l��˼[t��#w��B��vNRs�hP��"T�<<�{Ɖ��mח���e��X�[�I�.�c�>�i��%@����	�V]ƩD�����QkBWb>���-�b����#�J~��8��(m�|��1�_����B^q�����h��+t�����/^��!U�	$AQ��N3��u?��?��X�[[=&c��{�/'a͠��>t;g`��)���nR3�{3:��;�Rr��z��;0�z�t��01����*z��e���uG	)@ho�d�G�,!�h�DG$ٟ�@��B5:����-��y��Fη�Q�q�ȅgns���_�$�^qGno��C�^���6����z'F'�/¸�6�il�
(�w*�Y1��)�d��l8"�g:�g�{_;$B�9�Ѓ�PA����E�z? �D_�}m�k���_���G��&��h���/�w�4)�q=���uXd�u)�����̕�B^nEitSs-��e��4�Ib4���E5��F�5�$��x��4^l��.��T��2����_��!zh�※a��¡��iW�MľƼ��G �b�Kk����/_��w!�n�{�(��A��(q�9����M������)р����� ]�;��\+��[���,�W�1B�v�Ȝ��%��#��U@�3�C��2D7��:m�(�
sƑb�b���|�(�M��L���Td�&ظC��]��I'��!��r�S����%�$��j� <K+a��Γ	�c��ç>I�G0�=5mF�-2B� >�Ou�W�#^OQP����G�a>��/��Ҵ6�쓗J����{�����n��ax�(�lu�d�Gh�'.�����A�.99�,��Fժ�<1]�������t}����p��`�XMFϯ ��~��PŔ��8�r+8��s/gO�C?��CCH��<wT�QL���/��M�g��݊��D�E2����B$#�_���8A�o�7�Vܻ5BWM��\�Q��^��dn����_�7�ߴ^n<���|��]�j�z�F����i��"8F������n_b���z1�����hmf
���!v�ݠ�i/��1�b�{'�`��7M$�}Vr"��rb�Q8U )��R$�����E`	��k���8� j�fե�.
�`^p��
����"�D� v{����qZY���"&�B�*����aP�v˪{#�pr�]P��ǚ۠�TZ0�_$iI��|0�_������$7	!cW� v4�_���-�C��y�9�Ogd��W��x0��d�?s��6�u�4|A�w�+0bs��`����)1�8�nL���:R}�d]�@o!�f��ӈ�旘� ϕǅv��E3��F�W����U�UH����D��s;�y/��04��v��Z ��g	�ۣ!��(Ex,��O�d��]?�E�2���]��)�e��10��,��]�	pX�m���,i��;�P�"4���p[7�!Y�0\1��দ���m�9_{tA���v��47\��N�gk>��<�BL!����Y�����2:�͉`��;�Lw�n�u-����e�����q�5�Wc9=r}y�`��|�ۗ�P��^��a�D������0�b�tnz��F�(l��T^�o��X6��X%\���KAy���ݥq<��6x���ت��JSkGv�x�lV�`�y�x(����F�qqR�t�U�Y�4@S(t�Z����JQ��pA�Ӭ���ڸ��p\���Gn����j�.��A�fR���ދ��||\ȫ��E�wa�7���-��0\�!��S�%J�|��h��� �R�_:3��cXX7���ꭧqT�T�a�h�+>"Â���cA���� �hu�Z�5C��Rh�����<���r�$�Gc��w*�.P���o&/�����I5e'�l��FB���b;��J�N�z��w0ݣ��QZ�BTq���}ZD~u�x�a��
����_��~J��M?�7Ǉ��%�q��*�L��@�=Se�dBW�A��R7�fOǠ$d�妢[�,څ4{�����v��`��(���K"�x�C�헄?�p��F����p�'Ĕe�����
�DUʢ�p���[S*b�m��� �Hε!��P��˩h!�g���e�����9²��o�i�JmMl�3��j �T�?��|���:������B���p)�w��E$~l��M�_�ae�%Fψ|_Y��5p�s�Q֧!�[3�2i	`U>^��Z� ����J��?d�(zni:�3z�����{�m8nC)͠VBO�y��)�v2�;�I����fh@H"A���Ca겂�ܞ��fZqW1bg]��`����܈�?6t��`�OhYl֫:k�6k�QX�5�)%J<%�]�#_X���Z�c�J��")����?��uM6�i�
o;2�mz�4�V��HztJ�h#"�/ߓ��Ht�ށr����~<3�m�(~����և�Ki���Q;Q�?�ʖ+��W5��݊��������L�[���<�[Za�=T�)]�Q���:R��h�Vlw�*�8ߛ?�qC;EƵK�L�[��-��'� &��ج��9j�E����P�q���-E�O��V����׷�YP����򃔪?�
�aH�$�������s��q�~y����d�s����'�����K^M@f�ݟ�HF��.FY��V"��e^�����D.��y�7�e���I�Y���[G1��|����.H0F�#d���9�v��:�}"a��b�LQ4ʠPm�w��R�(�� ��J�v�K�3Rz�`R��-�L��	P�6K�"��u!�#�o2p�G�(�&ь	�r֐��є�
����O6l��[z��"��7��@��R��{�Bn�hY�V
�� ��.Ex4e������ �I�.Jك	�{�ӑ��X�e+|�OS�:xxh�y�\�	�b�]HK��¾����c��6)�z�g<�&�E]��,���sex&�U�ot���#�̖�;j᎟�íx�ӂ;k����!�Mp���/�hѠ���t��/sމ�z-�����R�Q\4o�d�Ez��/�-���W)-Q�5B'�,�(�$�Q���-1�L�B�_��"U�V?�r�WQr�:�AD�b[RI���|���a蚋o�~����h�G�-8"|Q�ug�FH�����G����Ў���Z�4��dprƭA;�'��jWv�FY����5��vt�uo�mf�d�;��BW��t��[�o6%)3e7��ꁴ�c�ޔ }�<w!~y�{BK�'�T&�n����\�F��a�vO�gp�����N�l=Uܐn�ͪ��'v1P��r��]Cq즴`:���ˍ�疮]����W��u.jFs�r[n�MB�� @[E�b�ԓ(}5ʹ�� a�6㉶���F� �بĒY5[{��.O��W�]Ӄ���҅5�#p�qw�|��F�XE��P	��=�m�?%���q��l�c��󼂘n������*��;y�RЮk�_����Q�ދw76�#D��̽��K@}�Î�\�?�%ί���I|�U0���1��6�?����Ǭ�[-5�ه�b@�^�q0���H���D��Tf�9t�X�繢3��˺�l�S������F*^�g�>�V����7�G���6�=�����~��""N�x�
�G�3㪏inD�J�Ԯ���\u=���)�H*�����W| B"�k`�um	=��`�4%!m�ɨ���"l�5��a#T�?�a�����i!���g~����amQ�3��ZaGk&��}�>Ұ�H�պ^��J_��@�A�B����@�hC2�rFI �YO}�~7D��x�Y�Sk�J d�%�A�d�O{�~�4Ĵv�^����E��JH'V$�Z�{V�(�ִt+�N`v�g2�h�:+�=��E��;С�.ގ��5ǳ|T��#Q�%z<�������'�յdM�!ǭ�ߜ���/� ��%�0~=\)ht af���<R��D^1�����D�������L\;�Y�Û�B��d(�B�_�����3��0)s�f�c����>�d��$�\�@�a5o}:JŜ~z�O_p�!�j�J���c�wL�6>_Ӡ��{}[�gM�jL=�۴G�P��ɡ��_|fߓʘi�H��f�1�͠�#��{W�Rƌ8#R'�`�V��P_��#X���s�@->f[5��6��LP��F��}4�H����fx%Y5�bi����E�E�K���B����ɰ0b�%���~����v�[�8,{S,�~
E�NcjE�U`y:囁�K	�9�ǆB��[�=�����6���Z�u@k�Z>�|��9���('���j�[J�j+�2qP]��r��^;�2�r�u�S8��z�z�):��g_��,�Re[���]k�'Ǫ+Ff�������&�����1���ү1�0<d`M<�F���j[�HQ��%�O�$�*<y*W=�>S	�s��x�LG���)O�������^�dX��E�tQ��Ő�-˄�V�h�L���R�q ��V�JS!���WH��&�B��|�`h����S}�zX�b�ǙZ�]�$���K{�������ވ"��=�W��>��}o���Ĭ���x�ߦ1�!RsW�=X�E�y�%OH�x������^{��]��L��:�-��]_��^[�l#���3�{��������$
���^�h.V8Z��U7F��@�ߍ���R�ϧ|:g8������9�?ʭZ��-E:��a�C���2��z��p+T����z���p/�"�u�����]>�:�G{��b��v��o�x��9R,�Q,Dew�W����x_�1Y��8sB��`�C{���g�<7��m���R48�=��W��C�s��H(�u�gI]��\e=��Ce��*�<��^��&����VȀ�tr[MEWkk(#�e��Y{u��%�,�Cz����P��.���#����{��;�12�䜶�=�����N�b�,���*����P,0�s��R	��<3��������_��髉������j�^���/���4�Q�1]�It����$:Jv�S){��!��[1;C9m\&�#F���QԛHN8	��L����[�Аr�]G�
��s��?}��Ӡϰ��`NX]��%x?H��}�h�����p/մ���+��/o��=[Y��j<��cL$.�ͭm�����"���Yet���7�k"����L�8G�'��2G?����z�-�7������=��F�?�����1�]<��Xy��}VX����7Q$�#Z�����^һ��a.������dK�f��:���TQ�Ώ�D^ ^�s��,leuc�n,o��=��E\�p�R��xU�^[{~V�����,���gb�*�X��ҩ�SilA�O�{J3�����/�6���a{�`(�s�o~;Z4�|I�P�M�ٓ�����a�$��U���& �=�6a0_��+_�WVz�OT!��꠩Ux�Y�]	ئX�n���Qb�Ǥo\�}Y���i!
c�����{3�`V�Ռ��ݔ��܆Xq���g��������rw��t�r���p�ѥ��>в�W++h~�0�H����q�x9�D�%�VBD�t�(y���l����s$��\ o�P*�MhQjL̙v���"e����	5�O��Z�T�����R�1gB��z��hRC�ۛ�di�%�f5���g���� U�����j�-��>mδ�	��Gc_�胎Ҧ��eo�2���D���[u��J��`�d*Z���ط�άl�!<[rb�8pm�2l���N�u%{Cq�ʌ��U�7w�D܌Ҟr�{�=�KX<�T��
�z 1pAı��Zñq��7���N��u:�����ֽ2���8KwȎ+��5x;��k,�� b����s� ��P��/��p��V#>�4i�����c�� O�;4PwEJ<�r�M<�A��8�)��DkF�ܭ/Q����W �sٯ�*�С�>���?�<�����2�o2�O��F�'N>z_ҩ'�w}YL>f,��o�n����b2Q�K>�(l��Z)\[L\��i��t�Ґ�Q�uR��H Ϥ~�g��YtHA,C�󀊨|�v�f���4��wL���'C���*�E�04�R�y�����L�2�x��ѥ?'s"t���	�!Mv�\����.�5��Z�8[�9�Y�T�4�eޥJ�m�@�0�x˜e󎠎8��S��/%2�-J�khgx��{yQ�ҝ��������-���Ħ`�&�D�E[y:89Z߮����nr�U޿_�R��|L@�C�sբ&_�.�!�Ǟ`Ib�W˝ hB[z��Fkًx(�X����ysqR꧉H�ߐ����\5��I���8�)0�2*�ٿ����qikʾ��6�\0^ �Bì��m��q�]�D�96G���p��O�͡M����"ҧ1��͐W���"�.�t�T�*U�`����=�!�6�+yK���u��'1@)��Uc=A��\��I� �u�P:'NH�#���3�����ꙛ(�c�
k��h9�&�L��k却7��pH0���5�[������n}g!��b���}�.}��g`�+6W>X�n�2�MR�����\�����)I�����p�W2LU�0f��-����0����:�m��&FK���5��Hذ��t�&���Z�B�,q{�B�m�2>�<�;s>���S����Z���.~�}f�k"O&���\��6ͳ5@�gS-�~A9�q���1�2d%��K�I�q��B�C�u�(�V�O�y����l�M�(+~�v�zO� �ۅ���]�;�j��	�k�.��6v��Ί%��r$%�!�O�v�l��I��ɐAW�o��.Ιר���)���j��s�h�6��
]@�8�`��RQC�].���8�#x�jZp'_g?��� �\FjŃ�<�P���n�"�Bm784��k1l���-����^A�q�_�iy��:v���=��Ub9���BU<dy�7y�E|�ޚDgH����2�#҃��mŅ4]��歊M!�� C�jd�j"D-�$��n��۷��j�'��<�B��1��<��<��>��0f[#�މ���"��]&��]%��a��b_��);��m3Zg�Z;�NΐЊ%��L��w��!��
J�/���Sk����QVQ�r�LGIj0L��'W�z-m,S���T{g��D��g�=����t��ѩ}C�j2(�$�oi��9r�h��s|)��j]j_u� $��#W�������>e�M���k��K�m�r�#.�ۥO�*̀�C��т>����vr�k�3b��%��Z�^4T>�@�;�g�S7 n7����'����Ob�3G}2W������Y>-��Ҁi��e�<��<Ƒ��R���ݣu�p���څ�b@��	�i�R^4$��# �Ǩ��RY�D����J0F���_�c�G�����@�4�s �����庥��MY#K������X�V|����:��w����2���C�}sG��y�\�"�H�X���B:̐Un��T�+S��!�9.�:��)|�e�foSf�<,�/�H�T���<�/���?4o���W{t���H��tڬ��4%x�`�.5�� �[��ԓ�A�@�u�,�,�YՔ�p�aj".�g��a���f��\X,��&�q�'���A����B�<� �~5|E[s�a�Bi|3]\7?#�}����,�Y|���0J���� 	N��̷f�ڒ�a����gL�2�Jإ��$dcj��41?)W�Y�yYPr`�W�'\l�5h-�Eq_����C����w�r�3
DF�:�C��ْw����n�+�6k��Y��&�o�h���VQðħ��O�����\�߬��pL�]�I	� h�`�k������U:s0ؖ�"Y2�����?G�ƞ.�n������W66lTi�S|��;8��؜�&<Y�.��i`�ҥ��g����d3�y����#t� ���u�_�[�getʌT������=8�*�v�oY�ҼC-ۈ�O�{�!��~�R�������+�GϋJ�D����`�g ���g7Y	��}<%U
H���1@�m�WK��5�fUҕF3�3a���?O�bn�Z UT2�c��@2�`�$���lO�S��Ty�7Ug��~�&��	X[X*�MsW��Ok7�����Yp�m�Y��m�iAZm�+�i�I�VE��u$�l��&���^h��ZQ���ϖ�����Ї놆�&�Ӷ�-Y2�U�?�*22<�Nɭ3Ւ�c�1�_�P���]��<,���Ai�ҷG��.�t��.'3��pc�Pm{��H?s`@��9�
�ë�~��n'����r+(��+��b��F�����㔯�GH@�wCj6ǖ��vݴ1W�Q�q �� �	k�0��P�!���t����*ج�eIZ���$PƼf���&�م�)���u��WG����j�N!��:�&kڡ�Ȅ����a8��u;��}��������MnW�V�5Q��ԣTN�}��5ו}�Th��!:w��d81�=��_机 � ��0��v��k��\���������l�zQW~^���y���� %:�A��$3���7�b̭���hCK��q�
�[�mw�}g!x�����������`D�g�;�/�\�5z�/�R���������09�A��ZF�5�kN�ȟ��W��5����@���yF
�jDFy��R ��M|��_#�Q�i��B�|���!Ѽ��vOԅn<�M��F�	֤��EB�#p������ľY��(O���tX����\I��=�k"N��V�˜8��4����2�^��1��W* ]�=֘`�=t	�B�=�J�K�Qa�j�S���(�P�*z�D�t	��z�Jq5]ѳ.�&���� �eef�������������f��{|��`�d��p��B��RhW����yD�-�#
�m��r�w��u�tC�����޽mW$6��p��-���u��Fo`
}���s6�[�n���kU�o�([�d2>8Zlе#S��� ���y���-�M%�,gv5w�E��tAz}�D��H`О���ݟ�ەe�0�@8&��]n�'h���澃���k��w��a���.4%u
&��LӤ�cTA	�ۀ;�t�
�#��ֽYwo<� �B1��";�#JT-��8�.+k]Q�}�B<�M�5��*���^W�B�tC�G�m�q��8��(����%}$_�I��Cʊh�H�@7��UT��x"&�q���{��D��(@$/�0��LuE���:c��)J����A�Ȏs<�L�,U����-�Hl�>����T��+�!��K�r�����P3)�9$�y�-�����	���M��֛�&�����
�K�,�yJA��/*�4g4ni����?3Y�P<�!D��8R���>��O��EƎ��~���kH�Nn@}��al<��'43�f~e�Ej��g~��m�vg3��Ti�*��J���
gN�u�����t<^0|xu���"�Cp�&���S�G�D����T����q\? }ff_����s*��"O޶�䳵�2j=O�/p˔G�Mٌ���'i�&�p���Rf@F���>���������>�>^�e��|7�N�!��6�8�0�FXyK��QjV�D[�6t��|�;���,g�h⒎��v!K�vi[�d��dR�?��U�^�a���k`(��x���ݶA-M�c�`�"���b��oJh�d�����i�����ͬ䣆6Y�l�'��(���6��/
%�/o��|-j� 	q�~��M7�_K#!���Z�������9<�6z�,�3��Vp�3�E;U���^H���~�!�h�%��6�-�P)�n�*�E�M�|/����v����v��J��`l0(�_�\��$J��1���V�\��
J���|��F1��ҽ�u�8��]6�K�;� ��9��%nG*��t�b���]N�*D�=��چ�R�-��.����6�Ei�Jl��X� Q�qs&Cf8a����?��T+����F�g%8�Hu�(�`�ρ2�Jl>�x�5�x����QEbF���~�x�[~��,��ĸ���'��s�[�w�U��Q� <� ]y@�qoܒeE�˔�z]�O��d`j@��̶Ku��K������-�R�-����ϳOɟa1&(��x��[�;�1?� )��ӵ�n�����Hv ��,�qN/���y����Oa+o�oR�r�h���U��%�Xm%ύ�bV0��
T-s�m�	5�{���t�m�Cf،��iC1�*ˇ�%���5ˎIz���#=7�)��f+�-Ԓb=�K�n@5	��!��y0�Gt�	B2 ��LEb���o�[��WS���xʐ{Խ+��v�i=r��G���c�#�w��K��)�2Z�p�M&��9~��W�p���|��0=D$���f����g��OG|+����k��]�d�wR���o4��D�iSl�چu�F�����Ȅ�ߣ�E�)CC��vg���F�t,Z˃�t�{��VMjEN�?m�ت�$u�E�Xp�f������j��3]N��<\z��@	�M:Qϕd0�S����wg�'XxHq��>�s�"�_m�f-�����̣ɏvX��KJ�W��a8<��Ս���
1��ʑ��3Qy{���F݀% �g��^�5yH�"&��)S� -ϳ�V̛�.є��㗊�`�?����}�djhH������ɔW�v�'�]�E~$��)
\��!�*�; ���n]�
p�z��L9�n��]V���k?]g����,�c���7>XU�b{a��@?�m�aO��p�fps�Eܢ�"!x��r���u�>�eoip����-`�Ղ������e]*SL|��|D2����_��7����4����|[v���SkZ��%5O�M�]I�XÂ+���F:�-5aC �C�0%pD�fi��A	ե�)�+;1a�IDp)aP�t�����|����H"r��I��eC���G2ә����uc��?w�z��#B�&�&��G�U��x:���MC��$_�h�)km/��]�`�D��OC�Ӧ��R��b�`����[�dAj;B$w,�߇��D��[���J�[(��C�Q��Z��P�Uɇ��$჋=�"�n�1�*zҍ�<�k�N*�{+��yx�����*�T 9����RS�=2�"\쌈�t�;�0�8W��'R����-�v�l�6�7�j!��|�]�3�u&����-Ē�7Q��xC6���!Fq��z+���ȱ=t�]��bp����Lh���
S���������B���]\'������6b&��,��O��yj����J��܉Uv�=�0�,x�%���PW[��F3�0���������˯]W���
��� �D�\֕���z��|���͠���&U�~XK����S�qV�.S�.��OJ̤#��Ksp��X��oF3��G�o��XdO��Y?5;;�Uf��yւa'�[Q������18W4R�D�%�墐������w:^,�fn�Z?�ӻ$�ފ,�5e��9#m�D/�Qp���ʆ�6���6�CLi����_9Y��Oo�����K��+2�պ���A�9B�I02pQ?��U{T���_2͈қpS8�K7��b�w�g�\0#��=: 1.���8�����ZF��Ɏ�<��*��ɼ�����G_ۀ�C�la���Y�Iy�[-L,r�@K;Z4#����n�gA���}�"D�&)����r,��g
�2�?�����<k�����0X����Ǥh�2�K�U�0�8��?�i��A�	s6P��A�M�`���n� ��gɛ��4�4���%;d4[�A�(sl�
(rJ"�̢^qQ<Y��x.T��?fM��ϖ���!s���f�쁚�$��IW�qf��^�]j�ߞ�0��Ϧ���v�΢o��_�t���D�M��3���#0fh)�#���NŤ��&8��!����?�`BV3�ey5+��8�����>�R�*>�����غc�(�)G��O=����y󄱼ã^�-:��G�خƴ?%Wj��=d;H��B�گBp)�l�db���aE���\��{�Hw��;���q�c\��5��?�-B�+6ӀE�k�����a~c���x�6f�$�w�c�����R͔�����9|��	�m�"���
U���f�'�sܪ��H� #�HT�kT��05�wh~rZ��G	W���8�%Mʎxm��Hc:x�E�q����%c�U��y6:�pHMv��:�Ȁ�욒v?4��ЮX�V
Zw'kXL���N5�o�k�(��]�d�\�"���o���Ng~�+��b�P�b��bE�6�Kaß�4/��;��\:���={�J��WRq6b�U��ؒ0#&-@]��|�^<�k��2�@��l���zKB�G�Ү��Nۦz��G��'͡��H���$��� *`�$џ��6N���TI8�=N)���S ���yݜu�ߜ�꿠�-"E(��$d�}��:A^�U>P	M����V��L��
�1����HsLH �\���w��"C�N,����Ѫ/�2�
���ŵ?Y�L�5� ���nJ�,gr�%d,���l3Haàm{ǭfOrzaFq��1Em�c�X�� " �i~�"/RTāQ-A�딕7�4ఊ�4���Uxs���0��oD�1���%A����\������/;���?	|̠�������@S����?'�K�ǉ0�'��b��	�Z�Fߐ�����_ha}皐�v�@9]��10��PQ/ϔ�A�������������,�8C_�� :8ʯ�2�>�c3��i��f[�>0��yNpf�On��-�:0�s��������Rq3h�>���c��^.	�B�ts)h��|��5Z���=H���\�8&��+��Kgk�� O�ha��%v�`���mY.:w%�[��Z����	�}���61�|0��yC�"
$�e�N�m�6L�3��V���c����҉��t�C�l������O���p)�3uQ��ά���n�ڪ"����V#��5"�i��6dLo#d�y|����+����Z��L��_�MKHV�(�X<z�����S�QU*��[�����)��C����0��D���beO�m(�`�9���x�1���C=��G�eP�����h0����#R{b��OsH@����Bw%�}-�X~���zL�6b�T�fv�6j� �BK;�H����|;��h*ô��O8��`��%��ri��}��`��Q�Զ�6D����7p��X(�����;��U�8�d ��IhK-g�~�(d�wB�p%]�@
^�@�0�&A+��H'�.1�f&H#/R��#DܙC�U��?.�Dm���{/e�F�l��(�H�k���Ɉ�gbAoAd�& ��rʰ���$��7juv|���VhS�^S�~V�ifD���mM��g�	FC6��:�dp"m3(*նO����HX����Q<~yVbL59d�t�Y�G.��E��V���}�������C�!��?q<x�J��cO*�?�n*�^�.��I�᜻�G���.�
S$X"������vL���-Y�@+lȘGJx�R�H+q��(�^�*�C��?Xt������\��s�wM���=C�M��t�&�t)�@U�/;�p�I<5Ul����d�BYB^�q3���?��������Ŷ%���VoC�7�N�W��C�r��Pj��$e��r�)kĔ�Ҟ�T}��q>���4�S�SC5�k���/�G�>
p,�-e����!��.��Fx~La��~����T���KfP���t���>Y�ë���鼚�xh�~¾�=_�wڊ���1��U�C��($�Z�un����
�$0��&����ʾ!줾c��]D6��^��2`刮;H�y�~�"J")�7y�ԧ$���=��Y�pb[pbG��!_Da�ݴ������u���+1^V��yV���m��g����sD���s����E8����P���%�h�Li/ɝ�oD�U�	&����qil"1~kJ��F�+H�ʖm�2N���i%��0s׃W���ᶟ�o�%����������]JJB[P*N���Y�[��x��u�i�=�_VU����~��g����ۄ6@yg���z���بw
)�s\5t$�Q��B���H�˂d���֑A�ʸL�ˉNa?�YZ��Rp6�V�)�o����	�&^���c�p�S�{��@������V٫�����~~\"������4թ�QR&�� l����8݃Q������-G���j�-�t����M����+D�C�Z����c� 0nh�4��s#�M'/}�A6��� rp�*���czÞ��i!����A"�ݷ~!#���\����c�"������g�$��6����1�dC��ΰ�#sW�	��T���1i��p���ڋ��-���������`�|Y��~�0����X�rL⧀�T)�
�#d�$���YM��v1�b�I�X!]�i�q\'m>dsp�؆ѧ��	�>���%�����6\V~�Ý١��G{FF�jqia��@=C�����!K�F��UԉF3�f%�/F�N��}31-�,���l�A��Λ�����|�8OIe���]��+�Dh服�!�]����e�'-%�<(��LF��t�.�g�p�*e3��)�8��l,��L�;�6FK����*�=̛V���#h՞&E$I��Li[@�]uE�	��8V�K�����U�zmq���ӹ�`j0�H�~ڸՒ�$�^ <S�6�+���C�Eܫ7癫���W⪓�Bu��%o9v4et�V�\e�8�������/#(����6�,-�S��%���4��t�*ȝ��>P�g���,��'�[Y�,Q}�];�0�6J�
�8#_�H��bJHJ���~�ٹ�c��AGCoi�e��٨�}��=��E
s��v�q8eOԲCƪ*P4�'?P7����
�>�?�a���d�\F�C�
�=�C��k^p�����T�RL~�B�,���Z��K��KK(�4v���@�(���um�x6���99W��l�]��~�v0�s��^��L,�7Ͱ��Z£端����|��rze%W�P故����!����5a���_�~�I�)�>ȷҟa�ێȆE	��$�w��-���i�c��N�Lh�ej3W���D(%�kjH9����5���EI"I���n�bB�2=ㄺ@L�j+�����w��ۃM�(��6�f�ԽVg�mhH��7y6&�f�9�e�t>y��>��e6h&� ���#�9n�.��D��/E�FP.;wm<��C�"���N�a����<lH��1��SX)�zl�|�Ta�ALn|�ؿ���B^�	G��n �Rs早���\�K�ca����Eˊ�b�	�4�R�q(.ٻ�w�]�o˞{dX�-	 `V�
@�u\~Hõ�������N}���B��z�xN��[�0�	v�	j��(G��//=t9�[��CQ���P�X�B�N�F��t�1�x�& �}����X�<J�&B��(���?�������Γ�\���ڂ�q��W�h�m�Cb��.��CY�m��,���^�	�!'_�5é�� �Y=���+�S��� �?��ղh�����ѡ��W�lNs�Z=��oC��U��h���U�*�M�5x�E'���KI�2�i3R�n����l�M���`h�
>��
�@]�B��Unm} �%=�4�Tӝ ��i�w�e+���t�Լ!Pd:>]z��wQd���b̟ۋaۗ��يĺ�A)7��ᎁ=�v5��o�!����V�<�K,{Rv���?�MʤD_��:���ˈI#nBU��R���|^�#o�s_���1Qo���H���gY��.����J5��)?���9M�C��:�n2��3n��) ���C�pK���$OS�bo�B���ա�r˞l��fO,@��lo;i�2���h�O��Lu3P��=��9l��q�`C=]�:�k��X���*�I��c�4���:7�;GeKnr���`s����1���ߜ����I�Y3�݂��S���(g\h~6_�+��c0���6�@c�\��j�h�(U`!�	�=��#*w�Y-nv7j$��\*��M
j�Q�C�x�f��ɖ�K� ���[Q׌r2'�R?��ѢPֵu�ٶ1!�����_*��f��������+p�J�UOA)E���Ŝ=Rc����}[pc��
����1�w�w�^����GZ,�1���R����[[�/�3(�b-XTd���R�:ȡ@ɽ�w8�Ӥ�yb �S����5�~
�w�#|Nچ�5[��	��T��m �3 ��<�/�3�c�����e2��8�7��q�I�f��e�(k�`9k#�2X�1g�Q�Z��l�V"U!�M#3�@�܌ c�}�7���	Y6���r,�S��)붽��k��gib��]����w�U�C5��JX�2�٨�g��e��0_ �yo ,��|�Bl�au:��^e�z,�����I3�ףt�M@�W(Q����.d��g8��$�X��on�M��%am��U�"���a� ���b��E�Y;��3	�=?�~�2�Kl����jB��-�t2S9l��F�߯�LX]�8�w�s�Ӓ؉��_Y�o~�s�P��� e��d��c�)A��2�!0�4�	A��]!��?ˬ.���%�6�i�J3�iYY����YW�۳�vR�`���&�Qj��j�26�[����+�&��G��3������i�����Ʈj��4,J��VK��\�M"�q��_O�33c�k:'=ɚ��vn��n�T.�t��Ã�ǔYX�� ���=�99V)-�gm��c�H&��U�h_�AS��D+�ws��9���%An�d/ͼNp��i΄6m��C^�3ܲ��af���0$�UCS����u�!���� �H�����L������_����$�S����v�w���)�8J�}��鞊�< +��Œ��I�,��L��n��Av9/+�pS]�!;��M�Y?���$BϑbF��C�GN�B_NT1�a.'�5n,��Ek�8t*FVm���kv�7u�UK��}�42 �\r��,�̱����:l�Bȶ^���0$uy�Lǆ䨿�]Vz�@�}�6�3[����Lڙ�E�19?�r;�Nav��6(��p��\� �Q�.S*�:?����՟�UNHJ�w~�]�M�#ߥ�����E�2r=۝���ݛxi$�!+P?�4�&�>M�u8E�
�#V"e�-�l)�T�S����:>��F��~����S�S���$w��h�����A4ڄ�~M�	�	�߾BzV��ݖ�	]/}�`���I<���f��ԝz6U���\��(�0�ۅ..�}ǡ�uz¯A��Y�M�TC�\�W3���Xlp+á��2�G"7{�hɼA��]����t�OKr�}��h�Ve���G��<�Ւ�U��fĜ��V$vK�/H���&��t#��pܱx�`���! �$.�#����򌜱�lr��]Z����"Oa_�*�c��
[�����C�B�jG�0���тo7x�
�$��cD��V̡U �_�W�a�	�!1�z�'�dkYTݲag|ze�����G}��]yOc�w���!��1Ņ�~�ОVB7/�/������Ax5��P�(Vs횢���FS��ݚUR`��0�j/��Z�˔��	�����фUr����43���G$4ƅ�ih��,����X;#?\.vE�eW<�F���Y��(�I���l�m���?}o�o.�!-��Y�����9��p�ʨ�����l��_M/ҏ��B�M�)m�Eʥ�0�)*^�����X��D��ȼ`ʆf��T��=�`T�}cFч��V<)q���NVi�}(]X�t#B
�l�Hn�yY0�-f/O��L�Rޮ��8"�'�Y��L�g���
�B��ހ"�[X~Tw��rn�$�z 1��� 쏟Vٵ!p���C|7�������*�	�q�f׺�Ͽ��o)�)q��W2�^�e B(E���������
���H�XE�Nw|$���R�H����׋�\�*\/���)��Y�m;�қx���]� �!@H��)��*�`�V���6\��^EH���ٿm? YP�(Sa<t��OM��bln;�T�O�3A��AG�-�W2m��ͥ`���/#(�A�ۢ��$&7�S�! �l�:O{��Wx<�{U�,�V���`�{�L�~q��Qt�ϑ�u�"l�������a�Q{���-��A�(WW��w/��a�8�v��_HE&<�ŀ���F	 ���8zC}����1�9J�w�T�3e6�u�{����xm[)��k����Wr���U�.-T[� � �������ťє��	8f�m򰡚�<`�,��*dg����� ��3$A�D��sk���NC�Wv!-ua�lB�ZEAE)��qnW��1g���b�ñ�ץ�_��d�OLD�9����#xb���gg�#q�}�Al-P�Ζ���,&��qۋ���0��K��爚��%��#1RU'�|t\�+|�,~�jkT+D������GDNx��̋#t_�]~-9���ه�>�L�7�����B�(?�SF�6���ѓIB��@��UA��R�lx���Q<��A�4�|��W��id�R���&J��3���w9���j(#�A���� ���e�VF_9T�Cȏ�ϝXր,+��!QT��s��FF�ֺ�ǯ��9a��3��߹r���n�[�$�iCև(���@3'C������fdʻZ����0�Ov��#hUn��!��R��x�LW`uA�qNE��*�f�ҡL����	Ol6H����;�	�L��������C<R3]�����`�=ð:�h�P��&➟6�}��ә#�3%�IZ�
\�B�9���L����a��"l�J��}߫T�9��	����wƋ�ū�}wwI���fq>ӆ�:��5�q�c1�Df���`1�`VH��H�l�Hһ��R�`��Y%�䪶0�R
�N ������3�I�h�_P(�3�y4LVg:58�]ţ޸����γ(c�ܛTcs1HM�W<F`�k�N� ��$��!r�aB�?+��2�����	1��������EzTrs��N6az�K�g�LO��ª�pgl����b{�[g�Ӟ`�݆Y��=��zco�������Ϧb�򊩜2�an���9�R�7��e�?�����}c/u���76���m��|�ۮ�����M���t'C�GuLo,;�����%�I4L~���e�b�,�Ia�1SB�F�ⓔge�r� ̞���$�l͘� Ki�lȇ���&�ѲV���幪tqU*x7�[J�رSsJǻ�g� �J���΅�V�F�ïL}��3ERE��S�v���H�g��q���{��q�B(J���؎_�S"_��E�o`x_4}�!�j4z� 'q*v�{�Y����rWm��#(�p�
EJ���8@㧂Pb���T/eR�P�5P
�i ����s�4��з�����M�w	Ƈ2_z���͵l�5���'�7O����"�֣��uP�b$hh��2������PU��Bj_WPM'�q�G�0J��?y������ޔuս�O,�)��4v�)���ŭ9��P��Q\*��3��q�B��#�5M��{�.���\ŗ�.�����F���N=�mq�ڭq��'-
*N`.z�{��Y�&t(���M>$��~�~Q��a�� �.5��Z��
���=Z����L����P�� /-� f���Uĥ/`"oH!>&�|��>@ۈ�	M~����<�m����ἕ��H�U��9���^�|�ؽ��7s����'��bw��j�
y$�n�>��⻯o�l�A���l*�!����z�-��3��W�Wx��ӉG����R/#�<�e�RM��#`��hX-����!B����������@·��>�pd�� l����x����o6�eN�2,��3���#�V]n��T홝~����dq���d�`MY'Y�/w�7ҋL%ͺ�a*�1j���;^�:Z��pX�{��7|��[R�̂22�pŊDV>̰�����<���}��ܻ�1�@��R��c٦o�"*w���޸����7��+�;��Ț㬻�U�@hL@C��QX"������T=ÂAfY˅�5��I����jI�Ϧ��Ϫ����R�baZ:S�������~׉���rS���r^�i��;�4�~L�j���i����u�	KF���Tni��2�űȫ��H�_�휼�y������,<o8�7|%%JGANE�ش���=Bݝ�Y����1 ��Jnn�=vW�>�6(m5M���P�g֡:�^>��<�krȓ�?z�E�\QAkfp�)�TD�0���ar�����,�������	�)E�	�,�f�U�%]ƭ�qO:1���R�[kK��E)ߍ>���I�+<X�n��̧��E�t,PyZ��O��b�r�9���t6��Ǿ�}���n�e>"�%�cUɿ��_�젇y�Oh6�2$���4�{R����f�9�ܶ6cgC�c�2C�K��F��8�ѕI�$�"�r���;�40��1Z��]0 or
ݧH$^r+����;�0�i[-� ��a���N�4�JL���ʬ	't����ɒ#,E��M���XR:��v�T�KC�b�'+��&�.1�g���rL r�>�.b�o#2�+����m;ݒ�CϦ�u�mI�B]È<})ZL-4�e�kl��dE���C}��y�w�����]�WZ�?�x��煮�����e������h�X8���`�D!�ge�%�B�}/�AE$){�8z&2rU��|����ڰ�eh���A��!�N_�O��h��;�em�b�����z��m�o�"��p�zO�CŐ�w7I2�)�S�Ϫ���6w9�,�"T�Y���݂�����1�e ���s8}���z ��?r=�ª���R'�Drh[g[{�jjs,�T%a*7F��ُ��)Tz%g�#�:S8%�p��i��)v{1p�"�T��;�3���=�{BúuE�R��N�U�\�s������"8u�&�f��l�aĔY�K,�(�ca���+��v{����gvo�Ы�eS���np�,��~��vL������Z�f�Q��Cئd�U���JS�kv&100O��hA�о�`�;��Gs��j�o�#@�ms����嚸��gif��k	��xJ�:���&T���k�5o�W8��$�`��9����v[��e����#�FP�p	�u@r:e�>����?mm�W��B��Z�4�)3:C����ա�C����y_��)�0c�
��s}��xj=�h����QF�b�
PI)4��V����<yp�E��8]�|E��PDw�fA>E��Z�cN�Ek{��M�9��B�
$;%1���;�é�vfie���3�.q��*��}>gNg�D��-��-M�$�N�Y�_�*�۾�8AeW���>��gxs�U;����H�7e{D�d��	=���*s'®���Z9s�����&�9@K�/��(�Q�(��d�O�
�<����i�t�>�����I�A���F	Lk��hyZN-�d*!y��"��<M%_*��\�2��^5��K��y�g���.��� �K�8�@���B-��e�g�m��-ZU��F�w����<�d�9�4��>~_��l$��.����׳N���l��G,V�0;V���ͩq��%0w3���:_�d����x�WC�3tl��nQ`F��A�:��L��F�@"D��f���4�O��%Z��޺��+j�vzݫ��I���1}䦼B,�4��cE�WF�v*o w"R�J%m��Ӂ�,A�9�ۻI���d��0o����_�1����"2د��Ɗ�GzV�D�Ï�k�S1s���>�i x�vW�����G�v���n��:<n/�_���'�;G��zţ{�,6���y�h�;������������ˉ�y��<�%�a����淹Lֈ�2�˖�H��´{�yߺ�7G}T���@>������L#G��0��,y��W� y��l\l�8Lw���
��a�8ܔE��u�q���'��.Z�B�Ў�e}(��Q�W債n����~��@=t�?W�l��J���֛�[g&Z�^At���sK��������ߏ�=x��G�3�D��;Y�#�3Ԧ7]�}�ظD0̟��h���9�b�<���&��ǧyS��qߧ%�����TT(�n�w��Ü�p�"�q9�lj�j)ð��=æM�b����C���%K�.�W����H���sM#@�1���4"��a]P]s���Q�tx�Z���ͻ�)��l�bc��#W��:3PO��r����ry�����&��j4FN�oK�����Ρu��@`�� ��LN}UT�*��سk��=#��ٔ�uV���.s@�[�}�V P��W��9�4.�E��'�2B���p��̢���v���	�l+������������a%��a_����޵
�$�"6������x��]�S����T<+lv�oL:���׊O�<_M�̉8����[b�D��#�H��V�k��ƴ��f$O�2���ƶx83z?G�Q�9��eP4��]�4�U��aْ�'[}l���2v�H(���5�d屏�8����Q�i��_S�N��\�l`�����j��~�5�N%c�ʱ�Ĥ��b�&D�EjR�i�n�vR�?�m�u����Kv���+(�@I����C�D3 ��XFZbw� ]k> ���(�+�}��tWE6��^YDat��A���J��aBφq�廝��'��Ao�+m��4}Fc,%:#5��F��AۭW��Q�e��F�Y{v�;��2���V���B��̈��K��ġ���j����6KTi̳�JG��E�B>�\�(���e��T�Z���42��$���h2^�Gd��ᤐ����z��C)
�e�?v�a=6R� |Ӆz�i����N \r-�-�Y�E4��F��Gi��?�wzLV�����t��D���]9����wl�P9��rw�Bt��//[B&��F깥��\���4/E��nĈRJt��h2g������������*���[��o��"`LX�S#�(�G�!�)6��Z�ߚ�A-�}Va�_]5G����Ð���6D��F>�i�(ţ�y�wMm΀��Ŷ��>
4e��^ʾ:��;O(&��4�TS`S�:>1&�Q6ĹDg}�g��	&���g�⵻��xC���� 0�����(�>��Ė�*�����/g�)sbSJ�S�j�v��o�� ���e?n��B�!�4��'����KJ�3��Q��p��j]�.\K��T�ݰ僑�u�4ٽ�����b"�e���1�moA�:d���C��<�}r@d�*)�<�����Ѭ#|���Plz�[���M]����Ƃ�a�����o��R��u'��.�/[�Z"�k7�����M#��Te4����[g(-����]�H�03�lO)��Jd����O2�U��6Ip��(4HΠ�$��$�#�� �,��f�K���,,6K����x@��ߎ����Y�5�Y��h�F�z���s%	5&�f����@���l�\,��<�b����\�Ʒ�Pw~�wɪ�*�Vx��`L��yo��>�I�{�!I�EĊ?����S	��_�������-�S�Vu��Kθ��C�m3�[Qw��ؙ=�J�9���f� ��]��7�D�`��vr��=����>ʭ=bT�Q��аOA��zI�yk��A����"���M�$z�f����(��f5Lh���W�〈Й���pt��Ka;� ��x�ՙ����$�p��ݟ��cB��Bj�U	�à���S�����?h�xM�|���	���s-
vх��;&�P(�����C�E7�/�}d�E�n�3�"�d�+̃[��M�P������k��?{�C�� �3as͌L)���*����>���D:�sTB�C�w�C*}��q�̵���7 !'S�E���2P!��� y�.�S��s�C�}����=��I�U�!r
��x�6��%��Yν�"�OY�������h �7��l��i���ؚu��~s�j|�>���d����:Q�b%w`T/յMi�fZ�{ڛF��j���m�R�;��!h�Tŷ�i��P+(�r�#�����k?Ҙ��<z�c鴆�����W*vN�D����?��zԂ��hn�X~۽�N��{���'��>B���+�V�����e��RE�d�M�d����7\�꿧pЩt��z�y����o�H�譯|�B0F-O��g,<��r�ü��LQP�$զ"���GDy'�e�F^~�������јˡ_�P���W+�6K[��p��ϕÀ�'9*�!��?���₲���[&�K�FVW��oM\{2���~$����:���,��b�h���������V����{��PS0A�"pv
M������	�Z��z{�L���H*;MW�1�&L�d���P���"��iD�e��x�lť����i��.�'�AZ��߷i������p�����yӘ���|t�Q7�>
�f��î$sz�Q��.��$/ �x�X (�L��Ӟ`&M;ġjU0� �oe����=��G�%ط%�A��L7�P�%N�<u�0����4�q�]Y �|�Q��"�[n#)C:if�hޗ'5n��;���#L܂�.l.���3H�ː����D�(���<�WM-7�7Z���S��[�6
>�YV�/���:L�)����e�i2)/�$cW�$1|x'�&�a�aGV@����-]�U��a�ږ�.�bގ�Z�������2Nq�UZ�aG^��7C�w=Tj\�b�R��E�bn�	+�L� �o�_:N����WibJ� ���>Ta���0!7@�w�ۚ��m&�8�E��!Aߠ�Q�d����Niq6Y��Tp���r
��Y)6QOa�Y}|�M�l�p�/�-���+���>����^S���s`Њϔ�(� �RJ�z}�-Z�bl��YcR:e�w���E �sf��]�Jtl��,.���g�)d����N!�oɏ�v}��H�D��37� (?��l:�f0�6�«Ϋ��悫'���|�5�5}���oe�d�y�.��̏�H���7��Lm��<ď�u薭�@H���2�֏y�o�[���]�hh�a-�GMz3�s�6GMN�!h:�c���lB��D�\%B��V*9n"�Ջ�l�@GGf.�2a@��(2�'�Ő��M�ȣ)��'�W�6��`�h�#�;O"�#��v�֫��6�A�%\Ί�;hC>\�k�n�����幉���ԅت�0��,w]��^u65�|���kKEC7X�UZ�k�ր���I��h����\�c�� 	V^���c�s���\$��"i�}��a"B�����c�,LJr�ތ�# ݢw*�&#�bŲ�fd����0�&:(���
ջN{W���� B$mߙ/S,01KH��-���|�z)����&k`�zAO��O�ou[e�O�& �`��1��F7���K��?i��L.�y�EVl]���t�T����s9u2�,���jP�����3��4V�������G�-����v�h$�:�_��E��r�h`��d#�M�s�q��� �qpRRM�L�e����y҅�����u������c���-`&fRp�b����@�+�8Fz�&�52��!��Ձ���j[��k��xt6޿��]��!�4A�f� m��9�&1���3�*�������/�i|
��B�N����A��#�����F�E\<+R��lI+f��p-j5X�o�����l[�<�@�},M�Ν}� ���դ��a������os��Du���4�ۄ<�]u�5�%B�ô����^��)�/ev���s�6�>Xʆ��Qi��Bl)�M�s�	�: ����]�m���6��_�4���V���K.����'���Տޓ��f-�T���������O�����v�~�)�/ԵfI��q4�~GP��@�%'>L�,�\��f�ߋ\ȮH���¹�Υo�ru8�R����� ��:Û�Ӻ9i��ngX��*�����c(.����^SV���о��Jh��<�Y�ߙy_��Pն3�˙
�}9�.�Zgbi��J0EI�k#��Z���U�]Q;ky�Q���������Ÿn�n����D3��µ!�^N�G��a���f�b�D�D�x͐Ƀ$~��{[]���T{� ���z`��v�y��d��9�3d;����x��2	v���Gu��,�9?#�e��Q�sn�(q��@��]#�m��f��r2�5�q��L�Ia�l��T��i�И-O�� �8[��.���e7-4J^G��Z�~g[�~�͠4�xqj��7������'�,���MAKz�Attsq˅;�4`�ٹ�L����*F��vY'$l����F-��w��F˒b_/ Z�&�%+��:��~ֺ6s��~&G�k�Y��|�nIq-d�d��Aw��K��~�s����U�5�R*=0��Ǡ�&�XoR�����$�l&E�y�w�$2�a��;�l
��������1�6��iQ�V,�p�G��݃��5B�1�P�N�`�F~&ڙL��vYw�O��1@��.'��] ��K�`�����B��Z�zLlcR �@
�K��@�}�:'�<��JK`^����(Dӄ���H�6csL���{����6��J��D:2�׉(J�ö����$W��\�+����i����ҥ�z�7s�4���3?�i
�^K E5(<�P��S:�����@�D�)ޭ���4h����ց�t�\V{�M�R���sӆ^S��>�b|I2bF'M�]@��Dg�'��JUU��p����eT�n��9����� 4����2��!.��������4�yb�@"����K��lXO����E��9~eu�ws�O�}\�Yi�B�8�T�6�P�*٩�^Iݠ�UH�(ש(m�/9^�F�_��������8DQ.:�U��̷�ϔ�d�U�Q=���}fk
왨�������'�&GK����_K�X׹��!qxC2?�嚤�#�J�!M#�2=[�Q�}�:���o��#FC��Ɠ]���X���<���(����+�d9�F��=�
>��(!S{Y%s��+�E��L���d�HrIH #r!�6U��	���K�E.��
���ve���ɗT�f�^����g�4�4Kߜ\y�y�ڇ��P��c�4tJ�����/�{!�SD�ifv���ιd/e��7�R�kk(.Gv״�]M���xLT��o@U������Qq���1�F�i1��"n�7���( 5��{��m��`dǷ�'�Q�F؋�Z�ܿ�o�w'�d
����N�*�	I���kwƇ�]�a�ʢh�a��V6z
�{f�7F�����S
�`���@C�,dq ��F��C&���Ήe:[�s�mH&�m./�{<h�Ό{����X��.��J2�}���28�Rq����M,����~~��/>�%SWz�趻��|�h_����	Ϩ�K_`<���� �A=5��$�J�;�jx=E�a��ÿ_�ⶉ�[ͯs�vb�w��YY/���aN�i�_ű��[�_�LQ���	UD��Qi�
�u�lW���h��c�S�^C|a���$�6
��K�<߭�~�0�����?)�V��j�X;n-t()o�ЊK��Q��J�nhw�!���@�8H�$��<Li5�A��mo��I�|h�7x�5�q�y5l��*ѣ�-1�B�ӱ��g'=�C�jk�����z�����-nʆ��=�ɔl �"?��Kp����D�Oؿ-x�ubI����P���H��$�ol�@�R��dO�a=���z-�xٙ$���8����@�5�~���,��D'��H���HJ���6�	��B�(�NHQ�"t@�*Y�сf��T�_ҏ����&!z��7��_C��x/:?�LP��"��uv�.õf�8c���;-��}w�����d����I*�C2pg	�i�+����q��\4Җv���3S�u�i�4���`M_��e�a�)jB�P6�%��#{�ٻ��U�a�y�������Ie�W3�,^��m���ty�����zy�?L�/�����h��zx<^84F��lm%Ѐ��+A�֦$�1.�Q]t�# F۳m<�����^v$��?��䋶�-,q��h�����
�bJ��^�/�]q��R���&�(�X-�?dD����I� �
����z������|$�`��l�`�O}A�I(�G������F�I�or+V7o&�r[Y@NŽ�\%~~�P�����c0�p�k9ыҫ�m"�8b�h����+��L���N���@���(��>y�V�z��GX���,&��l�:3fQ�	���Ǐ$�����x�[j�}��m,��g��	Y,ћu0c(!���L�o�e����?}�n�����c,�̘�m��R<�č��`����l^DcQ�H��+?�M�Dx���y��R��]ov�i�ӁG����ͩA����BA���� ����p���}�o�"a)oE��ǆ���q��&�W4����|�C���m��������^�7��Ί:��l�ۙUHˀ~"?XN^h7�p�t?���y��<������̲�J1ݴ��M	m���$��p��`�2o´&^_�n���<���c �3�������#��@��Z.�]�;-c����-���v�/�j���R���v���C�C��_ֵ��"T� �]��q�(5��j�0�A��<Bv�u�l�*�FU��;��^�@	���!|�i۲ҕ�����_��zp�T������T�?��j�3��U��0/_��y22��4Ԟ��9q9���#�5�{��5�]�߭܄&��5J-�Ԇ|��d�V�1h +��p5�_�$h�������S�DOz'��iM�j�ݚ�o�P3 ������m84J�<�'�N ������+����%
�]�}��R�T� ���X%&췵����6�,��a�_��#HY��t)�a0�ǧ�i��J��ס$�T _�/�wp�H���8�y�,��$��{��������ܷa
p�TZ�0J�a9��ʷ���Lrdi��g��	h���~�H���qsVO6�Y���� �x�͝+Ĭ�Pu��iDT갌�΋�`�di�;�����$�e9bf��EZRH��[W�"W{.���0��C \P�~&���yM&�b�T�P�P��� #~����Uw��r�8Ϩ���&���V���4ZD��QQ@I����η֬~��,�@�� �����y�?D�n\kICt\�j8ژ}�nm��@��6�����4g�V(��~ؾ5�f��>k w��X`���GQ�嶆,rx��gT��)����^�ǻ=yY�M����
�������	%Z0�]<z��u��F�GAU�� 'KQ�tZ�y��Q�Q*rL�;����of<�h���"��������u��٦qt)�lR���[��
0q�7HL3�y�.������I�j�aE8
�W���vt�*����i�T���MB���B�s�я$r�0l�ȉ<����[�5R{s�h�uK���h��ő����=�n`9Vh�so���Y���u,�p� ��r,��Ax��,�*�����F.yZF/���w�Q�i4�l����YQ����:g��R�
7`����yCN��C�l'r�R<{$pDp'T���#�<,6A� g4Q��ӆ���|�Y���|O:�=��T�D^�XyJ�n�,DY0�G��LM��R�\9`Ӳ�De��=l�E�����sJ�7�?���ծ��$�T2fi�z�;A�����N�j�3}c�$`����-{�Vs~b} �j��l�׹G4;��$�:uAl��(�����5�Oc���"ߘG�K�1U�ݐѢ�m����ρ��*���{z�U���I���g���:מ|�YK��m���S�w+��QK���_O�G�n|�"��������^�?�ϺlE�h��"��b��S�*Wd�w�cLvG\�d\�6���(��@�	�,�iq�R�@C�PZ�c��Q�QJ�o����y�^��p<�P;�s9@j+�j��S�4^�F�y�ț0U����0�����b���t�"���!�����UM��?�תV�fI&b5n;�A<�$ƳV�����
X������E��B6JYԑb~���{���ki�q�7u�o��SkM)�Ǜ��'�}��j#!����8m�L5����p>m�j7}Y���lހ^ܶ��'�5zn�E���@ܔ���~�La�j�xWJ]���U}:��z���
G.k�v"���9�}W��WF�n)��AX
$��� �ګx~(�-���S;��+��~/�q�te�� u_�jSѴB�w�(�=�2�e�M7�&�׷�C
*C8g����{�hYOwJ�o6��hKXox�c��I[(y�����V�-��Q}�ʶX�ݜq}m7�Ԯ P�-�K{żYl�R�P����?�3�hvau��EA�d�]���׌��r�F!nx2���>���rU�W��ȯ�M�GAo�O*[��Mu�u�{c����I��V����!@|k����q�ac�fF�F�Lps3���{Z`�ot�-����G�\iv�X���j�on����z|����c��Q?�6
Ԭ=�,�׆@�tJ>q^DsS `�db��+o��r�[o�0���PZc�S�Kz�u�VҨ�����Z� ���~��3+�U����wA���PØ��Ue	{�FNe��X ���?�no �,���������[��� �M��˃��C�׳TB��1�0�~D!�~�H�P���7���7xj�4\���)�<U&�ѧ�{O�:��v�hrA��p�6�])�-�'R/����(V�$��#n�ab�`�p��+�[|b��@�9T%#����n�
m�R=���z��e��u�sw��6a���o�+�E��>w�m�V��G�1$p9����v�����l�`Hx諹\�-�s�1v"��
1�N�S�Eԍ����	[U'~B(˳v��t��O��+��֎��)]�db�� !3��q<Xnf�lכ��_����^B�p�b0��K �3�ս��2r� K�����)�d��*ĺ�K���P�q��M& i̒���V�`�ǵT� 0�	c��'`��6���޲�84S-�>7��qxmn�7>u	E ܾB��(	�?G�k>xU4~Y�.�
�ܠn�3f���:7�+���J�`w��0�
t1���,��� ���a4���c�ے�6���>I������
�E�1y��0vE��P-!��[������(�����D�m�}svM ��#l� 4fŒ�0r��u�Wc#��A���I����0&��4�K+O������_��Q8B(����\���b�F��X"��k�0	� �U-֡.���$sI�0'�G7+���Ψ��������T���o�8����ο�{��#t�Y�'��}����;V�lm2��T�W���h����=Z�����O���I�1٪�7<2b[,	p��b�,RntiͣYc���";P�F���ڶ����_�{�#Hy'�J�@~]���к��m����Vc�ΔF@�xN�w�lĢdn{����QI4�&C��3�]%���]��X;"C���0��G/��g�@¸7fڣ�8�X��W���k��d���I0�CU ��un�Ϡf�g�x�*.�l�J3�5�@sm�R�a�IL>��P���i~P������J��`��]�R�%��[�q;�������ot���`�8��4�z�.�'�h���$��<E�uD!�ЃOrH�#l�f�c�ʧV}��zh�5�f4[��ڞ�>�rb�d�l��G���ꢓ1��@�@�i\�9��B���z[��9<�E�1|c?V=�<�hV4��W����E�ZcR�|�<SC5ϡ�� �S��kDg�A��l���1n! t ��-{�����(MUcC^K>q�2"�pǗQdrv�C�>҃Ѵ9K���(SD�@�N������G�%\}�\�F�.�W��Z3��TYX�(/��Gd;��t�#���Z�����v�Rp]'[�L��0[�k��w1ۇ���צD�͕	��B*���54mE��82��r�׊U��J�B:�v�X{lK.YSV�`oI&�Ĝ|g>m:�PXeZ����Rt�����p���;�X3K��/ר~_��O#��qe���~�JȞ�Ұp��w{��m�BR��4*Dc��'���W�'8D��˜'�7���x��K��\K�R��f���j���D$�q���;�;,dR����v�T��֥wq�g/�Xdˆ�~��T�u���[���D/@GĶ���}�' ~ L��W���R�G:#U �@'a��8|����J�[���}�1���ka_(9��!�C���bB+N�\3�G}��'x^���6%-�ar{B�����2��p�p(|�R2DJ�zL�W��w1��<�׶����w�1���֍���ĘF�gp�$�Fj2J'���jWV`<zme�I�<��eB����"|����d�W��3������1�M����e"Z������A>�ghOc���2�Z�/����y�ej6 ���f'��ϊ�Md�Ԓ�Ѣ�����^�(���ܝ������S�JG�Љ �h�� �hQ��}�s\Q<��1A�g�.��o���9[7:� ��4���m ֠���AA�>���\!�WWs��MǱ��U덷��Z��Y!��7�,�wM&I�@8�;�\�^���w���]7`�<�U�3���5F=��e�������jC��$J��eE���E�9����``fS;}wk���C(�E�hfX�����ع��o�ݴ/xK5��诖DD/�TG��Cs�Y�I�6�]J�'m��(IM����6!o=��O'�g�&{��
�.g���"���3�q}��~ӤݬrKp���j�_A ��ݩU�k�v:��%�����@�7[T�,����i9l{���#�~��ī�ڜ�J�S�<kT���ÝpQ�����;d���ӗ·-6�V�U�b��.I��*Lø�ף�S��˹����g�;�0�ST�g�/5�Җ��s<�����<�G�n����JK,gZ���'��r?+�u/��c��6]�Xn��@�4����C��BE��b��>Ò][����j��C������t���R�{����"Q�����7�V�0)9��=�CA,��}gx��:�+*�b4��2��Lr�����f׺z����p���;tI�¥K��m��M�޶uq�� ~+���pm��ACK1~o�f�A��Z�W�v �S�M$�Kئ'��b}�EԉKUCQr�j���ht,Qg��3Γ� �@ǔ��Y�|����\=u��k��<�c�]�Ȳ��I�X���~nM@#	���{��V�3���y�A��^q�f?��*g�͋����ä�T��NNk��ě����9*��c�J�:�h��JbV����M�m�]�����J���� �����N����$�aEt?�+\o���.�#M�I�O"�����:�4;Z��+V����(1�Xה��<@��g޿�i�4��T����{�/�_7�V7�:d�쾣��e|��`,b���:P�����2on���a>b�K,0���1Vqb�x&I�L.:���X��?��蟅���Ѿ*35f�aO�LY�l̀��(P���q�9
9~�']�@�=��[S�g����Z���Z\L�囝�ǵ�4$zH�ƤG)�#���K2�^�	@�D�^�5�㜖�<����?��A]�u��^¹e�x�UhPCf`�9UV|:�QOq2ѫlYY��L�me�a���1��{V]��<`���8FRn[���?�Wd�E6)�<�REx� �����������3��8�2Η�C~b <9���*�q�Z�>�9�' �ɪ��S2}A��(�D�9>�^�!��P
���F����^n�b`u�{��n���H��4�Z���� ���� �����~Y�W��Y��nٛ�c�2����'�ٰ�"bZ�`�B�����Zs��$9m[}\\Җ���|<F~W�7<lL�O'�0:\]<.=�x��y� o�A�<��ɚ*��=���.D����Z=��ꤣɠ�A���	�����>-�}�%��V�l��4����ا/������v���|�1Q���"W&,���3������*K��}�ڹj\�=��	}��j
P���*���ۣAS�<���,;<8�ϟA&�֧2�Ð�)����D3�{7p����[-���5�|c��}/B����j��[.W#�\����J��4���� r�]&��Q�ƌ�
����-�3���ѫ��A!�<�	Ќ�xn�K��d5�En�`���&]��({K��\N�/��~�����e���Rǀ��Wپ�t{	��(ۤI�����!�Jv햑@%����pO=�����̢6f�R�]J��[?�+��M-����V����޲�ٜ=v�����P������y�ϩ\j�П��S��s5�"u��(��-u[��7��ex���F]�SrM�eA�)��!o�2�:2�@��ѫs\��7Ɨ�I��XA�`B�X;�ZS^2`Fh�(Ï9���ӕY}�a+
ė�ȍ,9����ʮ����EoF�����x`�"�"������Q��YTPK|Oy�E��u�ߓS�k�����YEu%M�*J�x���eo���7��%�ɛem�Fl�s/Q�&�
b�\��Y�J�n�|"rHs��5 �W,�צ��Ra~ј��C�U��C/ۢlB�j�;����>�J|;�>ˆ�n�D�A)-�KR��Hd�0l�����xr�ef�ʠ����c��IS7_^ +ˢ���A�6jN�t��o$'ϯ"%X`<|Q��9�nc�QJ�����x��sg�t���FH���t�s�$o�b�kX�,��'Qs�uv��w"�&� t�0e�ݕ��MV�"'A�W��T@�߳���%�3�`��!mfH5d����	�o��T�x����.�����9$�3�'�-)��H-8�I�����(�L-MEܨYc��a^-(f4iu*0��Br3���3�r$���_�j�[ru����`��>�Ch�[ݻ��hi�Q+��p��wYq`D�@�yG�#5+7��Ů��u\S�����7A�F~zM�D4�7��q��ddʪ~��� ��p~��V��@�D�ˬt�	�E�i���/��KUx��t�Z �_�g��7����G���C�;m�V�&jp$���j�焆�Z4`0$w�5
�Dp.y�f�EJB�L��.��V�d�SO��-8�7d�m~����`��qJ��U��:�3��*)��$ral&�K2��\|Sr
n����Jl
�6�0̠��g<O�Y��̧��Q�z�%��g$��y3��q��J]z=�(�hr�6�`�P��j�2я��M���(�����@�� m����bf_�'2���,����.Ƴ�L�Ή� M���փ�x�&Z�,���H�YX���¡k�}J����e�B-�-��Q��Zۦ#��|&���n�����e���l0w��,E���DC�[
�~Kv��`M-B�M�a9�����jww�V��<���ꄘ?jsH�iX��	R�W�1��cmw=&�L����v&���dN�,�����pۜt[g�ъbUY���k�C̅�L$C��޻��[k�
$��w�a5k�Q�}�ݢZ�-�V����ݬ	�Cu������is���׼�Ε��|��pc¿�z#�N^�Y��Q����p	��/��]N�(���}�#^g��^O��oX�""{\�TW�\���M��Hc82 $9����i��(���*�9��x��-�CM����f������T�#נ	2�%���$?/H�F��w��?/@ j�F�@Y������b6h�&�c|��W;����<�"����k�Q1�$���l]ͪ��h"�3u.U���W@Q��`�����T�W�7HM�8�+��Pt��gid���:xS@�N8H�O���R((�`� @[�4 �� �� *K���];�{Y�P����^��g�-�Hf`?��'�q]%�{R^A�2
xR88�҇cI�-�*̫�'�*o<���YO�H�uÝs�Y��:��!���fG���9d��s����ׅT���p����p��hZ�6��+˄.��P�X���.I�XScxo�Q����A��-���'&�VB�Ԃ<F1�p�0p��N����G�gP���~zO���(��iK�I|�b!�x�����v��k���G�*���}N�B�O͕��'��Î/ܜ�]T?����3��ԪAe�7�Z�r;��0W'%�u�9��P�v���9`��BQݼ���J�4*��W��m�]�Eְf�B�>���:�,$�]6�K2�|�����&�i$�g�$�����eÀ���ыċ�?��Go���`S�/�(��V�q���8��y�b���뻻�.������1�9�p�O+�3V�As~=irA��>��d
u�LӸ�v�h�,�H�j"&q׈nu���6�)�1]�H�,b��0�Rg�RC�0���k���#9	ҧ��r��!��y���P�Q|,,W�0�)���z��R�FA�{��y�;o]}Zz[I��9��o����ڱ鳞�����;\dC`�2�ۨ����Ūڛ�-+M��A�! �.s��m�;'�rc,� �
��v� IN:��� ��������ށCr6P�K��*=��ң���th]|�Z�`$'Z��lӅ���p� 4�lf��+_7#~|��gk�������vdCJ�7�m�JCe�L-��,�|n7s�fŗ'[��k/�f|Q��僠s_����* u�5�A�+�
��g6�M,Q�����PVJ"����p�q����0:ӢEp���V�9������A�H�:��0�y��h��Ο��jۜ%ww4O.�ǫp��ˏ �n�k,���P����#���ج���t@��#�ܐ1�GM���_�Z��=L\O+o���T�,A��G=���.�5)�&�������V�ب�=J��P�zĎ�����a�敜L ���U��=�~`@�����-�tλ?>0�X��n�	�v-���
\������q���2�@��>ܘG��ή�D'�01���(�#D���=˂ٳ��or���A�p<�$<Հ����^����L����!��a���`?��D���H�^�D�n��f������Z(�ֶ�f���M���Gb�MV�9i�pjxYg�D�@���[�����LZa}d�=��XJ}�A��P�WN��*��1�ЅS�GP�h�-/<�},��rO���}H�S�GW�g�G�C0���9���a��x%aE���_��}܈��Y�� �\[~1O"�nd�j�{��wx���9�|Iǫ���J��L�2�jTю*���J���[q��t�:�,�)�;�\���kD�ld�A�
}�@����P��^ƒ�o �Y�_��Lc)����j#O�aκ@*($-������"�II��_����������Q��3"m\�J�E\>,p��Y.�<���=��a�s������!��*�'����m0 ǂiyz
t�5��`>+�ԄY��|t(&��/��Нq��s.��E*��x��/� ��uS�\�#�
cT�g�=0�N־-��a>1N��3��(s��^.
71��	��܇�Dm�(�M�=�Iɽ���-�Mk��`�{kiz�|8#� ���5����$W�]~����2�f4�L=+���S�c9:I-�@_�P��������d3�qp��� ��[Z��R�.��Q󀋩Tu�
�V�O�� ^#9��̣-B��s��&9Z��P,I%^�u'y4����aG���^�,-ZH���ں��4N3�K�O��}�2	�6����+�yG�9�Yx'�^�G&������63�I�V_\k�:���^���!����h��w�^�,c,��7����`#	��
K���'���^�$����Ӻ(�B:��չqZaB��P�������I$N�&��<��y��OYx��mZ缅:�[Y���W�y��6�1�H�,HK^dׁ��������Z��1 ���_�by����E�A�	HV�� ��԰���0�A��"�G"����F	a�Qd�O����(��i������$mM3��βOm��坧nv:Rl	mtz�T�.˼��gyȳ�����Vc�U!�/Ϙ���(_��6��a;C�a�;v4"Sxei�vW������7�nڃ+q�;Y����x�a�W��u�*�'#�]$A�ɨ���抨����Q܎d�����Ω���,�g�����O|�+l���;|�+���Fqi��M��V�7� Ci�4�+��=5���>����ڿ�����Z��O��$�4��2XCTT�-eƖ����;��k�7�)�_RAu�&(�8�e�������͓rx�]X��5Z��e��d��z%�\���H�}��w�9��F����}[E�\��(�14� �l������&00����sw�|{�1�A�J�$�B���
=��ʖ*iI��A���р!Y�V�$�O\f����m7��ORmuk��G'��7�n0��et�FPl��t��U(a��}���"uf4�u�
�4x��������b�CQO��Cp�G�v�uP���9t_��D��i�M]�Ћ6�#��q��r���f�T#~��Je	!t�*z$����k$���	*P�2�|#B��܀��DGb۔�s`���`3�H-�i�v���;�3u|N�j���f�<��	����q{&�C��<��Α���ƣ��e���2���F |���(89���>��5괒��[�Nr�3S��v�u4`���!��I^˶��?~մ����3v&��ơ�eZ�//��5*���&w2TB
���W��;N�W���z3P�%�,&�����Z�_��E3��?&ba-	�6k�0���Έ��F���HsC$� ���?��5H�E
\c��?���Z4�8������Q��-��K��SIУ'���F�^��BG(Ye�a�5�}g-/�|Ar�z�?N&���OF���H������
�M�F%�9���'�p��=��~VE�@�/ڮչ����iA�Ԉ�k�@�9�nMj����>�Cg�{zI��aGVi߈�w�"<4�Ż�g�R��¸�+�����緈����R}�h���IP=�=h����"B�ZE9��q������x����'	U�NY݁@
c޲���ɗ��M���RCK+��s��)�0u��9�4"�z	tЇ5o��B�{ �����&���u�`}[�-ꑮG/��$�����f*0u4Uԩ2PL0���)��������*�Zdq�5��,����3IQ������py�p囦��Z:�u��b�����N�'�Yx�]�(z���Z�>�|����DbL$����)�o����y�od�p�52�F����rl��>s�?|a!i�E�9�scp[�
ŝ�ոw=��N�;�Y�|;OM�CR�vZI\���73X�j�QI�)���F��n�!,N�n����i7�c�4C�[�޹��z�2_����벙�T UuNQ3�@��6��R�ZH큎�S��]ё�{ L����KE�p�ۡv����(�U\1.`7r|7sFK�:ȅN�$�T�t]��Y�=M�\����S�Vsh�D�U�U���Ů�U<iŸS���uT���1|���o�j�tf#-0�{�bn�>��ߖ��/�2�!1E�B��:�ه�7�B��0��]�Nf���, e+��I>��LҋNC� 3L�.�������F��r�d,+�)�xn�|�l�����������<�whf
Q�լw�?T��qO]K�#�~�軓��3Xo
��>1�8|b��O�ٵG=k��|7v��H�!�NG�A��Q�k�r����k��M.j��<s��{]r�4F+�.�%>�K��Z�}m_�Я.��x�0�T��m�Yڣ!��������(