��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
���ۧwѸB�;Q�)�q�ǥ̥N�y�7x�S���1+��Aҏk�A�hg�S����	�㳰SC�����Ylj�;��Ɉ/yl�Xь�}G�X؊����;�'��VG^:0�y��F�	���D�:j�k̷��u��F'U��X��ù-�h��b`f����#0.�w�N�st&C��Z�V���!: ���X���h��.�u7x/���,��� e�����엙,�Ѳ0������)��������in��&�y���F&�:������q�q���y
9���`�}��f��9�'S}�@ 5�U{�]3O:���[��x�+U���~�v�_}v)�>��
��%����:yxjD��B6���P^-��T�/{i�M�;�X#���"_lAMP���8'����e���d�X_����"�D[䄩�^�3�J���SY!��qq~�����T다�|�d�*�d��m��c:�n��^�+����=^6�zٳ`�H&`���5�[��t�f�o��o���LO-�Cم�_ρA�plX�vV]d� �710�6�')ߤ{޷7]��W��v��b����]ᨔ�3e�67�᱊t��V�V2��t�,��-�L��LM���4�+���f� �~�6�%	���9�NM�8�$/�^ږ��8ܛ��#K�tZ���	a�C�67�T�^JO���rB�M�$�^K��O�==�Dg��9g䴽�ԧ�3A��k�T�<�v��;*O��)\Y�p��]�c(��1a�����dPǛ�I�B���ώO�(艤�3�ão~k����\���~4���J�����)��55�&X�=���2��.��܇Keȭ~��[y=<��N���9R?>oȖ"��2(�f�!�8�L����w	�k�$��&�Q��j�&!`��&��fN��벌;���V{Į�x<���:��z9LK+���1��h,z8-GxIS�	�響�-AX�M]}�u)#�4T{�����â����_|�$͓~(�>����㴧���N�`d�II�m�,��G��Y�8E���'���.��n8�?��\4	˙�䧄Ͼ8�m�Z'2�C�.}UQ��]������$���_M�P�;��,&��[O��t*@R���ѿ;���I֤��ާ$�Œ��u?�B���w�I���&`�Wh�L;I���mc�>Z�W)��:��@��!�,�1�hVU{�d*�#�%��CV?�»�WD\DJA8(�ٛ�`�y�k�+Μ��!��GrI;]:Q�cԱr��=CH��C�����.��KVʎ%�^i��ls��2����yN�P��-ӧ7:�g%6�$��
���c�FG�K�k�/�|���F�g:�i���j^�f�~�k:L�Z��p8�J ��n����ewҙu���ݠ�'��=]�n@F�k�)*O&���!E
��W����b�ze!����SK��n8}�#�=�d�>�䳸�A���'=�NF�����3g���b�����q�@���;N�7��N�:����@OfH�LLb0h�;�!R���[�U��
��x��R����� �l�<d�!�,� s���MT��S�6���edd,��}��?B|�6�~�Z5�I|����ϵ���ϡ�:�Q��
�q�j�W"��7�^M��0���S2Pc�嘕~��|l�T��E$��j L;�l��2:�B@�ȠT���6�В�2[Ψ�:�O����6m0{�,sp�-1�ͻo��u��@��]��2gR7�Ds�s�n�[SL)��#��|L%�py$1Q�#��A,��X+�|��m��I�ˀ�K?*x�m�/2�x�<+�/i7T�)@�Zv��j���`��Z��7��q��� `ｱ���$C��ܩܐ�������T��a���������Ң1�h�l��%�O��$� �$C��S5c!�]@Ue��Պ,��y,:'���`��=���lo�2f�+����Jc�F	ښ[R�-�Bx<�$D��XY
�6�4�I����2�u>av<	P2���7o?
z
��7��w�@�/�����(D�A�s�[=D�;۫y2!��Yo�v��$��8�ȅ\�FP\��M:!^�in���z&}�����R'��^UP����~���ekPɗ|T
w�D�Y5��M��@e���7-�rN#g��
Y�\+���r�7?c란�t��j+�eew�<�@*{\�0N��Wa�iX�r�&]{f2�y����3���c��s0,���_�����V�39O1���`�c>l�����!}Gݺ��7�n�Y�Jur�{Šɡ}�������"�.�|�?�I}A�8���*�K�+����I�Ҝ:Y;$�R8��]��k2}��rp_?[�. '�-:L���tc��;^�6]R�̉B7­�2?y��2^�w��c�׋��U�O6��k)BoQ3�\���ǎ��p&�s'�+;ZK�,�,uɃ;��� Kk��y�Ѹ3�D�p���a��/m/�^J���Ӡ����G�3촬��G-����.�M�k���-�ZK����YCC�aY�׈>d�~�����<6n����)�f��+��Y!��X��k�\+��ﲻm����O͂�a�+��c󑯒��$�n��������Mt����[��^��ø�����f.ٙ�N7
s#�k4��ا5H�N�)��J΍j��v�� �{�`A�z��� тNXh�GU��k�h�Ԝ��G�	�ܟd��e��<���|���� �ʸ�$�n��),@�ҝF��l�ć�Q�og��K��
��VE�Kr������T�%�V���Dr8��S�=*!/m����c�XAȐ��ɞ�#_5�g˃��2֮�����Ӆ�i����s��+٠��S�3�%n��F�M����v_��m
��<�1пS]<�r;��q�8���{�nU�*�/Oҝσ��Z��=�`S��m��DuY���P�qz�x ߬^�<ѥ��Q'��O����Y�Yy5����q�<B���[�t���<'*�����T��2��_|�)ty�9�-i����\X��?�N��2�kY�}��(��uQ}�j�e��fٵ��x�<�����F�Շ���u�g�#��oǇ/�����j�n�q�4�\0`���e��wzݼ>{�W�ʖĲ����9�� %S$���2F��B$������k�*c� ��TȻ��o�� ���Q��=RG%����/�}��LG�*&�?����b���{.
���v]BewЂ�@L��m���\�ڧU?ʽai=A^���^w�(��\>�h&o�(��qנ)Wb�����	��q������T�'k�	�ч�" �B�I=��r~�R�a��ܠ�v���A�ƋЁӋLƱ�	=�)����~��"�ֱ� �Q啉�jig�����`$<��U�lhe�j6�ܔq���$�kPj��~�>��M<U�A�I��ZR�}Je-Nr��W��6.�)�uc���*�w�qm������T(�����aj3Ȅ�q��w�S*d�!,�=�ޛ����7'a�Dǌ\>�њ�lF�Sh���C̛!%��� �� v|��xKw�<��Q6�w�Z�J�� Ye��N�t��>?��f"��i��cxq�ok���5�?,sóiߏb(2F��o^��$���E����C�+�X�9���p��o��i�Qb��Ag�e`�ci��V��Y�sX?�d�[��?��P`�t�����h����]��m@A�w�ӻ=~rK��/I�~����(�\9y��F�6Y�F����K?�H��&�b�|�Un�kb~Bf_UH�,�4�������|j!3wp ����	T���}2f�'l5N��&�=@��������k��b5���f�#rc9��;���(��M�Q�������G9#�Jg�D���Uu�*F�w�<�n�G��b������0Tq�͙��=�zQܦ�j�a��O��G޻H(ȱ�WB��]O�(�{4�`D���;0�[ }Olќii���mڰ©T·k��ⱅ!(����0z�j,��k9�6��w�&�㞘a�Jb�S��5�͢��"��
��<�yn������Y�`��J��Q)��<q)���Gk6�6�N0>_u�3����;��Tm�����Q����A¶�:jA���[��XȐ�e���5�D��Dg��'���Vp�D�kf�:��nG��$�/�h�O�RjW�?2�+m��L(�p�@d���>+'��X�~`/���+�ew���������\��C>����q���20��V�� 8�.�f����G4�x��o��+얰˳�Z/O#�ǋg�
�a`tD�s�;k�5c�U��=r/��r� ],Ȟ=����ϭ?[�D{C���ꄞ�����7	s�!���Ȅ�
�9��;$k���?Э��b^Bn����x��� �3�Q�N��)��fQ�3jӧFX��eZ���yy��3QM8�V ����e�<ta����cj��˛�ۋ}�6��݀P�Bg�=��2\S㵛�xL�W���|]^��ׁ��'7�b᫤Y��T��I7`��b]Xxy���W��'
0�v3���9G5Ӹ���8�1���V0�G��,����-zv�V��Y��xг=�sb!l�j�+U5�UZ��0�>Wq�����ҥ!�x�/=�<���䟇M�:��5�cbW�7@J��VnȜ��9QoC�-#��~�@����K���Ґ;�M�P�@j�G��?G_�&0x���~	��>ZR0��X�".���5T� ��Ѕ�͈f�|?��V������_�҄���Wp�1$���)'�-S�4��[�}TY����	J�%[dݪ��[�Y�]tN\P�!�ӡ�Gd������D���4���.���x��C�B!T����`D��[}��I��w�n`��v��R_9�m��
]���w!�K/��x��d���/�����8)���L�Q��%7]��/�jT7�Y�Jk�9f�N��q1�����1 oh��	Vg������MW2��Q�6}m�N��-I�F�B���5$Օ�d�u̠XDr�ͭ�@f{QȺ�H��w18������ؑ���;��l����9��FәM�a*�Ph�:5M���z�P4E4�S��·֏B�������P�4���"U%č߃��l���G��ںo0:�ǯ+�/��
�7�3��~�@j���2�W�h���)Da���a,����8}"L^�9�9�aVt#�1���Z�}c��D���f�o���bw��(�:A�9mDr�=� ����=�1�ܑe����c^����w_�+P�A�����>��Ͱ�x�K�������Ⱦ���\=F�n��$�9t�j��q�Ը�|� Ƶ�E.�I��7�w����L �B�e ��@����P�M����Ё#����{{��gS��X�sԅ� \L�u�U�O�F��/i��U�ᛪ�Z��#)?����֊��������	��:�(������_]�NZ�-{�/�[��%ջK�9����A�NE�q\<�[�	]����0����k�_"6/Ʈ�M�c&�v1`Vm���9������NFn����h���j"S�D��H�q�5���0�'�3�({���i�-�~��E����h���<K��d�I �Xu����`P�����Ґ���{Xl����0#��m�T��[�C#(����ش�eJw??����{��Ê|#yV�[۷`F��`�K �cL!�E@�S2��Q�{�8��FV?J�[+[Ei`��_�3��U9�O2+~�XZr������^UF6�I��RlP\������4h�cߧ�8�*ُ0d��R��`Zr&�vH){T��ki��5n����K�c��j��-M�ھ��:��nV�m�X�K/��QĄ�IWH�*rG:9��wX�1ť��Q�/Cn��h��ƚ+w?�A���v��q����|Y>�c�E� 6�˄��.�p�^��4�yэ�!��3�$�bx~������g���;z5]�N�G	J��a�H$�6uQ�ޠ�a�z3t�̘��5>@BJ2�:�<����3U0İ�\�2 {8��oS�<��i�\�*�-���B��R�b�N�۩���SH��Eڈ������qɝ�gnK�y��z��ک�@��k�b�����cfUt�g�7C��YZum���HW�!sؚ�Af�B� ����/� Y��P�l42�8Shg5WQym�Q���i���O}��L�{?�m��IS������c�-�V�g�h�� 3�״��?f��0L��(ly:�N�y���&\��A>�W���?z5�g7F���c!�h�Fߢ�S�B��>�0�[�ԏBP�R��7�6Wb����&��]�+}�f��{�RVMfv��8�Q����JPW��s����,�n�� ��{>biofm��dK�S�bgAAomS�YL$$����AwW:���_���2gS��iղ�BXVS��2Z���א M�a����6;�Qn%н�Ch���`3���r"H��T�0!��epdJ��'���)�5��mNԁi���)�R�mS\����|L7�%>�9۩�Zh��Z�$&0�v��9/���U�@��i�i�ԥ Ӕ|~ 1�
���D񝧢�į�t��������8�O�^�3���J�����]/`�#4�e⬛,�i�B�١{�}��.J�w�&�����݇��W$�NՖ͑ĸ��.t$'�ף�Z�+k�㙺V.��w�CᏀ�i	qs�r���<�)[a_:O]K[^�����d����5X^),���!j�ep��~��m���� �ja��x����?rng���G�]�2�v[��N�#���Vs�ʂh��g���k�6v�ii�̣X�<�2�$���� 8�=��?KO�87��̃˭�w���	�Tpr�� �*���k*�ŋ�ʮd &^>c>ؤ���Yv�e�B�����ȍ ���x���=��rE�<���n>.�#��`�@z��-3g�Q_W��2��e1!1mP��
i"_��@���f�Ӎ�.�ɂ�OO�̓ŝ� ��pp8���ͼ�@]s����|`Ȫ�!S��O��к/�׸xJ��zGN9�@yw��#����y�){n�O�ʌ�>s�f���(�7��1�D�z*����7�)t\������Ϟ˩��	���l�x��H�OZ�o�WٞOĖ��B�1�cP«Q�}m��I0+�<��)�����҉�����=ܒ��I<a�^�N��.�5�U���o"@�I��<��� 4N��&��%<�b������CW­�'N��0����jI��G�f� ��,�J�C��o�����x0FF�g��䙄��Oy��a�4q5�j;W��|$�C��}�f���x��%6Gb��"C ��9&�^1\����x��(c�ԏg�.yih�,0�������O��fH�&N4�X#V�(x+#[n
8��}�S��D�N-/��g�UT����0"�xF�@���`\�����{w�؅���DÚ���� �cҡO`����9�Q�8%0GB+�nrLȅ�*ؘ\)H>��C�v��28�\�?�:���:�f%�D҅�1�FoT&`��Ϳk["��H\���o���xA���\~3�i�%���4Q�r w_P��iZd����}Ai�l�{�'���j�
�!�j��έ��eq���5�	�I'#ğ?�餕y�:T���pը�f;�����h�<��y���O\&[�9�v��/�Q�$)H�1��H7WBq�@�H?p#�]�YFקp���!O(�m�7�
w2<��nz�t�%]��I��U���:(��3x����o�kaή�>��ơ������f�¿	<ޘ����F��p�MF�r�R��z+��H����*0?m��m&��U����];VML���l�3��j�t�Vߖ�F,�c?C�b���G@�-*#�x���dN;����on߀+R���=`%�=C�.���X�9h���9
;_5��AYt���������Ԇ�+J`�ƃD({M�u�؛O)�䉟�1{���\|6�F;�qd�.�I�!�7�
����3ߔ���� %ai��|a��Ť]^k��P"�<��i�>��sY�hA���2j�%��q�:t3�����:��<���f��y�c��V�h&��3�S����Y��ɽ��(���t�E���ʝP�	����ݧ�>`����@\W�����٢: _�R:pH}&�·�W}S��t�Ǳ�f�m$�*L��^̍�i������p�!~iס�B�\�_��f�e�h��O��_ѵ��>&���L[�K�6N�0�ٍEO���lgF��{)�;��Is�G%�	��u�7!ъ}�8Ԏ%�E���K�Jͫ�Ób�;_a�1��#d�{͑N�y���^��,˦�k���=7s�AI��uIR�_�c�t,Z��F�T�:�P0�$7c����/S1���V�	]����91�G�����Aݠ�{��,{���|q��@�B��+�kW�E��ї�|�s{�meqg�28�~��=�wk��I���I���_��=?؝:��*8��:5f$��	AZC'CHR���fR��(e ��nh���#�_$���攰�C�ij痚�
�&�ٷ��[d$d����ųjA�HG��&�ih�xa�d��aӵ�KŒ)�OF�Z�|d���f���A_i���O� �!m���J����TQ#R� �ӂ�!Ʊ����N�)h<��B�x`�g����x��L ����֨$z!�M 
GM��gDCu����M���s�!Y�q<ܲQ̷�j��U�+�N�u�u��)�n���T��t?*l=���x��w�A;��������+w�5IO/��.��N�n�lL'yF�Y�|�\���d=:�Ո/E)4��4i+�Ӭ4>�K�M>�.,J�r*�a���G��=�+�{����9K � 9�ӿ6:��$0\��w�)�t�}j@�ج`��Nϯt.5�o��.��%�����֧�E��Ia�����w[y�h��w��fnX����E���cF�k�x6����@\�m
�v����ap2qk=1����i0�B��=������"�����E�����[&���_���,�����-�3������	�X�gs��@�Jtȍ����_#���ki+a��h���	a�i�ʇ��$���-jqk,e=��"4#��/V�c�5�y�m1[y����ە�!�N��$�[���J\���h���?3P�p6г���?;Pi��q<���**2I��:�qc��ق [@��(�U��q�PUZ8\��i����.d���x0��r���?�=<�_P`�JKMS��~7W͉��6$�I�ήs-e�qxf�OqD���D����>2�,�{�}D��u�p;Ͱ/Q�@��2�Ba�+oqW>:�$�����3�0����X�C��ѽtᶤ����,�|�!|)��8��a���՝d�����|�.�dy�:��@�	��;��'�Y?Tk�![i20hP4٩�72�ɢ�X�e��OW�y8VK8�e��I1<haOXW��:)_@�*}{{ɵ�}M�C����VO��d{Ե��O*_�
�"�$Z:�O8�Xcw.�D��؀�పI�/"-��my�g��e�.�aHT�+y:Y�Jr�O�O��Km|bNIm@2o�x�'�P*a�[�,�=	���<�	��������9��'�[J��X�bu
C6o8h�nӃ>~�D�T~.m(%(�ګ�5�<!U�ﲁY��I��d��� ���3��mg�N?~��ًfPѠ>���&�G �{����bM<��9��8���� �Pz�WE�#�T���WF�D��9DW���
��@\�9�\�酲t]�Lk���^�_��&��f���� `����D�-9ď�	^	�v��\Ӆ���j���Y #�� ��2CVz�x��4�.�c�����K~%���N�%#�!N�3L����}��G��7�V$I�a���>Y���Ĥ��?�DS4���G�HD��s�����7O�Ο:%���y3@�gjLծ˩Q��ܗIK����7����?ly���]D�qB�Iށn��Ua��~˅p]���D�נ��G�)�8�%�/��i�KT�vñ���E�~�ԯ���]t�eI�u�5#$s��Q���B�#���@����ωWX$ySj�@\��0JݳJ�+�W�.f���m+=r櫎.�6�!��!�o���+�jI�g��4\�6���4C��B�9jE�a$?�s�E��gT�� W2�*�F�D)����^(Q��߀�%�	�*��ܣԄ\�-5�' >i"�,�Ŀ�3GV�S$2Ms��o�N��ツV��ml� O�<*���Y0��4�P�S�w�L;���)��£� H��es*ǟD�J�a7��3����F.#�Z�F�U�t�%�
2���C�`����o��