��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��*X*���-�M�����}i2H�r�t��+�ghl|�w��񑚧��$��E�p���
�V{]�/쐗�oBqh'k'�~��]
2k�V������x�1�Vbxo4�G�4\h
<� �1�
�`�
�D	\hl���u�	��~��Z��\�S��������~�x�P�kU\�-���+��GT�5�w�Q��}H
C�	'���8�T`y������K�F��ԓ*������0�� 
�����C�v��
�$9�Kƺ������/r|�����ɑc��JU;��-�� u�5���p���[ȓ	_�05S�1�Nׄ8�E�E����.ǟ�[�7&*с��(�
��2����>U�BDVj`�1#i0K�S�]>��61� �F�{���Ǜ����HSsr�j����[�kG>����s��N��&/�q�L���տ0���b�%HaG��}#�@�Q����\���)Bq��T��1/�:=�A��#@���? �����cTI�.����0�r�峵@;^��Er!}*��_��a��),'ơw\��py�/�2�P�_T���|	2�1�
�_pѠe<���¯�CJ���8I�����s��� ꡶&DM�5��|��+r>�]��u����Tv���$
	�~�'��?�w_���g8.�(�v�*w����h�~֥��(�4߆�pa�{Fd����Z6J	1��`���ڎ�&�hmI�_����`��7�`ǂ�����@��u�/��`�q��m���t_ʌ�ؤ_�Dr�H�G���&��M�ֳe�&*>a�X8��G	���aP閏��9 Q��[�_E�-P)uM'��^^5gưyI	_��{p�p�C7�g�� �����_�C8�(y3
E�j�PS(#�ۮ`Hť���T�={�2a�tI��3�;����
l2,+��ń�S2<8`��^'��AWӮJ*�;%�_9_*z
"�q����{�xb�����* ��ӵ!��^�j;tY�l$~�U�����4
��n���3e�@���$�%=�/�r�4�o}�|K�ʩ�����'xE�t�I���ɜ�|K�g��o�\��2����^b];����V�d����0�T�Q��M�Ʈ�lste��e@pCg�5�[��/�(��tSҗh��qGj<1|zd�Ro�@A�P聫�-���?�n���0R���=m��-�ʛ��O�8��1�>��?u��S)S��
5Y��&�J!����m��ա�{��2nU�3�^z�C�8QF����çz����g.�_i:�)����$��8}w�^��\�E����X�B� �6s^!�tK�0��LjU$P������fE�͗�����rR�ڂ���FQ+�n��j,7��)�!�o����8m��_��
���u' �zN�9q�nƃo/���} �p�[��l�m����c(oW�
�_�� /��n�Sa��+FR�c?xA$�d۬�r���w
͈�H��@Y�V`�e���X�����`�,X��s���5z����y�^	��B����hbrϝS����1�a�V/�n;�¹bQ�ګ:�؈K.��0� �� �h��0prU���+�� J:�d�2i��#��8J6�Ru��b����\D!U )������JTJ�@4����%����Z�9y�O��67��(W�@��*��)�kHB������Too��p�q*q���= sfc�&[n�;Z!��w���hV�˄A���֡�[;� �.nuR�����8�|��lq��ov^�U�I��3�.b�Õaz�=|T��M�_�̵�~iզ�o��ޡN�]�n�)�t�� ���7F��i}v��)u���l
^	��A���Ğ���@DMZ�!��-+ H�G{O΄��ۧ�����N�~����83k��$��6��,�d���Ӄ��X�KLi�AO@xQ�v������Gf��ɥ%_�T�p%u@��P�Bd���'%����P�%����f���̠�H
BiT`����?W������i�K�T� _�Y4�>`�{&�¡U���)4QbJqx�yo/���{��w-;ސR*��X��G�f=%��6n�0O������֚b�(�Φ���
	]w���E����(f��#ދ��8۷Uh9q����H}�c���+D��dV:kBʧ�2��<���̂pdJqb.H��OX�I]�`���7V�N�����{$~�]��ed熌������5䂩��;S�
-��&>a��V�;Ը'�����Wj7���3\����O����6�1\q�V�Y�ED@�p���9ꍍ���=yq92=�Z\��[Ѓ7�T#�rR�d�IH�4�� #h������Z��"�Wz9p���=؝_B�_�;��.�L�i���b 3Ĉ��f4��c�\�zB�G4��b�t[��� ^���;��3�����B,?��	�؋:I��&�zd�씨.�D P0T�/�U��+5��[
Tv1����'���ٻ����a���&�2�!)(yM�������o�A��eY ີ�~'��gY���א� ~u�fV��[
�ħںQ-P;�"�V�
���G4��p��Q�9m�آ(19)��	�I�?��^����ӹ�]$��rOLkzGչؿ�]j�#m�D��e�N��sAj;�cGJ��ͣ^����t�ö��&���r:�f/`ױ7��=���;F����kPR�2G�
	�C�Hn���)�~��K;^>���7�ғ�L��L���;�ɼ���Z�Cl���,2l���l�j�}^Vs!�ͪ+s���Xw�Q�8�vO')��+w�����X�K�ޥ�Py?��E�;F�܎r��%�Ɨ�d�j�hH�����d���w~ş�<N�ɳ�7$d�3��/��^?�ő�l�����?��*%����ɔM<X���Y얯#��-{F��(�Ĭz�d4a��O@]����!ኌ���t��n}$W���_^�(�,�e}$#�d�B\�mDOt��,.	��R�,�9�ʳ(��R?ǪC�&%=e���f��t��@� �OK��%��i�����A6��G��xezx��T���e5���f�U�����.b+([�fN����X�v-6�A�~��Or\'zU��g�����*:� �u|�����ҝ� aU�g)<��;|�	]��^����R.���5_�)#�n�����S&��p/�匲�m,��Ewg���h�<4ӫcZ]V[�JE��c��{���l�þ�zr4�������؉���(���J�W ���+�s�5(-H��f�x�Sy�G��+\Ɍf�u�lop�#r+� CŁMb�:
���Œ���˄T��R�R������$mmnR��5���W��/�(�aC��ok��K�+wT��h~�cB3�9�eQx�%g�rdO2~d�,_�!�i�Π֮���v5dM$����R8*9��r1 �����r�x<$�f70_�@�'Q�\,̿�y�3��"����B�:�^� Ŕ|�2��~N�<�����x�sK <���9���f�.6��F��up����[��Vu*[HJ��kO�Sz���J9?��Wj�5)�����驺o��6.�?zc��?-�:N:&ù��%��@��g͇�����C4k��{�'�>��{?i]��4&�>�,�H��V�LfU��k𘁬��v�{�����
q�x�#��D	Lۉ��#��x3;���+����o�Θ �%���)�~q;{��R�/9��si*Cu*�����Zw�%?�8�Q\��{��S�1��;���vytp\t���w"(H��Şq �,#S�L�O�u�qᏋ�챽�P��Q���(�IW~q�;���"⧸n"�p�2�w�ۼ}���ͽͬY0_d<u�Е��8��<��C��F,>㏒W�W�j��my�O,�<�Buo�M{,R�Vcޏ�mȹ�D~�ތv]1�Fr-;�D���Al�Y�\oP������(�e�sMj�h��(�|JĪ��`%Y����|"� >4L��j0��j
!�n�o�N~M�RW4�����{̈Ly~�I��dH��~ ���%2k��2�3�C������ч�*>�">����y�4�ad�; <RMMb�"�g�Vj�I_w��Kn�}i���? .":9���Z����
����k)��1n�ZP�ܶ�d��'�K;����Ϋ�3�ޜ���]�9����o�lg�'�:Z2��D�y�
~VlHe���fId�{�.L$�N�-�[��h	��~P��� ����Q?$��,�o@`��{����ڶ ����0��v����I�̓�t^	n>�g�}$��z\v���'�
�!Ԫͺm��@J��#Z�	>��+����A����|�a�T<r��d�^_��D��ڊ���J%'t�[��u5�l�L�����^��W���Y�>w�V�W��2M̢��&��N���Bգ|���Z�>��i���c�I�5�)'Q��D-�O��!I&P�uf��"�8�qH��G?�	)zg��<j�S%r���ܘ�m�R:Y��iD�¨�V�.��9DZ�H�yI��ն��Su��)vK���E�
��H+Xw��[��nmD�h�5GBy�<�Q�<�ԧ�'���3%��!�h��:���8���^�ե�hH0z����z �ӄ`�ƥ�
3 ;�jw(AO�ejΊ!��5.U~��<���焻�Y�c
�D�0BZ��9>�����$zÕ���g�t�����R��>*N�"���X5)j�y��cS�aG���@���xn��7�j2l��Y?Y�X!�]P?�b�#}�h�Fc������T��h��j_�l*x��>핽s��i^���+l��/��s��yi�	ze�Q�_���Ʌ��;����	��.)ܮ}pl`����!6a�,������!�Ic��o����!UBw����Z�A'A>��
�D%�96�%15� �}9!�5c*h��X��+m=k�P�m�Z�k{�9q�\A$i^�W�I��@y_�g�>�yp��83���[?����{W#����P!V���\<e�.OW[��{����·f3|��A<H��ݘ~��y�L��7�\Ik��(��>�R���,TM^D��eQ�����'�ΨS��be��Z�r����D�_e���c,�ȸAV1�?��c/L8�4�I6���*O�*�ش�U8�]D�xF���^4�$�+�+�g\q���B�|ƅ9^�Y,o�H����ʠŵ�9����fO�9o������B�Y$L��l|��RH;�M�Up<"��S���̏�AUӓ7E��?Q�����|�j/3Ľ��/�`��9
t���Z�R�b�z*��o�-�a�������45@�>�`�_t� Tv����ۛ��m��
�V��3dy�m�n�>�E�(&%$N&� �i�)���#���h	�� �`�����f�\�;=Px:*�Ai<(�����:��'ֈ�f��϶��$��K��"�OkWϸb���w�'�7��eNW�(��.ʄ�RM�4�w:_\zǧ�MY���li�|wRkI?�8NUXȜ�r����4��Cj���x�"�:7)�"�z�9tW\�A�sn+]Y~0n��&�W���Z��=�YIy[�:x��Fٵ���S��f�4g]I3!b��f�#�Z�-�wS@�t�6!���]mi}�60FhLK�`��������Q�ӻ�DhF����8�A�<W��(�Z�(�L�A�*���O5O� �$�2?�	��T���e�_c�6'�w�G��
�G��3��hm��s�,(_�?�fnX=�<=+4H ����M��GRމ��Ӱ�``�٭�]�],ay>�xOQ����}�,��د�������*Ʌ��;�8^�y����F&ׁ�A��5��k`��cDb�n�/�����`�^���)��P�	��"�>���Ď�&��!���A.538й���s�F�gW��j�"K�jC��@��}ڠKR���j&����������;?���Q?!�z�:�����*)H�F~^g�J.8ˎyswDj+���'�zp��Aw�$��$q~�3��2��]�B�R��cCt�D��K����iK�b*��Bg�W{&KZ�����K,=Y����$l�t����ch5��������ZQ��H9I���&U���{	o)���2V�)�$�^Z���v�e�*�i{�k)�&�w�[S"%r���{%����������r������*��
��>5$�}Rb򥐿�\�Q����~����l,[���ojk �)mAP�Z�Kv�z@G(Z��	����c���6��߷qp4�����4I��!!ux�w4���Riܣ���[]�^C'����t[��gx���_6��x�_�KT��^`�r~Ӧ;�(#8��j�+�	A|;D��o�-*�w�ƊJ~>��C!'�NA \�W�j�9s�u�ς^�bU�4�J������0gU� #����UV��n���D۰�o��6�9.����F14w��K����6�3����d��:i��7�x��o��!i�ؒϏ���ob��#�(E4�\�5?j��&��>�O��E�>r��)��sE���^߂����v�(��3Ү�9�0��\A�H`[�n������C�J)@�C_v_!髂�I���oH���U�?�ٰ�9��"�}�߭�	�i3�g�NOF�.�[��b����`���a�����o!�=�P��}K���?qd�U�b�K�w��V�<���.��@1�h�ͽ��@�Y�2ύ��(�ĺqO�������1����!_�N����*��W6�-�m95���r�g&��n���fwNhL1!Y���a�( ��1^JaD���/k }�x�-��^|dA?(\A3���5Q���eX�N�5j_{�O^Oq�"�ϒ�&���{�W��l�3ū���}\�ݖ�mLK\刾y��wz�~�4c�Ku����c�$1�S-53��V��"pqZ|��A��q��vЉ���U��D��وC��7�e��Tkp�Va��6~Z������9���C���I����� 1���#g0�i�ģ�����k55�8�=%������	�/�g�#45`~Y�?�[��M��S�(�ew�Hy_h����穬':�H�k�$���;����e��ÐwϤ_�o+X�Ā����NgH%�-�v@RS�� �p��	�EqOd��p�!AS^,oIl�w��J�5���t�
NQc��钬�ݞ,k��ù��IZ<_MdR3J6��������9�:@�p��퐥w����r>��uz^��ݟG��(�N�Lt'TДf�^�'VX	�c��T߱��%��]��|`�,&�B�J��2�m0w<\�=�����֗�� jh-7���k��j���9���V,X����d��W� G'�*ɉ��v�-���#0C�#&��aɥðNoE��._D��#�3i��9�����)EAǧ�RK����;�"�IkCh����J=�W���Ň騸r^����R����) �OC���Ĩ����j��ħ�������'Uj�����>N�'Ψ��kJ���:�{�ī��Xi�*��jEg���/w�	���ť��u}P����Ȝ�!��r5�m���B�8xQ��m�i�T}"h�WT�{W�7��?��:�Pn9���[�.=5��xǡ��%��j�Pm�8=��b�lXB�ܕ`"P\���`-��Zt�It��[��ث�D�j����q����r�_V��Z*�DR~�=�w$�%e
����1[�h����!X����,���P>K_t0e��g �:�AiD�U�w�\�ʉ�媨�	�����[���&}��ů8,�.��h�jݕ���$a�fu��HXz�ϴ	<9�
�%G����Z�#��U����p����P|�� �7��<8�塗Zu�b��}�FDq�>GD�h47,�	�0f�Ѣ��t{��T���[����]�Pk�+82+�ˎo�+�YA�jV،/�S^�$�n�،����h�1j���6Ί�\O��t9��m��s��*R��tl��w��9ƒ�!���SU��|�D�_@��US�m�(]��5{G�	���uP1�ƕ���������D�4I��*��Dz�+r|e@;%	0��_F#ő��p3���6o�j�K�����|���@�����w�W�<O����N�~�:�X���(3��-~��RjS���~�0|�˕<i��������ׯr�sC o�֝�0�w�7��"����jpP�d�
-~&r�l��6r�l=���Ҟ=��9��F�E����J#m`�����C��{�I�X�|� � �u��`��)��!��L�̟�v��O���MP.OcV״�O��8L#�t���Vz�ʆ�$RR�����H�;,uS勇�*�Q柳���p\������H�CW �Y�/�+��D�"[���S�**����	Ji�0v��DC"��8��8"�T��JP�@��F�����4t��`d�r�Ƭ�<�1]����*����� �x��*��{>d �A���*amx?8'.��K.�2���g%q#Mp��;��1�F��}���Z��gFbD0��׿���^�w���;�{��=W�p4��f�]�6���P�R;s�S=��|�:@*���͜ĉ���a�S�Ԉ}Ë�A*�{(垸�c�_��:�mI e��_��4^iUʲ��P�Atj)�Ş\ ���4`��b_��2~�lp�h~w���9���	3T�"��U���N�6Vc�U����E��XP4�A��������m�؁�h��!;Z��B���zn�C�>	2�w��9-�s����㿗/�+�#��o�a̶�7R�i�t<su-��"!�r�:9�� �	07���]��f���y��)f����?��w�Q���`����wҞh����Q�N�	h���E�z
�g��XO	�nV�
��	?�I.7���f/��$��Xh5�^�7�7�݄�R$��x�q%1e�"2�d#9Ou�,o�(��B'&A����(զ�M��ݰ۟w�1o4]��*����A_b�� �(��=V|>�e��������.J�!T�r:1<s��S��N�����ɿn8q��&��N�2���3�aD��4�Jm*��crW�|��s��ޛ��Kyt^;)S�^G3��G[��)X���:�`���,ג݌�*tmi�-u�U��f���xD0�-�-Iۯ��8��u�E��񦜏�;,<����Y�Z���`�`#�X8$!�+͠�]L����K����m@�[�� x�R������������-����IШa��U�χS@\S��l1�:�W��f
���Q�v&H���٨��J�;4�QpY���[�#b�MI(W�j���dq��і+��GS��W�g��
�t�c���ld�R�0?Ц�Z0���z���������ez�-�%�����Na%��ы��Q�wjѤ_�C�:/L�?C/G���C��D\<ܔ��J�dE�=v�t���RD�I[D�?���:�Pt����t��cRs�l֭cX��O5U[E�4�ۿ��.�+;������w)�R�f)e��U��}��/$5)�zX�R�.���,dL"�*p(�!wH
��S�Z��=���щY�:M�KK6��v='Y���@3�,0i��)���ǵ���dR��� �ٸ��x�!��)ǋ����1��Q<EcT�t�>�j���3�����.ظ�eq�!���ȯ=,��EC������.)q��خ��	1��9 ���z6	ڢF��~y��b<�����O���E��anz^��y9�M���;s4���;@�s3ą�ЀX K��0��书Z���?0���޵�_���X�������U��i�~.p��pgo���=�E���/%MM������ԊAKLS�#=����z��p��u:�T�ļ��?�X�)+����k�����D}�ɀJlq�����M�\q��]nC�$����E?�Q�d�:i���d8�S��+P��~X��*r��Fwq]��g˃e�Os}�X��+-U��{%\���QW��IQ%X���FM짿�h8���
���͎l*�l�w� ��to1qx�&�H�_��[�,e<$�5h%Vy#��Sk��Á����gȓ��	��˰4a��%}%Q�
��!�r�������@�>F��'����|8��H��+�!��^(�9�N��/�E!�%�{N��%�o[�/�	�_8뿂r�q�%d�u@�"ٴ�B?�����e��#�1	��uZ���1��x��ׄ�@�;r�g�]�"0}~��*��5��ҵ{t(���'ym��d����M��6��9�$I%����33Y�;D��/p#�nI=�Mߋ3p:��-İ��z���_P�
[�x���H�K&��������e�I����m-��S"[OW�,"�V�~�Zn�K2�.L��˾7�Ԍ��Z����8��1[񺪺�@�^C�9�6.F_���$/K5_!f�����FG�{�]��p�8?A���$(�cV(r��4��=.b|ܘ�}�$�^F��\��UTى�1��HY��>�IE �6�`nh�s�/�U�FP�ڇw7 ��ǹv�!쩯��@��B���q����_D��Y��>h�U�B�{wC��(Y&�kj�]%�sv�;�����V�uŁ���������e���k{��Ⱦ����w� �^]-�
�/��>bA!<�,�g4^�"�gb��{8i�6��W�*�	����^^
:r&H���R?$�ڇ{Z�A!��V�RB{��sK0��D'�H��^e��6�qmͭ�+��m.5��U�j�~g̉�o�mt���7�)oMDH
ﱱa�G�Y�/�P�-@_u���� Q"�R.:���wL��\̗8L�dɛ_~���Ш�DQr�i�b�M_�>�-����$IoO�x�	zB����Cj���+<٘��"��Au<��`W#��Ҳ� M���� �����q*��&N��׆@�BX��ؓ���*@�)���,�"�>Ps}֥�O����
�u ��J8�{�͹� ���g-��O�8tw+�3���?�\a?n����r}�g.H�<=�t(�����hM%�@�$^�������.�e|�\�2,��a��GX�irm&�W��%,E*A~G\�C2 ��PV�y�桽�4j�������%�q�t1�4h5i��v{Q��.��yT��Ҕ^��8���_35�D��u�-P2!:PV��=>�u �G��N���&ws��N��k�\��8��|R���#!��v�����st��u8��-�0�ѝ�_�WS,�O�ƀa�%qy�tz�mˡ���x+~�(�_����f�g�E�&���S_tgR�S�V�m�0�'=bW� ���˫B���O�߫��R����P��J�`�Kp/Lc�-��m�pM"��H�<7�gJ4�S\�>S`\Aי5�&E2V �5=�7l��I��~Pz����Rㇾ�I��?4�;��w;�L55_������x0z�������P c(r��w;qnf0��@B�!Np�{ݞ��X�÷)�c  l�5'�!�{�/י�I% _l*	�,�r�"�v��4�c�p���2���+�u"������l����J�b���WM\E�Y!�c?��ۋ(r���8�Qd^����|(}������ZK��i҂VG<��>�!X��GL�P��ʎ� %���K�1�������4����H��,Is����� ���ȝ@->F-�w�Лq5���Gɹ��&!m�1L�=�U{l����ى¨�A��`
�'Q�g���c��Mr}zXw�|Kf�ذ�Ic�?��`ȫ`b���-�{��3��~���$��G�(G�Sk�lC�{t]
�b��n�xm���:�Z���s¼���]����::��������t��H�=Iӑ��-���1ݙ��<�:���*G`px���\BYZ�� "�BlWr�_�)\E+�w��z�1��6!ɥ^N�V�e�5I�d-os>��"�䛳K,�G	w��Cy�?w>5)4��/�Bv��pMB
�k���r�|�����@2��r���jbw!5[�##���'���]��|Osc��^a$�
i2���z([+٬]�d�E餌&�VB_� N*�ۦ��~Y����9[JC��`����<�"�QP���}&��ߦ`V�p����%�XAXX�E |�c�a���$e��ź[ٶ��LP�g-�1��ϫ�q�$�^�3���ڲ�2���x��`0���}W�f#���n���a6.r�w�ïG0c�Al#ߚ����o�ſI��g><	�{�������� BXDn�b��P��J�#.���l����P	c��5�ܿ�+�~��#�K�44��{����͗⳩��7y!���d�-�pց-�	ݷn�i�KfaʧC�,�
)�8��1N=�	�^4ڥ�Z�KZ�����B�N�p\��� �Vp��H��)Xc=�@qo���m�n�7a�	Oq{ 
�n4�+���p�B���F j�nQɚy�D�啨�
�o���Q�`l���Fޠ7*�}�Nߥ#wKV��t�� �I��QUn�Iȕ��D!��0��v��),�!��.˄�8��T���伊h�P�!v�P��X��q�Փ�u�0r!�I�����;Շ��"�0bWVmf�����ʏ"��CXMWU���鸃�be���)H�J ��(���-��t�v�p���X@7�Vu$�b��B�Mu%J���x����# <���/@�UhL��*���P�]�1s �^p_0�<�P4��A�v��y��\M�kV�9!��L�l��,�H��$w���S�pƱvՈ����ɽ��HN��CW�ߓ��aNb?��:��[���Kξ�\fZɞͼ��@��K�L���ME�`��G(�F�w(����1�=�lLayx�b6�}���nabfAӭ��i,E�׸K����!���S���u���O�=��5�Ի�� �1Ci���h�,��3(j�F -z(��>;p��G�a/������I#��"�O�����bj�e�!�
����/���\���K}�_�U��LA��C�3]����=ƴ�\����� W��K1���k�3�c��.��L%�^��L�VI��5)'��(��MF7�äu3�aJ�2��TG����� R��:܄�x�yDJ��М�B�����<���g�4H�+����Q�Tb�O�7d�����~�!�&l��v#�=m��➔�笑��,�Qm��"�<}�p�Ee~����t֔�ߐ1^Xo����
"���`��E'��gм��ds�v�P��.���ҟ���z/t��9M���H��W�;�A�
�Q��<��C�$Z����{�7�S�W>P��@׉g��9�̌LF�"��.SA�����ӏ~H�8#�΃���������F���Ϩ�h�y4����i��U�acB������2f}��enק��Tj`{.��p�,Ʌ.d��f9/�rO�M%��k!`�ؙ�

8��+�#�������ͪ<�"���x�ߚ���R�n�16h8�����pZ���q��ǫ����I�#�j_�������C��9�(��@�?;�DS,����Z�s�F�
P�RD���\J�wH9�����sP�e���f.�ﴙ��x1�̪�d�1[������;77��y�4d�en3e�2Z�)�e���O7>�K 	-l�	W?N:}����̦��!ǚ����6�ˌ��@�t��m���K����* �:6��p�*�������v�5!���>�B�[m ���>H�tl�=%<��ڭ�!��������b;_���M��d�!B�J�� c��!����e�#�Ij䠞��%��	*<P�%��!�(P:/E�$M����e. Oy}��gZ�,���!pz� �"X��-�� � r`��>�V�.��42�QE�v %�aއ)�G���1w��}�%L� ���%}�Ol+x�ê[%ᤦF,-�K��?�+j;�C$p�����ucr��d�C�*�|��]Y�$�LW��vʫ�%r2@�@�s��������l)�(!i�Y���&�9�c�~�U[X<�=�d��5	��X�"%*����}�|�M��{:�b����3AC�xX�����������m�"��p�U�ف��sO+&��Nr��ً�a9�_W�z�~-صx}}��\ M�1��z�<�ڲ��������n��w�34��xBS��!��5�.��3�{��§��@���|��O�o23�r�DZj�&��}�@R�!xW�,�<Lo�w�����B��%_��gh2°☒�xx��M��Zn{�ϓ��\�/�8 u��oĨI�z�I�uԭ��h���<������(�q��������qk��U+MK/i�5(�p(s��%G�R2L�� 	Jܑ^�aӋ�\���k~pq��|�i�1_�)&Vo�T��zȤ���3�I�c����!ƃ��d����;?k5�:.�<�s�$���B�z5�y��*Ҹ$��ԝ�I�Ձ]m_`���J[�;@� ��7�mYW ��V���o![���)� �̻��7��E���6�E��}m�)m��.�!�V��� �	J�Y�&`�H�򵔠K�Q�բ<�AJ����G�T&�T|e�a�c��*�7�4��z�����u|��^S���,�a�y~����9�]LS£��F;��Z����#i��S�|o�X0��l�V��H�[�YY��s:�0��xF����fa]�LE]�/ع=tq����|�����&�9u�#�����i�W	����&fO%�����Z���{Qp��.�O�/x�v�ކ�8����2�	�G��YU�x�Ju9�I8�`��zNtD�;�_y�DW�$&\V�є�g>,H� ��	��ے�S�]�6I�T�zAx]���c������_A@J7�OC�LyA�`�� ��[��k��>e���nս�\"��6�B���WJa�n��>�<) �~2�u��.�A�͑)�\��cr?�}��Ld��Nݬ��x�@H&7��8�E��*o�h��7����ՅŉM��R�C����l_�oQ�T��3="�*u�ޗW���ݓ1���c>���&c��)��#����h��"���Tfy��	Ah�O2�>�4�V'��&+��^�gr٪���'}��u�X<�l�i?z� �%Uyl�&9�o�c��ݺ�#����ұ�ˏ Ď�j�L�$��X>.��U�w�qݱ{|��� ga�L9FV�ŏl3zSe!ϔ�K�-
d��6��+!e�B����vҖ�Hl�)�d� ��"Y�b `�$�'?�	0��q�7Å���W�
ͦ�p�Jo��W�·3�����E�+���%�����v������AlUF�����iE��oTສ����t\~PJ��x�9���! ?��l&J���/�_h�{Lq���1��
B��O��.l�kn��^��xPF�Ŕv�[�0�?�};6� �FF�ۆ���D-כ�uK����0R�d7/�I7JX�Hj��x8	&��RrS�J�d�$-�c��u�Nʻ�kQ5[�Z�-���W�t"��7��S�34j�~�}��?���聍�V�H�4+䋮�}�C�o���E���bX~&:{��3���s���q�b^����f����ږ���J� ��="�e�^�8u��Y��@$8{�h��S�]�Г�Ƿ޿��u�fM-f�.��'���n���(�S8cx�L{�΀��H����%�c:
7*Y�>>�u���'o���'0"���4v`H�3�AKY�f-��(�I����d� ��� ͷ=s���u�f�U!�L���=K�Y\kt�Z��hl^�Ex$�L�IX��3?�I�|{P��~��Ņ��k�Xy�����S��99�R��!���Y�;��w��i������h�-���t�)t6�8Oi^�����J=��z}/�z������8� ���0~72L0R� r��-�����Trff��g1m��a~��Q��9bi3Ӹ}�a����j����G��r��&x��*�mCz�a3f�ly�)�Fr!��%��"9}{�C{�3i6�����`��D�F�TE�N;K�@
ʉ�u�a�,Km' ���K�Gn�"E��Ńߎ �\Lӣ0a1T���+��U��BĐ��RR�#�8_����F�QeHR{n]{N`��ο ���d���Z8)��s8C���t9�[�{UM�@rVBp`r�&�Q@�Q+̫1H��o�Ԧ��=LP)i8Yi��K�xЄ����W]{��26� U�j�ʂw~Ò3L������0
�7	�x�;�FJ�e:�g93���?��8��wY V@G���&G�i�>~:["��ɫ}b�	��I�4�ކ/g�Lk��;���R^��끇��~q���׶=e&f,�	l;����XC6�g����ow�t:]��&��8 � �V���jc:�3:Z�����'�w�vj�5=l��{��>鱼��.[n��W�_d����+��WU``sd!;Pc�;��Q�6[Rz��%Y�๒ zg�N���!�'�/(�?V-�@<���i0w���j��L(ߏ����#g��m,�Fsr A��ie�Kђ�-�ֶ�L8�ٌN�{	�J��)�۱$���LdJ�IL�ңΉ	��Ȓ�
8NY�2g�'�B>��1��A�%*��2�~�.�'@�-Z�F��E>m ���B�N&������4��]<ؘnP�l
�����[��{)�$j,x��)N48k���ׂC�'	r�/����O1�50�f�@�;_U����~F���V�5�Tvc��ֱ��hN�
����y��I��gT dd}�'�$yY��W�lẀ��c�	�1���3���})�b�^+8��35,z�g���_�B�K�˞6�a"�Kd߇C6�L�Ok�j�?�F+V3/��3�;��^�����R�DX~bY�"���+b/H3���EV�)���i�i�,���J�e{�[��c^ѴB�v��O��i&�ʡZ� pW�0<%z�Θ5#���!�w¡> �/�`r���*o�hl�����nm�-�ui�IÓ�Ɯ�ԡs'x�|P�� ˮ&���RD�P����>]��v��!��� q���)C�NqhTV��m�!�Tn��-��R�}���N�,~����+�R�MO���wiC�m�┪�G�Ýv5l�i�+�S�x�@r�t�n~�G��u�1bs~�=���3bݺ̑k�B`�&�/��n����J���}i��;�X�G��}�ƼC<NOOQ'c:.O*���Tڲ%�;��.o4�}�p[e5�i�	%.�5l��ƻ��>�iZ��=�G��)�������f�Q;����XV��EV\��9vk�nJ���"��Fْ�i>�P�Mrd�!Reb�l ���w~��Ro;�kj�
M����{������!3
�*��������F�n�(�j�trG�������;� o���o�X��� ��9�{�1�c���Ǵ ����\����@�}���( �� ~�x�z���+�	lzV��s�-��c-��y�R�p5�;7�G�b��=����F���]H�8)�6�L%G��dS4#��wGj:�I����m�$��#���RY�xL�?62י�,�`m��P���� ����B�+><�0�3I�Re<n���y�������f�̥/��^����<��IP,�p?�ض�J���/�򒥙˦3�q�Fӎq=5�o coH�ؚ �ǉ<B���If��������l��h�KwafN}�"�4��@�f��~�Z���s�ߢcW���\_J(P66:H+�?�Q#*k����╨Y3V�
��i�#+p9��@��.L��zO�w����ۺIn6��eא}tj�
��@>��p��=<�+���ӭ��.���������R�R�T�8y�pw���f�F�A�43b���PnfP��Maw}R��SY��A�ہ�� ��@v�Mܲ�O!���~�I+0��%��k��˟����L}BZ��/Vm��WY�X�W���U�(�',�zM�>�%�f��]v��"
�|�!��Gj�+����f�x9���<��{�����x�����`�o&�U�<_�>��O4h�)�t6Pl-���f��=�Saв��p�OOa�s\�Kȗ���J<�I����n�r��`j�- �E���G��1��`�pJ9�-���y.(��U�XE�����uڧ�>Τd�'�޳#�R�/��R� #�r�@^L�nf��??�|Z� �����j���ɋәJv���Vt��TrЉIO�ݎP~����H��CH���+���y������nc�j�l[~,�;��(SH�����!&�/�$��)?[�����Vj-�$=�a�i�Zf�)���Zm�yw�-r>/E�3�I!P���g}su�F�D�����uL�C�B�3Xq�*���17��n���3eg2O �Y���F� u_�S:c�(��G�P��m���s@1B~�\ZI�z�zt���%��"���qe:B��eht�\0�����N=�9?���6X�Sna��8�;(�ݝE_�x`�uZ}y�@P��xO���_Y��e���T����CV�ə��2���d؋.z=���]�Z�vC?9gP�'����B����ɤJ|�@⌡#�У�O���"bE����h� \F���f[����~��9'�*�bX��U�����'N��D+�91 X��\�)ƃ;�H�B=��b#('=�N�	�5������q[ɰ��z�l{�	U�5*9>a������cޜ.��;0���Oc4��;���V;`ȁ	y1�����y?�̏�∑�ׇ��E�o����+I�,=���E�4$��S!���D鈎Ge�A-��ւm�����^(7���S�gJ��;H����W�(�d}�x��EgX��q?$���y��doN�����B�X_�uM��lui�(/kQ�*�hx�ގ�K�۾	PҾ$Ӵ�/�P�N��Z�-r��U�B3)���g�ވ��N|{��Z�Ía�@2f�B���%G\�у#$"]���ȴ������L��1P`��U�-��m��ͯ��!hѣ�a����I�]~��h�n���N+�����V�8ב��&��gq��2�E����&�Z�-����ػ����1f�|��~���'�XнLj̉��Zb�K�YEW�U�
}!r I��͐�(*q���0��)�}��>�ef���0[�3�˦��O�-��.��a�X���!�q;�c��i��(��_�F'��4�~jt��DT��2���	.��ߔ�'h��<)��D���]��e�xnɿ�z
�I��s/!��㧀@L��,�J��>�H���n): ��M�*Y��I{��Qч�I�K˒WAI���4���D��-������� o(��\{V�w�d��nX}N~�w+Di�Gi-���BT'2����!�+�:	�T'�yKS�,}sv{����1�a�-�@Q�!L�委�ij���/>¶����f6�Rc� �D�sjl~�Z���v�KjdU��6�5��o�O��s�q,"�h6���S����+b��'�E纭*�E��JCz��E���o��%2l:l]M$N_$��DO�D��ڗ����C�x�#�>�~�^�dk��"�	�B��*h��77����-c�.^H�M5}��)�G�1 �w >ez���F����N$X-��la���Ɠ��zDSAႨ@�����d&��Y��)$ks#�B��	V�X���Q����8'ק��rE�	ɲ�&��ћ����3ٟ��X�SS�<֩���CWE����oN\vNoD�D9�I�H�I^C����d@4хy�:��_խ㟠.K�npP�簀��S@l��&Q�>��ߢ���k.v���6��6���J��sW�T���#��'_��OYW�XK��=��$��C �����b�Y6��sgn���C�1H����1�2=㮀���ޝ�̋>���9��t������^C�g�Ed&7�����U����g���њ���P�w��ٱ&j&��>���� r�[��%6��g3a!���H��~�ew��(~pt�����L::��|m�@
E�}�-<F�����߶�D4� ~�.Ȱ��+n��	}���������KuK)*��z��T��9�.���G�cp��;�^w�F�8�m��x��id�������ԛ�|Y�����<�.�vXS��GR@p�v����/�X\��^��{�3�&��1+���-��0��:"��D����v_���(��w�b�����H�v)�Rk��5��1"�]����v	�����yf�»�|����:��(D��$�͜ .��E���e��,a���Ws�A��,�1Sj�!g��-�h'IV�["ܟ��?9������׊!�X���7��pʿ�$~y@��o���/N�j�/��ęw��p=(h�Qv3~�ݤ�^�_R![|��Bs����={�~GW{��/@LR�W�XȤ�3nb^���yg`�fQjl�qǀXy�������N����Zʍ�d�d~�CD��t'l"��`���^t�S�g~�C��}���(��Z�GP��6����sĐ5/j"��ԯU�x�h�0��N�p2U�~��f�E���+?!(xur?)<��u��m_CKЈ�}6 ���a���c���fذ����P�h�.T��w�6�e��ʓ�l�
��I�\�ѫ8�):}S�z�a�T"��}�5��uK�v�GJI�;~���I��y��夋� 0�K�.�"ۊ�vH*���A��p���Y)7(���uG$m	�4i��Ѝ�=���5P�υ���Z�"���7��yw(k�\ �V�vA���z�d/���B�]s�ݠ����Ӓ��/i������?q�hZ�������C@���#�W�zQ����Ag�*�y��fm�}"�cuG�.S��!'/+(o�Z�TX�����\�!R/rC��E����͢�td���r����m	J��T�5���u��d)iZ)1���5�s��/���n�1 J����&	�D�䏷g��1�����#�Ì�"
�f��CKX稄�(g$�^i�:�K��n��M�q?�pW^~7������V���t�������ki_�-��z���F�G�C���
Q$ݯ��ϖ�Bg���e�=��p:������*^��z0Ǭ���ކrQ��|т�iZua����6F�P6��8� pw!%�v�Z�z�넮���	�V��*�^���?h�A:0��3�j�a��}3���_�!�, wj��
gHv�_�0�\h{S��D�|���<ΙVv4��2�	 �\YK|G�"fw"p��zѵv� ��7�(���*qjVdF�@����R�N$;b��}�T�g�%�IMpom�'�M��`3��uCN���q���{�~��Ƭ� 	s���s6,P��V�nKK7i�� HTT�G �¢��ւiI�}K��1/�'�Iٳ�}W�yi7��U �
3ީ�bN��Q,���7���Pq^p�id;��ߏDݸ/y�v@�"��9�.l��ɣM��%Pqmc��c58�����`�~tz$��%�{���"m�krL�"L�$+(K,>p4��{��m��#@?��"��k�Wi�^�3Y����&Gp�m��d8��P�̢ɞ�΄���͖=x2�A��[`�* ��� ��5;v<���]�lM�n�6,*7:�x�%�*8���#����2�Z�X4(W��UW�όp3+�S�%�^�:�KMqyE
�o�վ ������ ��%�������#L%�<��������NE3,Үt�t{e��	>�6=���������>|��܄2����0�y<ǂ#�� W����v���ެ<���[�﹊խ�Wm;Dc艸o�ryՒv@05.�w��B���H�S9�6��
����I���+޸.`q�*��m�J��|/�:ܞh��������w�%S��0���UPM�������$��$K�>z�cj< �n��P�-�\A�!D?u���� @�}}u���ߊ:nuY;oU�S5�oX��b�	��M��݄h�*1|l�a^��$}c'B�8יo�<,9�̅��/DVa=�u�n�S�&��ӫH�O.�C�lw+��ģ%y*xZ;��c�)��~�넽7��D�ϲ�"�b��c#�Y��q��l�:���D�|�����k���]�+�:D���K\���%ܫ����SFT��S�$�{�ܺ^��İ�$���I�Gj�~̻Ѥ�{_-.�B?z���>�	[�����¶dGQhz�<
�.���_��n���]waI��w&Q���T�$�P9�
�ɻ�FL��R�~6����J8�.�j �WFR���/U� ��T0ә���]��dw��i�8Ը�ĳ)�^�NQ�
�c�.����-t	�r ��ن;�q'��reQ�\QԽ����O���RFӣ@�Ӫ�1�0$Jδ��z]�(nT�[��aa�y���;��{쮿�p9ILDU�ǻ�ݯ���E���i_���&ef��[N*�~�����*���[mV�Q�Rk��>@�9>�y!/1��b�7��:��ɽ��8P85?��ܝ�s3y�Kc��%�Ь�G���a�Ci�PO�؀gv���e[�����&罃��S�_s�6pa ���A���lj������[dbZ�� ��gڢ��)���H�{�\���X�ݯ�OJ�_޹�9�3en0+��j�$�����dJE�㞎1}@Ɖ�g1N��)�6ҋ0�3�������Οt��/�\�s�M�!�퀁��R�o}��@�P�<��e�D�G[QvB�S��oǽ+�?�Ȭ�r�gЃ,�%d��������-��(�W�H����L��"�b89h�(�.�G��x±T_��AǄ#�8�QIsK6ۂ6�������0�1�":�f�����f3�@2P��_9I|-�w�E\����|�����D��O*�bP`���Jt�u�7[Қ�Ge���-e]wP)nq3s���g��|�{Q�с=��v���h���j�I;,��~���H90���8riM��G?W���錺S5���1B ���mE�T�����T:�������\q&�6��.7�.�|�U�ڃ�� �oY���s9�9G���lL^����/��z�򙨆Y_N1}^��v	�c ��؞��b��HRߤ��q}�{���=��)i_�|��t�r���7꿎w�L�x�J�@���(���7����A-i�ciX����\�rh�4��_�����~U���h� � �H���Nj�_r/I'�k���l�
����eP�T�S/��㢳��l��V"��팵�Ck�e��8���d]�G?���J���&g]��
���,�������W�y�L��1��I�	=�Q�6�!�\�Z��	'�w4�SwM�,���|��oh (���ll�-�sW��"�mLf����{�F� �,���݀ )gXz�D����߂h���?�A�!1K�e_��	�̂�3d��˅0JКh�XqLhrź	��`L�^�}�$0t�����jv�oo���.eu=Q���^x"�[����Y.����8��K\�=\���z��ww�j�ݐ�4OG�:���a~y0,�7�Te%պ�+7W�,�zQ"S�?)��?�{���ٱ����T���lm+px9��F�(MAY�~�B�B���6���ȎN��BG9JI��+o�.x�b[���z���3f�L��E��P�C ���M(��K��ߑ�ۤ[��Z6�$�Ⓝ쓴���љ+���L��&d�:ȔQ\z�[��D�tg�K:_��GLE"��Y�s�:Z�Z{���
@S%*B�kh�t��%G��-MLBK�qdh�ǹ��?`W����rhs��Y��8������X-��-�г��4��)�&"�Jq�PQ��d+k�����R�����W֛@�۬������n�~�8�����1`��X�jS�K�h�f���I��Y�m4�$Ia}���Tv�`�e�FN�y�ՠn������SH'�Q|��t��&������
=rBU�	��t��8���-o�[���ɳU��":�������9/&q]�mW��-�%��,�r�)� \��@����
CuX�'�� T�g���Bt�w�~q��Q�G��Pƞ��	�󩞋Y.�{�n��v�|,���"�S���M��M�Yf��k��ӄݍ~ ����ԍ�=��u(��Y�K-�uQ�