��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�6��y�̘8-�����h�lYY;h<r ��(�ק�-4�~��RX�D�����a���1����U���K2_��~�K�K�;�!BvɃ�ZA�]�Ozܳ��ũ�# W�c�/&__���;�k�,���(i����vz9�֬��-���D{Φ8��N[�Wuɢڰ��>��	`��XU<����JF7m����
�����2���z]��T��.5mQ28M��!�<e������������?,'Yb!�7s`����|`V��'1q@�K�=�Z6��5�N5�p�0�5)�dI��Q2���l�_g <�?����狳bt�Z_��U�*D,�4��>F+��k�q��@�1U^7���d`Q�t�C�ӥ�r�rQf�s��������,�r�4@�RI�ȣ.P�q-圾���X���O},x���41��,��٭�8���� 	aGE)|]l�ڀX�;'VKu����f��n�J�~$6�V�L�z�n�ك��q��ch�3L$b/I�q�`?o}�

q�;�E�u�_\�������H5xC܆9);���-._�!�k�+g���6\�[;0b)U�=�C�ʠ͢��|'�i1��C�m�Q7�O�`D�8�3QĭZOs��֥�6P�Ч.,9d	x9��jܹ�x�������?�����c��^��
�������p5�F\�cB3pݫ��X�{]L����q7׵ ���b<B툋"P�셒Lr�q�ӏQ����0S�<6i�� �g��	�u��[Tb�qH�k��1���Kxdmɍ�7���{�x�`� ��\�Dr���� *IO���FF��$Ǳ���G��4�C�9T�ږ��"�Z�&tY5�ټX}�8���aDAS��lɪ��+@1zS~�#�s�2���l�A>Hr%z�⻽���oH�����З�����\L[i��Ѽ�ڨd���������D%}#G�����D!�z2���K�66�d����塮��\u%�_���Ea�C���F�G\�����ٛD�&E5�֋�k����U�̅��|���[$��:a+��ch�fT����Ñ8�=`}����6B�$C�<q8�� #xH>�0���+��ӹ�!;�A�Ja���]�h�qR'Z���`�A��K�Df5�3��v\�%+�8��Ms�24v�6��X��r|O�Un�IZZ��a��yp���t,:�A�OE��W�!�?ۖE����X||������(knf�فw��`����3��Nkv�]�E��X�(���0��.q�p,��h5����r���,���ھ�>��r��&�p`^�Y`����z�B�bT鬻�N�j�"!��n�\�v�`��o����|�/��(OS�o�xe��[�jr����Hǀ��렚�����d�aFk�HT���K�w	�tH��0�+@�.>�k �:�`|j�>InHqҿ��Zt]Y�qR;�š�hR	M����/f���g�M!�=�L�����E��{u���"��>}���
<+"������"�M�,�/? >�}���;1f.��5�+�v@}�U�-�l��&�1�pn��o6mڣ���ώ�� 	N+y��)��P��<9`a��&�=Mi�Y�S��-Q.�p��չ,�GBp��̥�<;>�(�(���ak��`�7��A�kk3�sf�C�ֳ�(��-��v�Xs;|E���#�,{���᫡e�~(e�AF���e�9�|�S�Xͣ�5�H%{I�aP쿑�Y�Q�w�D0zib��|YY��l�Dn�j�s-���/��KP�a�>�����(��v�J�c�$�������R�(�><cI�i���n#��;{1��ef^���U�F�����R�Լ ��6���<���D�NǠ��5�K{B�?�,S���)=r3��k�8�����!�����S}7<u^�b�/��|�K���V��L�A��*g�$���Z�<Hm!�(���L��	AY��9�s1o N=���������^��v߱k�ɖe *_a�N�tC���l�u�?�|����߲�lǘ/k�F#)����`<�]#j�z�Yܠ��T�P��t���TUR��l��PCm/GIy�*�lD�?�
5��0��5�%C.8�� c�޵��`�����(c�]��!�V�f�5	|6�@�����Rϼ3�<Kw�ˍ�P.�L��������μV�mkӉ�&���H��
��'�[�s�^ٷ_ˊ�ug���}�d�>1v�BX$��sIzЅ�7�$���b1b"EW���_��Rw�vz�>46	�;��GE���.G��G��pG�*����gJ���t�_�E'Lc`�h�8�I�����}�6������/It?��h����#� �,�L<�w�di[�g��T��+E:z�;��+�p�[�1�Ȧ�m���-U��h��(uyE�gؙ17U����J[s��a ����'z��Y��}.�ZMi\E3�<���4%L���ٝ���L���/m.�B\"��k����Fm�
#�}!����[�����Is��?F�2C��P,&'�~v���:��(Zk��s'K���9w9�XmG{��5�����d��3I��ɲ��Ɗv+�N��z)u�G��+��}YV�j�"e
���乇�n{;���lo��f:⬎/+�L®1�m�7yQm�n������J�Tw8ϝ��bGՀ��"�IG�R��S����ZR J�I��u���aEܣ�.&	Ъ񮆪��1K��]�C�Q��!'�A*5�gX�>��-�M9u��ڨ�m�כGlk���Rkq_�aʽ�Fx'0����:)��!�$�m�\�i�i��+ן[��\��фL�L�j����	��7r���0��(�M�Qb�G�T��5�g��Jy:&~��Opd@紬�GX�J��ݴ��bn���s�vm��9��[/,u}�6"0T\ax�}?�'2�\��c���D�Tx�uA�JO�=*�:#۞C'�_�_�	�ѥ�a�Ҽ ��]X�l�Jt��w��$�\�+ �Ko��U�ŶP4��;Z��!'7�[��£�\�O.œ%^�.�[;�ɺ�w�甑	ǐ}�G��A�!o� �P*۲K���(��茅� h���*�$�	�	p]8B���8��7��?�kgA�A�YP(��YG�Ҋ�~b�EB^�~�(��8D�l�����'�O��

b��.6|G��g�����Y_7"���5��v՞��U�qK�Ia0���Ƣ�t�۹����K��ֈ<���C\��~��6[�Z6l��9��s\��3ط���><���p0��1Q}�`�l@VF���W�������OV��Ug��*�*]q#'En���גw\i^0	��`�0��eZ}���
��0�r�|�f�� ���u@d�="X��b�u*_�	l�q�u�F.Z�uޞ�Z�W�@Ik��S�a!|1i�\z2_%�+�w���a�y��0^�q D֑�e�_�'n������M��.1�i��_I%V�9��/ ��I�w�]%9�2�O4_��;�E /̀��S)X-�a@U'�c4�.`�2B�I�q;�締�f�y��oH�q2�Ny K=�P�G�tR�X�5D��)�E�;""�`�˭A�����?��h-�f�<��$��q;y��t��W�?����g����������M���-hL�:�������q8N������1U�~�b(n��w+��X�$��jU��x�%iZ��. �eIs%��`�{߾�[��UGw�ޱqt�Nu��>c �$q����p��sS���q��1�)��v�7����E�]oɓ��1Q���]s��Z6'`��g�Ɖ�qdяK�CĒ��wv.��)���S_�&�p>�����}�6�Y&"��9�]�:�<� `��"�)/�p4�0l��������)��57샢E$[q~6-�w�7[�f.p,���)�S�b�����I�$f�e�G�OS���W9���y׺5�^LA�BY���L�s/�۶dnܮ8�6[w�]>�uK[��\��PnV�Np�3�����]>]gGM��pCH��z�`+��>Dm�酠�PQ���9x3����wJ\�bP
���<�|6��`��u/��;ն
e��6�qC`�U�l��Sw]	-pl��?#�N�s!�͇��y$t���� �8�j�
�ʡߊuD��BTGE�I����q2�F��G��l+,��l1L\�cW�!nPġ;*��Kk�@�O��dJ�,��V�t�,Lx���^��ۡ����@��8[;�0��H���V�!>�u�RFE�/�RY)�#X�|��d/���Ul�/�qP1�Q�S��*�x
,���-��ڣ����6��W>���!X��F�z������,JS�]�g����9����d�vLԱ.S��fU��g��N���r��i�Í�x�Io�L)����tĿR���$l�زKT���XB�mQ� �4<{��i=�Ԇ�¸]������j۔̡�!^%�����/6:A�U󃰶_#�L�E�̠-d%R�p�����jO��f�_���iw�ƅ���H��L'��99 �D;k�� ?Y���f9��[Qk�9��C�/�����h�詛 4_��˩�P�B�g���'e���8��%�d �:z7��N �p���� ��̸�B�����/ �nu��y��n�WW�Z]H<W(�����#�]Z<�Oٲ;r�o�����B��k1iϠm��&U#��U`�lp�y��0N�	r`Ӕ̱o�{#m�CW��.�4�>�N��
¼�p鈪�wW��#$J.�G��G��{����<0_���uƘ���
�v�L�j�.o_��P�/��ƹ�Ɉ���_0Bԅ?i�79"3jC޾�������e�[]U�/C�}VDs;�%�}�:)yg~��0��t2�~�F�㲽/�xd*���������ޔm�>����S?�F��4����\�j.���!�\���V)��x�����%$�5�7Ib �;�"l����7~n��UF����ꑑO"̶QM�j�ʎ����$y9]F�v�ٔ�L�zx��UF�CV��G�9o��>D.���J�j_��2͓�2߷E�-����&�����3ֽ%ձ�r�R�P�w��Os	�ߝ|�X%�>@�E�2��^���)����NA��z/�K�-x�y��
b]�OXR�[�@"�Šx$R�w����s����d�%�j#�BآM�d8Wy��7p\�6�m�(͈�Ҥ<�01�Pa?�L� j�2W�-�e�kࡖe�w�%}���/Kl˥(+>�k1�=��7.(��­�uK��m��\w��=s���H�D�f0��:���e�r��y��Tѧ��r�	
�3�S�L2sx��+ ��?Xܨ�)[�D���"�Âgn�y� ,�價���S?#y�P�u��l9�W�#pw��������l��K�:Yj�us�չojrj�d�L������������쐅�+�E{�d���"�x[_C n�X��2�V�U�̘�US�JU���em0�����T0=\����Pze���f.,j�*��0����7��s�եa7�R��cbQ�~�i���(����U�����R�U����80�*F&����z����i�Xɪ%V���IHѭ���;�_�������Fn���>3��}KC��gv�Gd�|w�r)���A!�P��TX����^&i��h�v�k؍v"��'��VT�h��'����/sX�}���h�F:�+L�d����%�,�h/��l���sb�оҹ~���j8e/�@�z�R�!Z�Rn7*�*T��u�UW9�C�g*X��ժ�&t[�<�Ia�S��m%���%6��ɋ1��T���{x��K��5��&�f������9�d0\��'�
0�����<��Ȑcs?gv��_���6Vi7*�v���w׊."`��!�w	-���ki�7j8�����j�P �x�3������hV7���L���D���6�I�j{�4���`����B���V�,g9 I�F<h#�yQ��H�D"�x[A]�13��f�9�V��a�����&�(U�qƛ�%�y�"�t����ƫ��P��<mn�Kŧ:��'1D��)�t���1d��{�V�o����r������Ww��:�gӦ���bdO�&��-�
,����L��3JT	7p1ժD���q	-�ޚ�� ���Q.�"���:C$�^��6i�^^<��<C>8� �61��]��{�b2?�<&�Fũ۫CЕ�7� �v�b3����;N��+�Z'��Z�8�nN�FK�|쪛ǁe7)eɠ�*834��Ø�n
W�����r��?�x�eh�up�cO�z��BQ�������Z�$��e%j��U����r�+�=�}�Z�]�2چ�&7(�A�hHX��0�Uy�Έ�o�-���[\㤆;�������vf$�FOt!��&r�1��r���IK*`'��jᡄ�QIV�%��zpV��-0���P
2c�=��
�p}�aN}��)0��\�y���҂��s���ؕV:��}�����hCy��}�3�Ѐ��4��^�(�l$	���d��i�ţ��/�B{h� �Wj��#�ǂ��~H�������i6.'J!��B�E�
�L��Z-��=u4k���'I}���
��ΐ}�k�Rn2V��Fm֧PPmC	�H�_RA+�? ��_�	[{�{��Y$�'���a'�^<�t���@^�����
𐓊؅\ʠ���[}����q�&r��Y��C�x �~ˎю-xW ⴱ�i��_�d�;���7��=����f�9�����{�&�^��y�����}����O�gS��o_�� �n���#]���kbG�'��wu
c�C.O5��r��az��IKkPa) O�&�`ˊ�t��J&4i�x��P�R3��X!ZA��gE^�x~�w5�2�m�����A�'ݪ?�NY�z�zZ�	�ӵ�Ɠ����H� �2���۶1etZ�*� 2$u�m������ޡ��Ζ;�~�h���I�KY�(��4F�#ۃ��z+��iձ�p/P��߷}��_E�2����+�b���ph��))4Fp:^k3��R�_�vX�]D��nβY)�<[�5�Y�)&�f�.7��ק1?�4���9��`F����{�瑋� +h��k:���Nr"7�#1ѣ�竌�N�(��D�����$��:�`M�S�G�����iF�c?_����S�F#
�X���fއ�5T7ｉG�RH��s�����r�tb 8d`�64M/5�R�}���2���c����%(;�ł
�bg�@P̟ײ��,R�$��cܫ��j5���)w���
Z��B4rj��Ǟ����k1�@5�[����O���uAiǯ�3�Z�.��E�HSc�jH\�|�o�TN
-�g�go�B�}*�c�r�l��m�,[k���62�J�x]�):V(?1xgv+�IS�k����Y�Ƭ	Ŗ%�:G�'�!I�#���9�B�6�<����<��GX��+?���!���xZۦH���VE�����I	�S4ѫ$�L7�j^H'|�d{%P� "%�˺�܎|�'%��m��P0Y����.x�Z-�9sL��_%֞)]/'Y���o5����@r�!��<���S�zG3��)f� 'C8��� �X����H���6}%�x��vu���;I�ϻ籧�OI����O�NE�/���{KW�!����
��UP����𦣋 �G��xa��߃�?0eo�vP�J��!����"��ί�x����.C�eɞ὇Vz8�T�j� �g���Q�䍸��9f͕9#FPa�j��{mg]�������:x����%���1���$\.n�S�������#Ф�"���T�8 ��~cG+�S5��I���V�:w@t|�mf�, R
��W��T4]��M/pL8��\^�H7u/7C�ʊ����� ���%D��*T�z�X�|5ñ�dW+���a��gI��1>��F�����9Dq[����I�;D������.dS�s�:����+�C��]Uu�c>5P��I�km+�z�1���FH�ʫ��M�	h�ծ�K�Ab�����h�����9x��Ϲ��8�I Cg�ᦉ"X�#s��'��&x$����H)aE#%[���g2:׿.3a5|#�j�?9�5�byM��ub�?�+�w~ν�����ĳ�������M�+�#d�0�O���qF���&�vf3�:����k�QE@k�ҩ_d 1F��Ԇ*��Elt�Wk�n�}��;�����1����y����*�M�^�Qh?�.��z?moq%}r�'ɟ� ��%]�+[<�x�A��*�8�fB�>6{D��I{*�?��vVF��a!?jI����i�g2��?у�ӫZ����E$l��ݡ�� Ⱥ��5Sq�:���`��6��+��7�D@���X�,d�9�`�^ӽU���oؗ�
t������n��g=��6�~&Ί2�"p)\�3;�$� ��!������l�Sz1A���Ew�8�-?78-�9��p����8ɣ����N�!��P�x �K����}�T$���Y5�G���x!]����L%�\���:cAxV��O �j�
ؗҷ��?��֓)\�����8�j��`@��v��F$1OqU��4�Ȍ��p���l	�*�AC����v��'X�B�9���*�c�Ww�S��ܝV�{2%a��ٯ�;�ɺ�ahv�V��D]q���h_�\/G�?�H@@88�l'Ҳx�C1�M�	���,������y���%*�w��-i����ڇ�q2���ZH8�썍?c��)�a��.+�|�~clcZ��}�j�ڈ���(1����CW5*�`��x�y��th0�4	����w���_|�/���%�+��(ч��Zy��	B���$o������ ����G2mdzi�J|.���{A:R�l5"���=4���;<{�x���hHP�%�ou����m�ԏS�E�V��Y�P<���`�8� c͕8f�?�.ް�`텁�B����v얆	�շ�I.v��ډ��r.�S�osSnA��A��� �'�%�(9Ȭ��7d��5'V����y�A�U��(3��|;�����G�\T.mYf���鶣[jCޖ*JҕuID�j�	X�r<O����j+��nļ�(� ȡɱD⠟��gf�,�+��Y#����=��~�Ia��X��MS�E�D��2p�b(����l;
����G'��L��\�v������1Qw�9Ca�Vʲ�ڧH����WE���#Oh�-��$��K��9H�n��pn��+��=�rO���c�Ne�|�TQ0�C�R-��g"�Z���\��Xnb�	�����==uNM�E`�b`��ޔh�F���/���R_mέw��_�j�?��;'�R؊���ys�(���g�ܦ��QA����[n����V�h`K4K���g��х�.���;@�Y0��n�R���^PQ n�	6>��gd����"�jܼ���5��GO�<������츾-���C�*B�ڥ�{P�����g�4�75D��x�xR��L�q���f�2f?s�,9�l�H�c��,B5���
LwRL���8��x�9p���00c�|a0%���㹟��i����Py"�Kw	��h�^����nǰle�n�8ݦy���<���
5�NK�L.,��&GoRp��!�I��Z��Q�بI��bB`�ݮ �ȅx$��T��t�Б��vu���.&r�	�uO�O�NU�{���ʢ�1��@�9js�B��p�$��-@�u`�@�jdb��v�����C`��ټU��4��2��滄.f��
w
�?�s�H�k`,������XU�󦭏�`4�v���A}7�$�q��y�f�mK�4�e�:|��l4�0���>�}��bj�9�氪��ʚ�fד�&��ȘJ�d��u�\�U�b͌6wn���	�)�$&[�Mz��֭�3�Ym����1dM[�P\k�xr`������
U?��3-.(�N��{�j�R�&�Ƶ5�f�k&�D^l�:�oB��L�3�>�������q}Fk?F��Uw��DE�7]Ї�gꙁ�j�A�^Ý�&H�H\7�P��-�,�k�8�=�gj%*����)T��K��㟓��0p�K~,a�FNruy	��L6uŕ�O��[�"z��9����r��%5�6�1�/��,�.k&��Α|�I�b�ݬ��&�2���W>g#��V�予!U�4�)�A�O-GԚ�������CZ]�I65�~V-b��Q� �T$�t��2xS�"P�j���{�>�%u\������+v���Y��kJ7�O�h��Xj#����j��w����L5Z\|^�"��XoPF���q��G�4��^/�E�1�����?#���N�[���=I읏�IRB�k}7r�-�(EyPMp�W�Ҋ� c�'��n�ۢi�� �ة��U��p��$N�
�c����J���� �q�`�����h �����~�EփuE�8���&�_�ɑ��'O( �� ͦ��V(n��=�Щ₽���hw|r�~^��" �i��߄@����Dи-�)�[�df��Sq��5X�g5>9�It=�;����'j� ��[A��%����f��O�bа��T�����˚(�/����O����-��},!��@:r�${g^�<�Y_6A!���q�Q��K?",Eʋ�E;�ܘG�zj��
Y����G�'mE}�4iFV���-���^�߀�-�b��Is�MKZti�Y��+�l�	;$`3�2��n�y��^Ƿp�)���Z��=�_�V3dN��ܷw;�t�R[���q��*��MU��Fzi(�i<��b��k�
���+��l�1|bfFO;���(>șI��<�r�Rx�����%b]s�ma's��c+Α��VY>��K��,~y~�PQ�� ����������I\�A�<c��k(�Wh�þ��*��^+Ѝ4Xo��IL�r	��㒾��<Gt���ztPv�}��E� \��~qۇ5��lG P���0*����o���6N�9�������r�s�M�=����rjz�����c�D����?vr���"��g��nQlp@ɮ4
���rN��A%��:��x��:�!�>[�G�w1���8.�DG�⫎1y 	�=�=e���כ �ʺ�K;7@K2��	vw��(��ua��kG)��h�r8bs��|�?"�(��� #fA�2�=tq�p`cjy~��=����j��Z�3��d�<�8��nK�~�K,�8c��v
��uJx�.����eV},��_�
��nUc�ec�u�5�x֣2���r�@���}��:> 'Ѣ�84�ivjb�}�|�7g���6��?����¤�C��g	�o����{L]�8:T��K�<!?yPM%d |�v��>����j�f�>� �SN|d͟��3����0���p��r���2(F�U��ٳW�%�l}Zǈ-��t>��_�t1�{z�q��y�9l�#�t�R4RX5y�-O�A��~�ï�VT2�!2!�_u�C���"a|���X�z�����Q�k}y�͑,��.
'ho>z��Is���%�v6d�P�����7����7�=�Q􌝯�SKi�<���#ɇ��5�i�u�,�q�%?�@䤔�^kew}�" h�x�;���t2 pr�$�>,�5��r��@u���z��A�����w��q��+YF˩B�&c�[�=G���	��i��;s� �:$u��8z�0g�F h�FD��n�"(+.��51~�^Ped�Y��j��?���o���Jܧ���f�L�vE�[R2�-)Y��rw4��Y�B����0$
�+#a0g�J�,�ѦF��@��ʨЃ"�]��9�"6L� ��Y(�<�Y����N2�,��C2C���j��������j�e����L�p_�>���Vv��t^�+�)R�F�p(?�ePLPR�%m�pyE� ��PF�v��JF�a������7����6�A�kC��s�է�e��	uh=�WK�����Q�6�Si��&}����V	�q;��֏ш�e+�C�Ә'��\���R�Y
���`����ցz����1p��T���¿4����QOq6l��6꧄�y��O����]��.C�-����h�WzzF]f<6,l���6&h�$F�%F�d5ᘅV,���bub��4[��+�;��1�z��B݆w=��-C,;��ĥB�I�X�y�U�u���prLǨ�j������4��[�Ybw����v��4�>�A�o���"�"���WU�V{��(=S�7�7T�4�p��)fM�����JKV��'ـ*�������o�}�.�FD�W��z%�>���+���F�ďe�ۓ9)IZ���6��{?:�z���]��m#�a�����[}r�3�PN�x�|Q��j3q�q��G���ԥ�N�g!{5�&�^R�.�W�`�M���������ϫ���ˎ�D�A���{d�|� ,�8K�u�B[� �lx>��J��\`�d�o8��m�:�nʊ]G�fG��T�Ġ-p)/�?�a���H��&R/��> ܞ�/���M#�Y_�W�)����ӑ� �)ƭ�9o�p]���+�D�/beZR*@2���0��!kM����Ę�C�g�����
���R>Ds�i����r�Lqe����r�	�s|�L�p}���Jwc��x����y�FV�|M@Õ�4��]�P��$��Y�z���"�LyAQ�bkں ���g�o�x|N UI�^�z�=
n?��h�����̴������!��XHM6�+��?�&�1J���\�@
�DD��d��F��|)d�{��8�8���N?��ɰ�]���K��:�)� �Z��������qP[g_��UU��P�k�T+�s�f�N�ϧ�R롛-�j������D���;vm%[��C�����%T�dJs�wv��P�ڙ"��P��������"Ky]��)f�L�9W讪/8`��V@"v^��p�š�"�{`��ڄP2�7�[s�]�/���W��n�������F]�l�jsntb{�o#\���4��P��7�.��B�I�	���+�⎞[=ڮW�\d�gN��YD�է(8gw��cq�����ۢ�8;6��-W�oZ�С{���/p,�mR�����%�O��&Ęt��{�$ӧ$h�峃��wyȤ��"�U��L5�W8�N��7
���0���z�EV ��]���f�,i@�I�qM���P+&l�}�Mqg��ġ��b�"a'#�#a����f8b����v�Z~R�x �[�kRk�Չ6\C��B�=vQI��8gL�㋓�ΈE,���<Ug���A�E}���l���Hc6�c��G��L�k̢�a{�u=�a��c8�>�����,��wN�brCY����.�'�f�����g��veSՑ�;!������' ��tU�k�<q�S��YxD��=f|�!�e��Y�0,�ap��U(�#󕹂�"��X����n����`~z�E��rU�;x�0�ۯ0�ߑϕ�����y���@�wۯꕛrR(};ݵ���1K��@�#\�鮬N�1�	*B����1���3l�C���z�H|*�A+��+��NҦGP�HIҳ�Œ�$���"�J��{R�!����
��q�s�������aJe��'g|K!��V����t�BBV�"�fy;U�/6K�Ƴ�Mڹ����pz*=�S�8�~�����sW�k73��)F�N�bf�8�Q��� D%89SQ��Gu���C�sn������ ��l�Ơ�U�����u���`�N�ZE�E{z����9��4s��]��� �Q&���编�������p,C�f@�s~��΀�߼F>*��D;�Ջ�G��&�|��r�!$8�X|O*l�0���Z�� ����00-�n[kpo(G�Ntj�!`�Dam���o~϶�W�`.)u�4���&�G�6#�7X8ޟm2%",�PeV����͇�r������Ҡ�����X���.6֤�-��p����%!=}:�eA5�O���5���*5n��c�{nնg��hb�8�M'�Rz\q�y{�� ͗�C��/\'�4����0��?L���v3k� �k�r�}4��Կ�zs�z(X�����E��5���UO�BL�z?�����[���}��Fb/kL�^�
�́�-���U��G�V4��[}ܨ-tjÑ���
>����D7��/b�:�k��:�����K���c�g�"k�mF]�~�|���V�� b�p��$"u�z Y����n�7e+]��h[��k���Ҭ���5)�Y���J~�I�+қ�E^�uHinbi����ڷR�je��ة�g>�F�`g�Ig�2�5aC���L�1�̔���.�$&�v��ѝ��yv������+F��?j�k�B�z��m��T��]n�u%G9�M��t�#~���e�(<)��N�%��b�ц��߀K��۪�^�3��SZz� �m�%ψ��-��^��hLU,��n��2¥����i�: ln�؞�1��#��#T*+X�^rX�N)�	x-N�f*!�.h�:��@-:e�t���8��N�^�DB�n�Fa�ֻ��ɖ���О��f�^Λ�������5�a�BΆ+ǽ�<�0���-��_4(�(>�u)�eǤ�Ks�
��Y�b9�m��8��y��}�U���H�u���Ӗ���M}��v����6�wY23T.{˽ �d�����A�vț'�sĕ�H�-�jN��Ɋ�t���hiA%��L��/�\�� />�f��~!�T�]X��)uNp��7���O� ��S=��ط��L\��qL㕍����+9 ok,�x�������\�~��M�P��������N��0�����R����|?��|�������m1�~.��iC���=���� �cu�`��G�6J��6%p��7#;>|����t�*��!���zl��S�`�~q��s�WJ��9��I���Yr��-oR�y�Jř�یgl)�"�a�����oZ�wW����{�i�9�������9��E��'B+2���S��"�_P
	4��u&/
q��p����jQ��ehB�K����ԓ_1��/h׶�A����
�|ߎ7�{��$�s���e� ��k�����Ŕ�o��A7�.|��Ua����˃~�H8�BIS1/L���ɕgZ�c$�}��}-?U0�(Aj�A�_�}�3�t\�+���4�q*�XQH���+[n�?�������G�J]�g�y��]����v�o��$�����&	r�Vb �U�h���#�y���E��t�=�_�^��{��ȭ��O�Z��J�@�M��7��lC(l�l�{͈��oL�Þ�*���5q��U�bA.6�1�6S�2b&(�����z���T,�s�t�JCY�ƿL��M^�S;�*��>^aM��RN��<���p\lZ��:;�i�3�4�(tb�o��r��]L�����L�h��h@}���P
����!@�U�����4���Ė�uBT�`�i��'K����;_�8#=��w��K�-e�m�+k�p�Z�^>^`�p��&��	%���2����?�*���6t�GUqq�3#�B��׋�8��f����Ućc����ץMt햆�tb@�!sL)����\׸ME�A'1�ւ�̰���P[�E���Z;�U�gz&Q���tӔy��Z��a9�ᓁ��*gx�eӔ���w;ϙ��V��?��쭷������9�z�0|N1�n|��ziR��Ѥ:> �aG:��a3v}{?lA��^�?A(�b�g���%����4�ԱjJ��#������kd��n�Jc���,�L �{�K��p&*�[����<��Ħ}""{�*S�h�?�`��
��
��y�;�=�A��-��L講N�Ц��q����F�R��s�S��Д�.LK�9ckIP$�Fb�K	��^	�� i���i(�$5�q�s;f���ϱn�Rk��1�ƅW,�В����(g��0k�T �(��E�I~0#�8�D{��2RX��^������E@�n��j����Kt��/j��e��Ǡ?�FH�H�˜=L�d��=�&4B�`�`�#����KJ�|f�AR�gj0�釟G��$kL�=KC��ٺ��|buJ����d	d�{3�k�"Gך�~>�q��Z�U��KR�)�� ����� \������?�S�"���s֧E5D\Ar��(B�ʀ_pʀ`���,���fTt뉂!H�[�����e+Z`���a ���u�������
�"
���׉M1�z;P�y��_�B��j*�G�M�mJ�p����a�������+%����F:ȗI��d0���\â�J;=�3��U�t`��	0����jo^��͡�	�]t����>�}����u~�3���H�N�gX�X����_�*3��I�������H�����9�hd � ��<�E|"%���N$�UJ��	�6�h�_x1s���:����0 �t��ͽ��X��_�:f�Z^���/,����f�D�Y~P�cR�,
���f.��K�O�m�k��݊�/�=�R��N�<3ཀv���x���� w��sk�:,MІ����-¥�v�pp�C��/TB&E��d�:�L�j��nB>�t���}p�V�����H��<�4?��W����س����T�T�����.hQ��l&�/��y�G���؇�������3�`��=�B�lY�#f��~�C���$�!F�7&˴`Q���=ۧ�rW؁!O$�[Ai�jl��|�<p?æ�:'���͵�v߁I��������m㍭�#����ȝ��=#2{��T�w����1����HZ^����\q�qi�M��z䀤�e�
o�˗�?B��5�-d� ��"�t����O��Psj�D�b�L��e�E_pO���*�V��mEbHM�Q��͞�l�M��C�
=�Qxb���,X��w�0��Z�+Yl�0�E����m�J;Ŧڟ"^�LI��U����JQ�J��f��Er�i����9���40 �[�́Y�@�̂��Њj3~)��>����r��C�%���݃�Z ����%u��F�6�����Ȓ`	�l��ۭ#p�sH��ݖ�s5�x?��e�ģ�Η����e[�������g�as�2����2��0���b�&Tl����3x���sD���Dq�� �������`�g+/��Uq���b�.�����q��I��!�N^�/�h�͌������]_Bb��ar��2��R~�B�{� !�
,�	���'l�d�dU� ������hC{��->�c�
$-����l͝B��V�����j7-{s���G�*����Ez��l�����s݃�B={;%�A56Cz��Ĕc�@�vp���O�c�\�ʝ���R[����/�Z>��
�dB���|�_.s�7��]�6ɕ%�DR���	��B��1�լ�b86��D͘[�uh%�r���B8�F����4��Y1X�����j�f��f��1���Vo-��9���4�jbR �*�M����W()��[�"���l>�6 $_��W5<ޯ�Yfû��	��.}i�����GO�X\�/5�VUkҘ�F�뺟���⢊��振�;�aaCQ��B�[�Ir=4���\a���+y��X!�]!�{y�s��i#�I��Yi'�J����{��3 Ҹ07'�-��%��M_%ܢ�A��� 8�a�.]��jY����YWE(���:�[h{S��:;��gnX�k���h!
)˂@d���/���A�+�hؒ���֒6a��	@�����xy�h�?ɓ�م�P����܊�L��dC+Y�K�mf~%v���o���>2���?�i{���P���Ji��]Fڱ%OMe���~�;pVd���1�m�:w��P�g~!��m@y�u��lq�h,�9�[�o�!!�b�f��߳�F?QѨvە��8&y�+X��G�H�c����S1�a����#4��.�b�1<E��]����Yœ��������GjE��dJ��@C�R�m����5)_��u3��>��������k{AP
����8��^�v$�^�>+C�����Yb��o����F���_�z�h�h�x!ʚ�}��P �Ϋ���-J_YP��T��'w��Ώ��.O4�a�kT��ײ����6a�v���Z��u^5B/*���/n�AHc���L�HU��� �o3w�`���In�e���@mʏl}x@`A���l��A�u\�W�!M���:,�Gk���'5��S -��>��۝�{@s0^T�/��������T��j�VLK�@���=��o'3NB+^﹞�x~�>�;�1$ò��k�ϰ��ѭGy��\l��]�mV��Y�1[�C��+K�K��O- �Ƙջ�N�SJ�:��ܰjm~⋤��fД&�Z�g«��|&{��*��� �۠'G�Ȥ��ǋ�s��7^p)a��AR��$K�='w8n矙���'>k��o��7kP�yvG�C����C��sQ#��;�����<V��E��]%����@��Uۿ�x��ط�V�q��Y��>��p��S�z�)!b����5�ߵ����8��KI��`�є��9U̮�t'4�a��Ф|�������(�$%hn=���mt��l|1d�.M��B1yu�8QT��z���7u�v�Vu����A1_`�'c�}�E�08�JV�$ع���ZuK���Ϋ�<Fh�9�[
�"L+:q����Ib���̓j�C�̼2y����N>�΄_]U��v�e�d}��8U���%l�k��x�-��u|*aV���9�N�c�1IN8G:�]"X���(H!�ʝr�]pq�[ɣ�N�98Hv��r���VS��޷����#��b�%�P�Pu�e�(���*�ԭ
j��3��僤��`Du�;�&Y�%�٭_���M|<hLP�����Pi�>��c��YՍ�+;���0�Rp�{jy`( �6��M�I����ۼ����r�y@�_8%�\�|/3��b�{���ŕ��	��
`�ǾAS�������xMdUK�`�;���[XѷѲ���8�w�[��+.$=��CWaa�p� 9���v�����r�&G֝����3�k���<MD�A���A�nN�N��X�\5M���"��H����Md�^m���ȱ��1:(Ы�V���E!G�`i�����p���-X���;׀=�X�;4rP)}�l��FF��sUD/2	3����EkЉ�ҝ���A�����N'WN�Ⱥ�9*��t��*{�C�RW��#��rEyb��b93t��k�,�a��Y���-�aR�܆�i�!��8/5�`���J��b�⠞q�o��%N��4p��~B5ik���%x��sub8�Jok�j���k����hPLI/�)�"��A��By���Gȅ���S��$}4���{����ۙ�"j4C
|e��t3��L�ۧ\�Ì��^��%)>OjvP��h��_�6<� �O���4�Gx��H�+{	�U.X�ܺ�vY|���M���EO1��˂�S�SGq��d��z�ǒ�0G��*2lܓԚ�Mp�����:���v����c'7�|*ksjGG5c?P�ۺ6��%�t��z�UUe�Q�3�"%9Ka�v`,c~ᶕ���Yi7��>N{�h�i�;�Ww���hYT��<��	
����0�{�0��ӕH��c¸�ʞ9�k �ع��6x�q������O

��&���\��.�J^=*k܊7:@�O��� � 7�«p��kߎ>�	$f��T2���:-�����;x�а<^��V݌4K���df.����9f��������>�nS��CL]RѴ2x0�FZ��,X�T?j�l�b&ST�Ԫ�̉,?vw(�[����3�@U������0b��"k@�ZN�X�9���TA��}�ȾPD����&�4oe	�־�ępb�����V��ȹ�P+�*r`�o�u�f�+�5� ��Zy��ՙ�|F��I�C#V��k�z\�ܣ/J��ۈk�[��<b)4�FOcH�*��A;�:ACI����(,U��I[�RC�q�#��汅~<r��(P��ݨ�3����5z�1��O|�b ��H���4��d>���_��`^�N_;���T�_ϡ$������R�>�`J=�l�j^�N�υX�QR>�h3�����T6S�^_J�:=�{4,��̮�D%8ھa��"%?���/"WX��>:����
�����ƪKCYyMJ�E�y�����veۉ���)=�3��r��5|F��j.q;ȸ�أ�6h�'L�VwC����
��Mܼb�]�-� +f&�J��~z]�9˶�{s�D�El[}���Z���t\�k�u�/ ��.��oz��V������[��v�.*�������@�DJC�� {f���#9�h�$>���'�0��"|���w��w�_ުj@�/Sl3�o�2�>/���[i ��w���o:û����W��cu4������&�����h|y$.R��j50�AE��1�7���d��_Q�L!�����(V�������K���1��s0Ul6?��Q�ӊ%[,�r��|>��Gt��ޭ�S��ntĶJ�wh�6��y#��e�+۔Eag����9�V,j�_Q�N��&x��i/@�y㘡�պ��h(�	=�GH,rZdj� �?'u�$�wآd�ȑ�Zc6�;%D(�ӕ�}m̺�
t-��4[P���0%�x˻:h@E�z�s�%K@�*�9̂�B(Bٻ�Ћ��r���ŤL�)��.���?�Xk]J�&C2����_�g΀\�h�1��vu�Z���9 �tl�!NJu�Zv7N
�`Q8ّ��?��;\bS���TeY%[�άBk���J�5��B���W����$��M��9'@,���Mׁ��a0L��'�aQ�Uq��vꠌ�Y_*����]?\e���v�f��6���8���^��`gF�_1�Ă?�6�Ct��E����.��^�oq�/�и�Z-�k�����SM%S�xX��I��6>�Q�6(�bf���:�����r-:0�C��fr��p����s��^����
V;:���D�4���i�M������/w�t�_QC�_�>���5gP�8 �8M%�_m�-�;��u�����PPqSsb��<_��ڛ�=v�	��ܙ`y�#��M���Dj��E~kLP-��K�s��h�3����?f
��/���lR֙M+�*t�G��Ǻpy)�Z��#�n����"#?�9��c������T9�{l�vd��%�p]���������$/c}mjUwD�#�,oh��"ʵ��g���bοG��	smq��Q|_���]�\_���u����1�o��f"�f�*�)E.[�x9^��5��<D�F+���H*��s02��ӄ[^��D���V��K�~]::ȏs�h�^Z�т�C0�O�o�,_엽�L������Ss� �!1�D}�T3W��z�o�
b�����̰��-d?��M!��;��*�[��y�	[E�#20p~5cuG+j����Ѳ��R�!���3��(#Yty�)pY�An��?%��,]6�Z�b�,��U-���FC�7�h�(Lڨ^�c@L�B�i��,1����JB�g�qw�Ԋ	�/6��L@vx^q7b�V#vfӵ�e>l�R�JD�J�R7 ܞ��� 	�vQ��q s��������f���'3��9Yô�D�A� R4oY�+F	�9�N9A�������A��b1r�	�2�y��dW�:�P�i/iv{�=;���#_�8z�O���N�m ���w�G���pJ��؏7h?�X��)ߔY�N�����6�zfQ*�� ���cȠ���;` U�	T��DI\c�Wn�o����Z��!C��5r3�bTB<a�M"g�b��m�D'C��(N��D��#@[ϖ�
J��'	���G�5����g�(�#I����M�8���� :n�bV���c`�T��5�
��a��g p&��w_� n+j]�p	h1$e_G�d�\�7�*�`�b��1��!��͓�6PZe	��-�7��彟cƿ�XP���-�P�B� -���Ċ��t��pT��3�N˰Őkt���5� ��}�&L# N7�P�y�#�k	����?�Q�4�H�Z�h�2����-}���A�)S1e�V4P��M�-��_f=1	�����0� ���\��T ��i�l�t��)F���7�z�@v��,ɐ�V��)�c����(9yb��$/���F�px\b�]�q�h�}��N���ݖ	�DQF�L�l��9ݔ��x�sn���H���������f��������M�1��K�(�>�D�1�M��d򍢖�͊�="���i������}�;�}��~�'=�S���\�f�����v�=�xJ:��	�H�.��] ���񏬋�^ŧ6DT*V�h��G����//��E�r ~5o̳�)t��O�W�M�Y�7r� `�!6�u���;�8B��;P.E:����%Ð�3a��FM.""�!��wt!	�c���& ^�;S���2z�C"��t&�l����TPK��|�}�c�����~l̼� �^�B^����(0���I^2v��?r��KbA�jqKA[,���v�G���2K��3 ���3��$�Q�ʄ���{�Ф����i�q�Q�e�xB�EM�S�p�y�_�1�}jn`��dw�� �������q������h�	�E(Z9��$.1?�r*+ŋA��s���k%�$b�9Iҝ���A"��c7-���D6yn��#��''��������\�^�x�N^��#��w������Ys$#��.l�����_�f#���L���Q��:� 5q��J��J�zI��*�C��c�D4ϐ�Q|p}�X\���sPc�<T� _3If�#L�׊+�0:��r=R]���#H��u)��n��x�Yy�`6L�_�:����H����y�+��\r��<�Gj�����Spse��<�h�Ӥ�3"z�oJo���0z/�7�0�8��j;AгO�A�i��"�̞���ιF��&VvV��5N�v^��\(�¾��o�"ʜ�̺�>3�P���t}d/�	e�q��� ����ރ��p�W{�r��Vb*��/D��Ro����a��½۬���g����B� ��';��C�L�C�⾏�Rf�ˏ�"�Q\�����0V�Be�f��$�2K���6%�quu���0s�&w�(�/�5��w�@�1
1h�2%�@����+�X;�7� H�G*h��Җ���k�h���w���Me�y�uL���jrM	���ɰњ��B�zK���C����r�7{s6G�y��6e7�V oY�F?��Q�:+�1�Ų@Z_A�>��;L��Q���Yzo����*�"=?�^1�s@�[���ބ��6��s�ZF�9��.<q�4������F-pH��C��œ�>�����-Rv��Xp��@R[@��M�ܶ��ބ4�Ƹ6��F;�;�qҞ8�εD��6Ϲ�Uo_D�V1Ny]x���~����԰^�\:j��V�^S�xAs̑`����x�(���"���lV< �C#����5���6|��(��-��샟_�3%Ǿ�6~
��l��c�?�w)��Kg��	��BcF�@w��x$���r�z����ҕ��j<}�e����{PŽ
N��9_�|i�c	�Iv�5����¦ %�L����~��m}d����}�?>��oi�:���'��A�8^�d-Y~���l�Έc���ؐ�]��M�5n(��zO���g�J����x�R|�CT+�	U
���Ox/I���u��ET.ń�&�n�MUȄ�;˲�+�#&5�pE��K�B�S9�4�q-��?��Vhq��O����I'�����ے�d�ܢe�ʠD�Z*2ٳȵ��Bȼ���{�t>G�G���5��j�vQD~��I;z3A�D��8�	��7�<�a��(;��R6���p,Pֆ��u
uV*�S��.��z��X
�D��������R}D gA� ��-"���Vÿ}��,i��r�	$`�?Q�%�Q3���:�j�VXz��T'��˂�'ך8���$�3 �b�\�su�W<�!I@GXr3=j;����c�_��@e��\�r��<��}��a���֨�$����7-�_S����S~	�s�I��8o/D�"�k�ڊ@� 2�;����E�&��Bv]r��W|Jm����z�m�7�xd������3�nj���c�\�g=( & ���z���P���u������H���dQ)��9�v�>������Δt�d���sk�8�S��bf���[��k$�����G�Ua;F4φ��M��! ����mu��JǊ}g����_��K�N�����x��X�W�z�3$�l�=ph���w`�6f\{*{���QNs�Y|�����cK�'kΫ�	�{A3R���AFɗ'�R���3Ԑw�߳+G�f����P΀T�=�#� *�-�F�r@ 29���bŴ
h���'*-����͗@x�-B��g	?�Or1mf����RĜc��mj��Y���.v�etO��/J�2�h��B��.��=��%>y�ϝ�m.��f����^d}sK�p/h�a��QHf3��;_I�3g�*Rv.+�]"�Sh�`��tȩx��|
�2(?F�x�_�����=��.\T-B`!�������G��ⁱ@ONZ�ɗ �V���i���~�q@��sm�C
�2�ci���#�h�&,���NIpf �	�C���;!��1�!o+!���q4���fdM��+?�����2�SI��"�6�6bьm6��)�{Id^�/��#S�Z��*eﱟ �l�t.�����.\�Q�I�e�G�5�H�++oYK7�?���e�����@ MI������ h.J.����*���sj���!��� 4��bz�U��Pb80�R�c	�:��q������7ȉ�d��К�{aj��Bk�`�*�ӹ�sJ��QSJ�k7��K��jf<��\�X]����UzL��U��\]E�G�,!��XWf4�N��%�c���M{�L�~���ݸ�/���v���Sc��ܭ�q����qr�2���C?cv�Z�j��S��]H�g2iތ[
����E�>��Q1�5����yY�i�cI,������c+V��G�@�L�"ЇƑm	� ��\�2�_:�%������FV߱��A���`��(�}7��^�ͬad��h����Unp�rZ�7� �!g#"����q�K��i=�ۆ�!Ry��{!�N��5Pgd��΅:QN �#�� 0F@��c�9���3��擬��[RM�5�,Qt�_[��v��=얈Gk �_��b��}��I^�8<�J;�
C�T�pD�y��J��Ry�{K��Ecp�z��}Q�ih2:��U"_���׬b�)�Š���<��
`��5������'�q_�����X���1��p�=Y�%�hPho>S\�vߪQ�����f�Ē]8��u�^g@�g�R<)B����M	�NѺ��9�pj��w�BCEJ"�PQ�_���Z��\:�kz�$J;"O��m�s���S��a�y��۽�Eo0�W+�>-�b;�Iw��kp	;���dq�i�ߣrQ?�]�2=*���������Wt?Ub��Z#���JHy�}6�7�{��Y��w�	=�C�;��I�nޣ]���8徑}dSo:c�t��z����f�YO�'Yl-"����xv��34�U��	B��T���,�$%��
�x��o^p�Kȓ$�v(��`�i8J��,�m���9�|�򏺃2�0�4���p�5�1L��)h� �
C��GG��=��Þ�/_��^Cޗ�$e�*��B(��i^���a����Dy�9�~�r}۰�}ꕺ��Vcޙ"����(W:3�ʹ�~e�K&��~ׂx�<ѭ������`������NHL��P�l}�P[)����$��,�-�T�ap`�Z:�I�@^�FPm`}�2@�zz��=��ۢ��dJ��G	�jh�%L���k}-a��R�'�p�n���M5SZ1�H��oq����� ��+�T:w'���Q��+��,�ܨ��ZW{���Gy�)x˝�n�����*�goV�mb���;e��)<�!�d�˿�}�x�x�t�Ȟ_H��f����=<Xfy��q ��*5D�����������,�9X�� �垊-pc�߷��$�:�N���E�v�޼�fh�ִ��4J<eW]#�U�r�t��{�KmQZ���r5����'��g����*YY��}�)+r��"��HR���Sd�<B�n1=�(F�	�d�v�Q�`�y���eluU�?��	>�G�3m��l�`�1�O�ۗ�ZfvA�<�c��>�8(=dV�j��1�G?ϋh2�nWfI���g�	�.�m�F�gd�i�E��)8UE�9��F&�
f�#��B�>�E5\քO�4��)tq��D��D>A��ލfA�D��'�� �sO����ڴ�Qt��m@�N0!�	M�YZ`��1�W||D(�����^�V���s�'WUq�Q�n5�5r*c	V�b	>�!�pP����_�h�y?�\�O�k%^c��[��.����bnpΖ�o,9�B<ۢ�琸隺�t�}�y���S�� M��9g�����NA�
a8�M�cٗ����p���,�H6� ��}{�Rs\�ls�%��m�ڏq<��-G	&��`��Ϟ��//���ߨ<�z%8�!��e�W6��:�@����{�����Xyg$���{}q�J��J��k��hr�X@ƿ�:�kϰ�|�n1DQ8�?��ѩ�s�4�]�9ܑ�T���ٍ⼝�a�2���:���7ZI�lX�UU���N��<�6"3�W��*Z7��i�f�jڃ|^�B�*��6Y�����H�n�KWű�գ߂6#�-�@�
'���A����y����bF/a��/�
�ݔ1e���8�!z����,ꕬ	%��:�p��\Y��̜��ڦ��@���vZ�YW��],k�(������(�$���al�>�̣#�Mf�5�$���m+�A�����k�=1ƀ^��\�3��{��c��k䏀��n�?!*4�4 +6���7,�sP�50��OR��qRd��H��"�h���x�Cu4�%f�!�i�("�
QR�����ds�)������S*�xXj�(�ͮ���NĐ=�A��wx��S��|�9?�<8�%v�y	٫�3�ɡI���e)q�C�F�#4��q4�v�I6��X�!=;(ZW��I>�5!E.م��;6:���I/LqH��j���鶾f�B�h�)��^すQ���{ɢ�p�uf�vM�5�iF#
��ȝ��@�7ʉ���Tb�𑕬u�J�z3�/؀�7d�/��n}{��(/�҅��o��9���.�3�iq7����>2�ؒ.�Jڨ�|�����Α��6���*��eB��
��gwy�:�ܷ��������j7M�"��#����ݓT>4�$H�}�����a�����L���/�� �	�	���GA3�dm�5M�ylCV���5��Ӕ>j*	$4��"�H�dč`D��+���/�r-\��\;Y���^rp�r�!����SY�&/��-a� �U���,�1g�����/��g].�\�$���p��Ga� ����LRqJ�׋�c�0�)�&�>n��a�'���ab�a½���Y�e��y�T���;S�N���{3vL�����O�9�-5{�X��)�;��tC�W��s�r�oɄ;� �.����V����k�)?�渤l[�T	��J�R��m�;��DAx	\��9�j��9�k�P�J�aD�U��l�ɀcR��Q�ń�>(���{x�s����'Mƛ� ��#�}|5���L�4b!�t��5Xq�ZG��S��&� N+�����̥-�s�z��O`��g�.Ű6&���Y�AB���lBO�w���F�m 7���צ�G����#Z�=h.�R�yf��}��H<dr8�)�Mjq�6��I� ��c���U�q1�M�~�D��h��OQ��]���S@�&�ʒ����E9�/�)�YrA�o���!��p���L�x��4\�e�.�R>�m@��(;�d�PC��a�Z�i���@���YZA�w���H޹2��<x|���\�2�-�׶XU�]p}	Q��)ZԺ�:h/�(�Yb�r�(�w:�u��,z�ߎ��gG��v�e!�P��g����\���@������P��y���d*|��_�E�1*cAv��^`��uXq�L��2OĪ��R�t��6sK�1���x%�	��9A|�SB�^8�� �����9o��U���ʀA��o�[�w��+�v��	d$^�h!�d�x�.�2h��6ù������4��ipț��{vԶN��X.���r��m��h�H2���'\��x\�mfyߩƙ�����M���פ_*���R���?�Y�T�BlBmh!(��	+?/e�ǩ\G���6&ڏ���'G!�|E�b���X0�G�����\��s��s47Q�*!�;�לR��a�t+=S5��L��{mc��l![�����YA�*���
��.��u���Q��VH�V."O�OΌ�A@��䘩���6�-�t{���p���P��1��~%b^�r�W�ì�����xζ,VO7)-0;��دn�By<��|`eP�LG�9*������C}usE��j�5���X+*2�P>~Ɣ~=~�o[�w�����f�>��#EZ��+d�m��'�Lg_�bX��Z��4@&�
Χ�]�;�Ͷ��a:(��/�@IR�Y*��J�I��a�1�����5U�>���<eB�P�*�۞S��2�
O��vfӺ��Ԙ)��'�4�\TG�$S=4�c�i�\�d�f�l���!?SR�#��<Qo�ܚT�\X?u���Z!	=�o6SI�0\?��޲b������S� ��;]^e�SŻ����}6i[���ȵt�j��x%	�r%�$|e,��XRz ��j���T�%��ܬA0��EO�����M΃�k��x�1��(���M�ȥ�z���%��N�6�]w�V�z׸fs	^ �u;���a J\�g���pG�i/�<u���F��B�7dC�� ��;Ѝ?�N�7��;�곓bҕ;^h�QWIy��(�Z���q��e�\U!�=:Ⱥ��%�Q�Ӯm���=����R�6uuZ�� ���P�R,'�����~��u#�:��Q}ឤ�P����Ժh����p�x��v�3,���*K��̼�w��p��H��@;���ܠ��g��&E�@����$�`B ����V��>@9G��ߝ�	����J�P�NE�׋(��_�:���뺠�����aḳbH�-	�'vu^�S��,O6�[�� �m�+�Q`�r'A��������CAk/+?N�zI��Z���!z��� �&�Ք��Vcq�-m9}��V(
c��\W�Ո0�������*(6+�>�A�5�E�
��_�EH�l��.�HT��Q�y�]��'��QՎ#|�Y�.j���y�}�>Z�B>� W&|E5�m�}��i��t��dr�{�{�2 ��l��N7���ѾY"5w���b��7y�o5��C��E$gG,D-m=?����K���|���k�W��gg2m<3�y�C�&w�;��'���kM\��s9�D(�9)�u2����X�{���̍SA%/�x҅!�a�t�X<F���e[R> 2}�W�f�x[�@���"��U����s#U�����+� �G#�J�
2�r0�f���tW���#&ǘ�J�|�y��]��#��~�R?�PȮ@���?iP:�6 �w�9�C�V�ߨ��-�.�+��5�x_�<�[��4*��;Zt:a��-G�Iփk�DͿ�=;�a��V%XT_�k2�5�鄆����Au��N�7޵qѵ�? 	Q�H���.e���P��Ax��cGA[���*MT�6=g�RDd %�9��w�4ܪ�I�����{7';�|P� 7��*�m��@��c����4H�2s�_�ʆn�ځY���H��Ѧ��0��^��9e[���2m��Lȝ�o:�D$8�F�'~\TVԠ}N����"��J��L�Mu���y����a��K��$�[60�8q7�sGY�G����K�޴�s,	�<��d��0?�)ZW��H�(�Cu_ٲ�c���eb��Ҫ�E�� h���X�֩��TZf]���(���џ+	2I�L�'�{�.�-���g�2���W�p�t٭�3�2�_�XUP��\�0��U�'I���^{����V<�أ!U8�'J�=����ha�Oz��_Z0���k�B�B�S�9A>�p4�������S�48��FL�.� �ԍV��X���" �k#M�~]�=/I���}��#S@��8�_u��FRi��J�#Ra�`�\?@$�;�ᰭ�_^�ԸC�͟�((2���2c��)�M �||��]hl���Rh{VHP^����x�u��#�]�p�i��-UG|���x2�QM�r�0��.��vc��?�u��MB�)<� /�OI�`��NW@A⒍239���3�Oԕ�4~����%�.�9��,�4��A�`����/l:Q� nc��/���?�D�|�ë	ۚ)aK*�H&��B'x$�6ր���f����X��O��i���{�P��f3h؂�%�G&��i`)�y���V����e
����'��@�񮌳7�d*�9�AFć7l ������L��ad�Xp��{�εS�&jZ��Y���X��?0YFx(Ef��-V�%�n\��M�ZVnrc�\|��C03���P�`j�u
�xzϯ$��ʍTҥ"q�x�Y�����c���������(
�K�F�������v�;ϸ>r��8�� �ID2�@�	���������7*͹D B>���)ͼ
F|��#�P^"c/;,���B�a�Y]	±Rfz��e/xmtwK��4�٩Fk{����ǧ�{�IU�>�;�d\��h���#A;�W$��4&�NB��)�M�X����=a�T��&'�Nc	H��ϵ�r�������J���g���|b�!�>U~
�T䆰W��[@�c��w�E:�@�Pj!Xp-�,#\�4&ﻣ��D	�ӪH��m�(Il���2�PD�V|�1=n���7x/����Lz��G����}��s��#��t�Lf̧gx���)�aCqZE���d�n�I/޲_F�%"3w���Sc����f#x`'�(�*s���J��jψĒJ��&,�Hh�f��5�DS�^�c����s 7�l��ր��blo���oP|_�xq���:N����dG� �LU�a���ރ2$�m��Mi�+{�'��b�hecA1c��n϶�'�pwy�{1.U1T��A����]-����A�ȋVnYV�(
B����-�&�ڌ}3�� ��+ex�o��Op�-��\F���u�ow�{�+-GM�2��+��$9S�� �/��@\ϿGըFN�t�BLh.�EP�Ute�2��P�6B-�~��i�ރ�s�̥q��o�NR���C�����}�
�x&^:����j�@�PPq�ô�j#��+H��vzp�8>\���Su�jg���p?9��x���H|0�G.��f�}�3K�B�F`>,��Z\ڦ�P���Bf��2�}� �zӖE��3aF�-*[��5ِ�X�� w�8�ǁI�f�S��(]�n}����(�)�-�v��|������ЏϷf��;]��#R>��Ȇ�ی��o�����S� ��]u<#����}8�˛�	b���xΎ"���1���7n�ŷ3~ț�mR�<��a�]p*�kv\�<$�+��2���v��(sb`�R:��;_���#��N�j�a�� bg�Gԇ .���e`�B�����g����M�T:��Xxo��̽��E�@�yYGɣs���FeV����V�I�A��f(b�Y>�#�`�)8��;�Io`�1ݢ��@7�$0ۈ���lS��e�ⵣ4���N5�!~)d<J@�s�	�
�K@��Zi�q�J�AnYLv	�P�]:�t?#�^�6��#�ܰ�m�W�jk�n�,թ꠿��������.�ʸ���7,k�
�����7�ټ x� �˔T 8��w�k)r��:] Z��6i j\�2��ت��C띢��Q��Z�sSk��̘d��GOXx[f���(��{���i~f�9*υK��T�yC�ڇ)�`ՑPݑ�9H�\��ᘯfN�,j����� �����,�ě��WfՃA*l}�ԑ[4�E��v!{:�B誧�������;�M)���B�P�PQJ��3��c�3� ��oV!=��7w��Xb��2���4����&�I�;�������sE�3���"i#	�vYS���i������Nz��<m���GąӔjU��uh{�gx{��D�fU��\ ��/��c`�k��dA���-��K��L�'��E.�F����Q�~���D����/Ɍ12�#��Ejyk5Ect�Q���Ĩ��rP?�c�O�kjϭlc�J�u;�F_���t�'�s}^�X���I({9�ѩv);��Y��m����r:I�f���DYk�Oom!a�j���J��Z\%��]v{� �j�b� R�o�-�R��i.ť��~�tDNf�~�\��A�r���J:���m����*�3��|��e���:g)PtYqjm�"����}�ΨH��\�Ѡ�H�@��e��v�t�N<qh�Bѣ{�N� 
�B��zד�p�A� �)��`
�:
��⒬��E�"	xz��ʸ����w��(�ޖ�7H�(�	�Z<c���U��(��\_������׾�W��C"�A%����&͵v&��5���Q/� �/�֚�QH6źp�h����/1a���P���R�@j���)��;�b���{���MI��&�5�C|��i�Y� �	�'wK�4��lq=���;��aJ��/�F���;!*z��E1SHR�_/z����hP%T�
�?�>Nc�& _�Le�k쟭Pϙ���d7s���X��wz1�������E������u�!��M�2-E](�-c|<\��病w(�z�"��)m1Jf,#��'�T[���9x�
S��DU���9�&7�9]S(�X��H+H��� ����Վ9�}���Ϻ�OՏ��E��*-�Ʀ!;��	!D�Qb"R=Qr��j���}��XL��u0�d�!�d���)bL�<Կ^��~o꒠�J�Q��]V���1���M5a;�F�P�>�19n�{'C�ѻ�n��B�X��L��;8�H<��A�{S��cm�:E&a����[�������N�&�h[J��d�D����V�^jۭ�o�Y�x��k _W��ޠ�� FF-���8��̎D^;p� ��e�j�N��K �b�#��^��e��-9�k���:�jH����
�8�513�ԫ�"3��N;�NnP)�^ɑ�������-Q�z�"�3h���My����03��%;��N;?����|+3,����ܰt|X6c���ň�P�)�%j��eUKQD���GW,��o_�$,��L�=����+�La�d����6 �|xc�i�G#�Fw.됖�M���g\A�T�{C��K�zp����T���b�FmD)T>��BoU3�@v�������0C#怟�9p�W�rK-��(ME�9����	X�"���A��E!�H9R,3�i+Jk��K�;��
���W��`$V-�O��6˵�0ͳoR{H�C�S�N��n%U7p�����2��x�)P��-�E������P>&�@��}��������8��nו���Tf��EU��{�:�W �/X�(��g2'�?�5p�b��_���G�
������ xY]U���_J��k��BHH�o���2���-�Z���t-v�C�5�[��h�qi��L�&<�P/#%2To���	�W�᧶2�.O��ވ�FS�2�Ͷ*��&�X���zd�ఔ
��݋6���LM�У�B.�?M�b&J�p=8ٌ� �'H�������{Y�cDՖ*di��6�X��"�Pـ��Ou�٘��
.�m'�Xo�z !N%���%۸�\����|O��B}�0�Y�5�/c�Z`��0=�-��ئ�-H�w��r�/+Uƞ���Ř<C��J8�8��
�5�ʩ� 㡩���9����;�B���#F]e��q���
�f�X��_���,��Nձ[�(���ZC+�1�ˉٻC���\��|���H�����R�ÐO����rz�,�n
-��e#LWK��ӊ�dc2O�ɔ��?0"4��u2X.QY<Rp߸�����-8#~o[t��q��B�=A`��H<.���G�}xZ,tՕ����Ǎ�������4t�0}X�E�3���.�Lu�2A�w$��0�<�T��'&N?�k>�p��S !�n�]�=�!�������AHm�H�~���9�vHE�KT�ly�m��"��B[N�]*�:��i�Ic���9��,�JU���>�\�3Q��V6j�9��x5J��;�S��&�F٫�Z�G��Z.����>Ca��w��
:�]d�S@������q�Cԣ�����V�#Z���o��=�"#�c�X�='�*R+!5��堨!�����h&&Ѵ��譻W֣j��Md-��!A�n� Ps�L��/�"RW������;�]U���<����\�"쁨xD
w6&��,1����l�$q�m��:FQ7_{Gt��SQ�цh��.�0d��1�m|�^�?	�v����8�-!�P���[�����蚫x>"�R��I?�"D������L��;9 �q�MZ��������7�F��Z���o�u��7������r�x�0�2���b`���߈����1 W���u�6��)�������w	y�tZp��Em]���o��:�}+n����Fq>��3���mG@��x�ޥt=m?�2Sk<%�oRl�Z�;��+��o��F�ڵ��r6���o��ܗK/#�sэ5����^�⭂'%V,�xJ�A���g�}�ъ�q�Y�P�m�����u�o�P��
�k�9�(�f���x&0�C@~��`	:�L�J�z
%��c\��e]����c��%��^<'(�^��h���0�k�e=�O:+��$��"ÅA���v^�,ȫݮ�N6�v��Э�/i�B~��C��B�h�ŀD����P�e���?U-�?��͢�X�ɜ ��&��N��`qk"$*ȕ���N��5�%���z��^�F�魊:���IW_]�Ί��mEFO�9�K�N�9�����-���C!�� ����_p���!{��QTi�jA-qM�Y���Q����Br��C��$�	q"����-�;
���"��Aw��L8$�r�nt+mW>ڜz{F9և*�[�)�j�i�����y'c(%5��qÆ��H\>���׎��u wF���d>��]���z�#�
���5=9������?�d:B��a�;���h�hd�vd��b9J��<�0G�t%x;fH�T�u����6k=e��yZ"�z�"E�ϑ�O��C�/Գ�C`��f��|���^�=�@O�^ {�'wi},є��[�b����e0�y���� K���_�V���"oS�/G����s�	�;3���#��͟���=n��*1����|���0�4 y$/�o<�D僺2�Զ�B�]]lO�J Ԑ�RJ>>3���3�?b�F��'�-�I�	�'�u�8 `��MA[������|h�^o[N�9�_�;���$�`.0��S�%��w#�l+E�F�?鼑�q&d���A2-S�R�ݔ��3T������MZ�$����z�5�I�S[i3C�4�a�7A��=Pɐ�,s���=���s_$��!��at��$������&�74�҂hh�⊏���R�C�:����I�w���	s��xNN�����T?�i�	Xd����EȄ�� ��?��٭�����t�1���H8Y8e\&f�}qA/9�o��?��aͫB�Hq(�1��`p�	�jX3w�zq_6=���}�EᕁE=^�t���E���PD�>7�JY��({*p�sd�ˇO���1|\����"�I�?C�f�ܙ��T�����G=���2��<ITz��D�lv�ⵂ��)�	��f<�� ����8�����/�=��ڒp;�Kw�������"�4�Q���m�"9�T�@MT�M�U��:��",�4T�o#>�t��N��w���V&���κ��O1\S(Ȋ)lǈ ��{>�WC�|���1�<�ԃ% ����i  ��M9�"]����o��ɳ�ol0�b:c���]� l!��l"R��� m]�	 ���"�^���+޳X�����h�s������`r��V��Ő<�GH�5�]R>��b����<e�n*B]G��.�BOD�z�L�*��&[[���+T2��y��}�8n'��6���ۓ��*���s���w8���{VL����+yu2�oǐ(�{\;Qs��$6���L�_l��ُՃ��m1����K�1ۀ9N3�aisӬ�M���ݑ��ϼOܐ>�eK곉�		�Մ�^7yk0��]k��97d̅��[�ݷ��ʐ�Z~\��>0�hL�ؾ�܎ў�"�����8i�?7
W�|��f{gv��y"���@Ҝ�Et�!�� �j�ҫM?��O\t�!k�f��Ӥ�I߭�A퐈������y9����´��yXJr R�&�:����i����&���V�*����-����uH�o�*�ew�s�h�[�Ж4T8�\s)���g�z������t��`�B��}.�d1�q��H��u�xGK��)b-��)����ᙽ~BV��/loWT���F��Fp��G��SD��܍���R��
U[E�a����3�v'��׶���w���]g�� \��К	���4�Xҍ�94��MmHݾ^�3�/.��D�{�IVq�xz��h�,�6٬-r�ؘf�m}�Q��J�� �vv�r6.��I$�x�����B�J�D��-��	z�f��C�v��2�NN��Y����Ș�ڕF�����!}?u�#3+!�
K4n]��Ӗ_�F����u����Ͼ��3�3K�����-Bb�����z3��K�-O̘SE&F�̌����Ѵ������_S9c������;�I �<�T���$g��\��8���J���g�����-[?���@�c��Y	ؤ)W������Ƭ���	.���ޭ�"yT�v���Ad(P]�v2����!!o�q��[���-����T�k��"�_�3�yg���2V��8m�fw���f�Z��<N/MS���V�d�*����^n����F�JJ����7�ZP'����{��͡L�	!i����-�6���F^(��glǺg$Xllf�_ψ�k��D}Ny�$d}�;T����e�mK�/c���ќ[|���+���Zc��mr>A����*1��0
��yY�w`�d$�2�"�L/@������`~���m��$����)�,DL �'�蟷&<�%R��5��X��^�Ծ{�X��0R:ye�P����QR�"�
�eIw��Dk
R���Q>�^�mbԲ p�p��+#�0��\q}�I�8�������}��'���ay�=^-A��4E�Q�C�V�~p�bCm_��svV�4�J�Y�l��S��xTo�m�l�����C�S���7 z���b��r+R8�>��C��l��󮣕�ϐ�d\t���\�ǒ��,/W�`/t��|������0�a8�C#k�HqЀ����\h�Vn��J�l_Y�̶l�iծ]�J=��l�����h���n���_���N�	Q_gųZ������*p!�r��X��T�����r�ø�,~��*��bV-[�� �uZ��@$��w h�G�`��!���hr%��s(֑Vh�z9ыN�N�s�c�}�MZ�	�ы���0��ud��8R��9`� ��_HU����̜�c�$�p�H1�f�/��qjJ_���
v�
"��]^
��kP�\Ϛ����]H���n<������r��DK����\'��RрI�^X�\��T��O�޷��t��Z�;��;���+j��(����$�0��A@��=��)J&OI]u7,��xv�Vɜ9[׎qj4�C��S�%<&Sɰa�;��i.e�.l�#<>�]������;�V�0�[",��+�0�;�8�,5�.P�-�)ji���XȺ/�2�̿�k�f�|s>C�[��Ra�:t^���,�ں!�+��k�SG�5����C�1�"�� Ƃ�#�H?�>�B-����N����F�	^��uZ,�C�R!�S��ɤ�*>�|�Ĩ��Sg�b3c�#W�h�Ƥ�c$���6f^�Z�Z�E�ݽh��/�ʠ�]���?1O��f��]�q�*�A5K�W�$���B��Xg�x�����N��!�<G�*�ZxWk�?��JC�>�d����y�����O�I�vD>L��.����]��:�1����%ft��|���Y8�''�a�0f��F��.iic�ʀ�XzOyMM�{�҉�Ԯv���r�vx&���|d;���
enZ��)�`v�����j�d+�zaujgY�<�b�h�4��!�#��[��y�ޕ!,&+PI�u��y��p��o��X�=\���g7����o�׬��V��C��m��ʧt)N��m��|R^wL�P��>u����l��aAΠ���ͣ���3��;bϿ
>�~۳��Ġ���������9���<�A^�U�/0��7��W�^�	C�Zu�S�(���r
ӾA��d�١�g|��RZ��j�Kk�����)���ZDR�@��+ˀ�K<�-����o٧�6���q��7�26W�c�ٌQԤc���I�һ 
�l_���fW`O��^/,a�i��bH�in�<��a0� �����V�ʀ��,��0u��W܁ʼS/n������.��#-�� hy*]��̀�O�u�Iv,;�4B��5�0�k�q0ū���^�� �ɠc�Cl(P�J"*�t��ߞ��*�Ց��|��(u���6�l����dj���)sWC���7�)yC��x2��F�G�%g�4�����
���0���q2�6�c�I�)9�4�tq���g�Dw����bY|&:+b�͍�l�e��GA�#���Y�� �qC��X�����=x2��Ō��