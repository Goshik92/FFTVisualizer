��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�`��ihۨw�R	���K\�P���x2�����G�s������?_���M!Nɗ�K<�&�P�B�S��\/�u�D(��r��V���]l�g
{���ӭJ5�S��(��n��W���Щ�;
q��+�6Ұ���1��nʺa��y��R�#ys]�.8D�F�~���=nX"����_�Q�˦^�K�	w���(��͸ ������)���\�7M���7Tk��m�o��~GF ������hmbW\���afN�tZ����KLy�N��/��a !�KƛQ9g�h��s�Q_����G�93KۓF���z�V��r+���?��Ivśx�ПMS?�� �ri^��_�Dh�)WZ��lf�Ks#w��ڻ�86��^W���j:�ɖ�'�6?s��?҈�l&�/�ȵ'}2)ᢇ��dK�q��3��gcBB%-���d%"E%La�Q�>�RT-֭��9C����00�p�#���۪W�:h`�j�l�K6�1aZ&���+3MY��(���\�朚�ϏV�c=N�u�袅Wy�.U���#�Qd���y��S�$1�&�j�YF���CW{Yr�S�'@s]��s�1�H��p5l�2����4����/'f�8x�b�I�c_bغ�I�����Ȑ��wr0ʡ>�W�r��i��nڥ��Kv��Κ�MК0������*��{J���4W��Vӛ~�^�z/D4�i�&���Bpww�6!U�P{�zA������c��L,⯙-2���k��r����t�^?P�;�_�l�[�U�[Y�7��A(W�AX`���2��S�bXٳ���br����VO5B���黟�n�2m�/Fu�c]���^�s�r�v0Fт��־tz1a���~��Y8�7�7E`R*�L�9:F%��
t]��H¶׾a��_�2��Tn�k��BŷF�������ou�^a�9��.@L"A���P0�uk�����&*=T�/@ѪTC�p�7�q����ӹ�̋�(Xm�#m	e	�z!�o+P��/�=$C� >���y�)����瓎 �ⱂ���S��b��x�0�[�y�-޸e �Ҷ	/jT��<Mǧh�T#!���ě� �� nr�1�!��C���_�>(W%q�K�����%+��x�0���_P,�p�,/qw*(%�	����w��8u�⫳\�i2u>��5zx��߶�� ��G���<���nQ�=I��%���D2UYݓ��D���a%!�2�;�x]����$u2271�$S�H\Bvcr���3<Ւb%.�ì��!�T,o�+�O83�M5,��qC�>�wA��=[��DF�_�������>Wc5�f���9E�2�#F����D��g��#������v�7���d�^���ߪs���\6EcN:�`������ǟ�= %��Xרn��e���p�W,ܤNf1ޓ�hM��k�x�j����o�Eb�-���Y��#NViE���0?=6(P89�u���LZg�zTL������2���`&b��!'�!Y�ƽ���ͭ���������c��#re|> 6#D���p!&) DoC/Bw�����F��"ݛ�2'�u��4�R�<��,2�� I}���1���np�\����9��6�io���S
������<��A��<����Z��z��AE<l���0�[�
x�����7��v�z~��oio7����)W|T�l��$>XNu��u�d�����)��������rJ^܋�BK]�{�`'.^
zM-C��cޕ�(q���_K}
$�w}�΅�0n�Sg-��>��;��NY� ��o�>�-m�(¡DF�'&�����QNL'��in���BH�[
��!%�'}~�]�^��$n��ٖ�����X e����9]>t���p�X˸�N81 $[C_<�,�<�f��gf�>�q>ة���K^�=XB��eQ<\I�+�Qn�+��vP���������z��I7T�Bb>h) >��Q1�\y<��vq-a��+ d��_8d�o!���R^�����8���w��6��&SC#�O]@9L���RTܽ�������V�����
��8�'��3>p��o��R_������7t^�y6:At���322ʷ��n����h���f~P����y5����E������:�"rn�(r�����_S�,�.DY�Ƹz�O�P�?y``�8�]_���"��Ef̓gO�(��C�̷�@�r,�*�t���`�1�I�O�l���H���Ǉ�W8e]��aT��b����K�C��\5��ևsgf�Z[ڇ����%q�P����;�M�~�{�D z!��݊�$������N6N|���B���&nM}�,�R��`Rv��ދ�\���ޜN:`�l�����hmZ���iA��2������}c_fL����m��m�\��R�$ 	|�O�8d�L�����7LvW,W�����w�����IvjS�HE:��~���lYO�v���T�`�Vh����p�J8E��
t���
v���:Y�J}N� ��z=*�u��Q�~/-F��t�t>�'�i��⼯c�j���]jv�=�]U�#z
�޼|�Um`}�?�ʩ�2P|��M�RS[|�� �� �Um&���6�ym5��
!3��c���0'B�Z�ߦ3��9��U�&A�D���bw�M�5G���@&L�}�Ƹ	�|ue�l4pg�W�$L�Ů<7ش�h�!̻{�@�a�8���QY�I�VÕ�C�[Ū@O��q�LTp�@8^�0�>ª�H�t���)�j`x�ɬ�ЛQ{t��'@=u�7���%@�mf޲5��6�`H�`M�9Et#�y�tT�D7.�_2eS�V΢��P���1e�'̘8��z!�:��mjs�(�B�(���G���^��(�$�����i:�`[���hF���(:P*�o�t��\����[�s���^X���U��L���>����di=�y�o�Y1c����1��������>��x2�'�N��k+�>����'��q���w��w�$Ȭ�y���FME�=R����������u��|LN�s^���}�����a�`G�>m�<�Y�i�v^b�v2��U�Aϑ7b��cG�r�����S��p���P]�:��RL��ؘ�׹n��￵�!���-W�?3����$1��&:�P3>J�@�m�m�1Pn�ĝ�_�fis ���*�z��Z�<��c}��we0qC�s��l�j[�ǯ�]�A��u���C��)�?�7�~�KD�&�7���K���~AѸi��K(q+��9	�Ƶ�a �n���D�.ނ��U:��-r:`�����Ç;���*����5}il/��F₍l�E��PE�}�P���w9�Ϥ���x��n���A��Y�Z�%��ɀ6�תg�~�a�3���jQ!9��Io;�rZ�����.%s� he*�\�]��Jb<��w��AdS��(y�Q�Q��Gլ� m��ͥ�╜�O-�Vc�j�U�
��Z�_H�/x��lY�KMG���~C��j���s?�¾��H���� Ic�:���6�~_PϷ�	�D�yg�C$�'��#��ۋ;�q'�ԃk�q�vo�Kny��Ŧ�ڽzP��U�:C�_�V���X#�<�*`{>�2�E�<=!�g狜 6�(��&WC3�ag�(���r_�,�\Yw?%�TRȊRB�����c�Q5 �-^��TK�/�8�,/�g��~�>���-ħ�;��JA�.�K^�XM7��17rĤ�No��z�}�pƤ\ �U�1�:�	dP���$uT��qt�cY)yנ@a�4����DM�H�,��,��~����x@�s3��/S��O�8�R��>̨Bá�	?O�Q"��q �
�Iڭ07:�۴����J��
��f�Z��8d0ՎR�P @�Q����?�s\�3K;Y2��"P@Pڒ�%ǉv�Kۨj]),�DMsWI˱�D��ŉ	Ir������1�\������a�Ɉ.��҉NdNs���"Kle�^�Ob��I��!�q���Y���!�z>U7mz`�C�gâ>B��ǃ����V|��*�7��8V�Y33�N����^ӑ�1�7��`�����0>��Z�%��aE�j�F�P���ܼP��p^�Ǖ�a������s�N����@������)���~�zP����v�]�U���Y�|�1�'3�q��/��Xeh���b�o9ה�{E/�V�t���0�x��r��,����h��p�a�j����569����(K_���͗E}%�X�<(�\����C�A� ֝,W��̊�Ws\ �Z�4�+�I��E� ���p�;�Z�a�u�b�D	��Fd��}`=ٽ���6����_�g���^Ū�m��2R�v�����>��|�T�Ծ��q�RQʼ?\W��Us�z�r!`�u����}�$��N4���՞��Cȏ��3"��sC<���B���������M��ZvhS-�!�PZ���Q�(�*6�)�F����e26�S[_��ꪤ {W��!���/��\
wvdE�YL��ѿ�O=`mȓ;����+�Þj.v�3���^G��t�� ��~��f���+G)f���C`<PH I�I%��~R�}���BTJ�`đN�&�v�,��:->7�����k�}�n�W�u��1��M-ӵ!-2�E�;��nC%ie� ,1�2��&��`ھF�Z�w ��+'�e4~\rn��BK�Z:��Q �-ki�b\�2+<8	3�k7̞���h��%� n��������%��&�~Af���T&��H�S`�Bb?~�K
�߱<'Z�̛n!�O@��
~�ެ��#���ԓv}�������#��:���&���Tt�K11��i��	�%�����B��m����bLپ+i�݄d���6���d -��d�y]k�>7�.����p�5�2��ν�Z�ͅ�W$ާ�!-e٘�"`z?��a���_}�.�F�(Q7�'��[n��p�L���3S��a%�9���4�P>��̵L
�鼃�ǘ�/���������zI�� ����
����́���6��7|&������2t:���,��E=�u?��I���b!Xc'�y63���2
��~���G-{�[�>�e�(➴By7�� a��7>���[d�g2z)�'[����Z�Q��8F��MsD����WZH���]�Ezo�����+��3.��x��a�݆�4�y~(?0�@��s�?N{��]3g|��v�~���u)�N郍�����o�Cj`o
��YV_ʵ�|��Pr��8|2�{'�ۘ�C��f2����Z3�Oe�*�Z`KR^K%��Qc��p�1��a���/ɪ\H���#�4z�(�s��Q�h�	�z�w�}=��G-O����_f��L#��n�i�^r����;�ź1w��-:�ѶӕFP�84 �j� -��]��v�el��n<�i_�����/��[p� Hcg������s�+�+rqjZ=�-��y�2�ۦ�����^�Dp���Gh e]5������fI\�Ō�����ۡc��ۈ��~w�И(r\��<tCh:<��⛲>}����&���+Ǽ�K��"�,��`��m[�8k��u��=	�(�4M�7ǋ ��rl�hI�"��O����"qfO���X�;�&��}��n�ݯ�s���KU�Ax/O�����J���E���/s�k��т&�)��>ҧ�
��w�u�dK�)|���a�D�fs{~�f�������jE�����0<'I�nQ|�v<�%��$�EX������q�fC��~�H1qGg)��]1����n�t����ᶲ-�q�$z(��
e�U��>7������3��}��1�a��!�Ȍ���@ ;�lv�"�`��)?Q�`~�6��a4�r��	�f�ـ����Å�ĮwG����X�R�,/�>U߶�e�0�5n�vpO�Y=��,�.c`e��$L9�2}#��'�}y}��3�j��`8|oW����JZ&]�����80[8l�N�������rq�m��U��VN?����-.����= �⣑��J��7<�E����#���z����2.�K8�'
*(&��TyU�?v���n�Z(��/����5��+�(/�6��Ȟ�7^U��hT�1(�{���$Zx���3%
w6$6B12��5�<Mm�0��������&V������E�X}��B<L[�����~��<�_AZ�B���'�U���Up�o�5�%��o��{t�\��h�E�[��:�Ǡ �������^7�����H�(L�"H��,� �e:�,`y�u�� c��]T�B]a����֘5�Ǉ�ϩZ�߯��15��ҏ-<Gnt��~��I�xM#�;?���h���P�8�Xݕ��;�T�Ơ��Ja�J�V�l���6�Y±�TyϽ6�PHY_<H�)U(��;��h�r�b��r9��.�u5%�㘣N4{rP_WkIF��y��N�|��� .�7�,h	2dS��)��#����w^
��؁J_H	��N=��L�d����72�R�V�%�ׂ�d �Q�+]⺺Ծ(s����A���-�؟s�o:&���Yt��S��b�)o��@���M�d�QuSS���꾧�r�X�o�j$/7��v�tJ�8�x�H�X1�E@s~f؆�R�C7�0^��O�8�LQg�6T�d��&���&�i������U�Ki�m	X*�	���l��E��(�J)x`��<�q7M7;}/��^{�J��l���.�TޥB�^�q���v��Tf聛oT�on{�	x����>�}^|��f�1����d1�6~����;�����<��;��(�zh�|�����j��ٔ���Q�qa��$+QϞ���t�d�,�t����+��(�:�UR�1 ٕ�K��=Cj���	;m�FA�[��~F�|�9�c\�ףaUܼ�"s�-�D�M�O��?_��G�$���J=�u$���p�Bf%<n�~������H�����]-s��h�N�-����E��rB�RV�R|��~Ȳ0�Z[��pZ������	����n�6�G�7�E�H�F����Kg��vl�r�3��{CK�$d���z"�sD��kD��9ѣ���b��t~����Bahƥ�����|fG��&�?�����Sn�)�l	$�"t++�?�%,�Ƨ���ޓ��TN ���e�̍�&���럭��?��S���u�>�l/�hR!�g�#c	�=��"}[2���Z�6HM��(:������ED��5�,X�bRoer�1>3�X�B/��P@���6���ñ�m��h~�F����/����'/���"!����� �N��}<BR��4&�2?�K-�)Tr0t�w�ʰo��L��%[�M�I���S6�̖v5ka>E$�Y@D ��?���;�b6��d�) �vɌ��:���ogT� ��Uעz:��Bco��U�#W����NS��b=���D�����6 X-Wg:!�q��?MQV��Tԗ�1�!d�ʏ�����R�O&������`�T�C�p���1����!�Cb@�W��Ux�O�VQ�*id�#`���oY;ܓ�訛���s��p���3sHy�{t[o���)U0�yRǏG�E����H��sBED
iԽ1� �I�?5���l�Ә����Ep�_�P��_޴{�D��}ɀ�˺s��5�Hd��U������
z4 ]���8*���L��tj�����!��e?,S�l�Z1I�q��!W ^"��U_�JL&GK֥��sA�����	�;*�eo=�$�;��¡���JO�-��"�rN��#�x2��-}g�/G�0���u�Ab��{mε~��;k����	C?w� ��/��ۏ�F*G�J����as����'¸�>�E4��@ZY����"�:/�)�P󲈷�����@��4��a�����;�ȑ4�"��Ì��]�В���#8���oF�:�-.E@��0$��8���f2r�j�z�ڍo�N����>��S�qG�q�������,'����[^���;������h��"����]��m-Ō�kE�Vn��Qo:�x��%Ҍޟ@�,�	' ����!!jҡ]�g��-ɑ�{�4�+����b���b$�k�\Q��.���:��l�(��{ZM��&m�bHY3'_�g�}����p��ǖF4���7��%s|��a�N�ȷt�X[*�Y	�,���,Đ�oxF����֖8;db���[\K
��$�|bQ׎��=E���:�"����% <W-����l�0�s�/���t?cd'������O��D:w-�lO�A�M.G-�9L���3dd��=ǉ��$�~�~�
�i���[��%�v��Y�R�Z� ͊p/ w�yi�`[jU��X��:D'��;�'3������_p�����?�]͟^�ʛ��ɻ1b���F�N��<�<��y�|ّ��<�tT;JerV������v������B�άC�=J��Af�j ��Q��r�j𒚲@��������D.Xk�OVDc���P]������?�$�Ֆg���T�C;�$#`b��P��ӹ�<���W�!t��o��Το��Q�G���%�3����P�3��]pQt���	Y�$��UUsJ*��."����d�8�w$.@��	д�	�M����Zu��*ٸ��RY%ϫ��,H�yG��h[_2l�$x�6JyN-��5� U������މ|o}�{Ѿ�{uk�"��@���qm�׿�omǪ��-(�ϫ�F�^����Ҿk�J�c���η��	�������X��
i��<G��8e��U�����׬`�?'���&�/
��52X:�Wrq����Z��e?�����D!�gޚ@�"G�In@yv+q Y��$?U����#AfJS(UH�ϥ��k$)��M�G&V�xY��2�aM �T�ێAJ����2y��l�:`0^�����������^Ҙ7���0(���?[ MrB-數����=	�|�$JRP��$t/+e�&����:y&X�ۮ^�nM�@����?g���ϷᲒ�Z���� �M��
	P8\� �"�Q%~<�ﱌ%���w�QӏOQَ�hǶ+b�}_`P���4�?nP1?�'�RL�6�@wR���:8��9ω�|�ct}��w^
���OX��m�:��$pP���{��j�� f޸R���9c'�p}��4O���������!mS��eR�yB�m�_I� <)M$�����Ɇ�������f6��"�(�/8�[y���w��JUG���+j���.X�]���W��O!TD�{.�&yF*ڱ�I�l�C޽W�h�����fBj:p�Siƞ�f��ڇ|�#�}%�P�2n&���P��<��O:rn�a?�7���lBO,�������X�2g��5�x}�C0a�{[��Ʀ�)��#y���k�uL����>�|�����T��)�S�qlI�8��Vr�\�Rwx���Mb[�*Cd;��q����r9�*��>6�Kؘo�wͯS�񊡔 ��u!�S�ޛ2+x\�R�K3E�#���aL��O�P�I�[���M`~:�}�r��ȿ�S1�G(����7��s����ҳ_� ���nRÍ���'�D�y�}`� (��	�Ka�
����d����J��U*)��\r��f�d�<��-�\5NPw ��Y9[����#�8�����(�#���-�Y�g�.�\\��pT���ƶy)Q�~�VqDg|����qL{q��"��UP�`l���	9�0���^���O�`B+�v�c��k�Q�:N5�Q,��nd�wT]���ý�C��T�it2���5I#	g��]�(Q�ULN��Ը���.4V��"
�_Մ�_sU�B�P2>���\���[����I�ٵnW��+,���["v��C�v�T�
�X#r�+��ȉ�/;_'3M8������v��$�-D�����A��B��W���K�\���v9�V$����}���CG���]��6ܼJ�1��M_���y�%��D[�K M�ۡjS�]��e�}7\��� �m�k
"@d���]Q��:̍;#�UOE]kgZb��?�:$� I#��S�v�=�3�d�/��A�G">�  �v� �8��q�#���n��җ��_|�	� �v::_��*��	p�����G�&���yꪨt��nt��ݐ�
�ܟt�}�+Y�q�d8�".�ax8�6�螄�ă���&�� ��5j����09�1L,xD�C%f��"<>��0欧�NOGs�Zp�qSS�d%��)E����M�z"%PNh�x�c�ǃ_>��M��r?�����Aw��pnW0��%7�x�7��	��6�|��U|+#v|����Z�<d����=y*:�� ����i�Q�<��~�i���3�̾�P�x5�\M�FAOXr=S�[orYg��ynlQ⮼\r�����q��'hR������UO��0J(�mX�ν�G�lk����&�q�h>�!-9<F��m���O5�U��]&��ł�d,j�P�>~�Zd�&e�� ��'��g:㱄���j�>{�=K��ŖT7���&�#����Ɗ��i,V�^�Ҝ��>&�	K���J��%��@��&^��q�u�&R�������tٮʅ	θ�T�t�7���qX�B�\2��P*Q�/v�L�M���8[�����	v���b��,|uHu6���۔�&j�d�7��èZW�����|�6��5Ƶ�4���TI�����;#o��F-�H�)�2�rp����$����Q [Io�5����C����Z�@fzd�~��g_�� �7?��T�!6z�(n���D�*��$�p���
�`�L��SGW����܀@&�c�Y@q"���^��I��\�T�/�a5���&B�+,R8��d��_��u��F�(�D��M%��/TW2ي.����(��/%;�ێ�:y4[
~���o�1��j�0���͡�����;�Y>?C��(��ߖ6���PP�֦ܽj��xn�F�hY�]�xn�l3����fR9��)Dg녾U0O�E�Z6�k���I�Ԅ{�9̴cJ���?,D��������/�5=t�
�n����t1l����ˉg(�I�ч��e�*>����X����CI�2@�.�27��6n�G�_��L��s$֭	b��"�`6mc(��8��%Px�CM��_���J�>	�$
(��Y�
n��������!�	Qk{E��06wDj^5�	�E����;j�������6U��S����0\�_���l�Ď����Ur>���n@�˺��u�3{$�����4k :>�0�Č?�&WO4(Y�Ϳ= �PЌ#"��0)������B����,H:��*��Ȓ�����G��zi��`۲ѽ�w'���b[d��V�t`��"}����2���]3Q�"��7|����?��0:�tQ2��u���cү��|9G�S��s�0ւ
��^��e�?8���yC����.u?���G�ṹ�p󁲿I+r#f���D����cAC���M�
��8��]��A	qB2��>U��dY��"+k�]�2ƭU:�4���=W�D���g>�q�#�\��5��v����� 7fX�L�?�ps���W�V�������"b��%����A���s�ӳM�]l�.��şj�s`��uQ�ټ�Ϋ�X���8L$�ْҢ[n�����*���WֹÚ.衏^Òs�ȵ�o�)�6�x��y��=���n�<�B�} ,���C\����SG�}5�Zc�(`O��������??��4���D�V+�[x���D4īG�6�����G���)s'^o.Z1<'��7���m��PVR��\�ay�ͼ���%���&]0��GK��:@l��@>:�?\(Bf�)��,S�"^�L���A�dKb=;��J!��԰��A��r�|����|h@O#��A�?��䢄�)q��b�o�/�PjU��T,@�\�F����g��}��Y��N�j݊�_���0{/=q�%ՐB�L�	�x�x���χ�9J�(`��`��Q�e� �~�Z��v����a���
3t����vd��}�E�t��`Z���1�Qd�:|��3eE�����7+�|`�  ;��7���C��-��\
�
j}�gу��XFa���:A��AUSr�*��$O:��|�N< ˌ|�[�u/q����;��l�]�o>��T����;(A^X�D�S�b��;����RwOMH��'��ظl_ѕ�^�ډ��p\�HR��e���ST��
#M�n����sG�
x�'S��\�������(hB��#��c��ʒ�Z��~�P��Q��ʂ�w�O3wq�adԵ��o���L�ǋ����7'Gʿ��ߨ���{Sj�h)�$���1���0����3���߭���hT]L�=7e���[ ǆ~��?����E����?\AX�Wu;I_;�M���|$֚d����1�U�8��߆��ۢ�O^x�OP��*�K�K�!� �4|��{�k�1��Н[<�S�K>��Y�}~
�r�sB��KƚZ��Jw}����$��xC"�>�t��e�U��_�H��4.�, ��~�\o���[��[ә�$�ĜBr�ܼY�Z&�&e9[��xr6B���A#��øL,�j�'�k���=3�JWh:�S�-O|-r]�_+�: s͚��&�4\J�7}����(���M`W�3��Mp����5����tYW_�:�v�>)o؆-�Qh���_bR�F�q�;���J�xM��]�g;�	l�xV�"���(�cv)9�;^AJ�>=��Y����4͒=�=g�_���O��J�X� 	ߝ��Տ��k�s�Gjf7D`5ܧ�i��{�R�쌛�!9�b��߽[lҫ�D=9�"M�ξB��;M�R���r6t&\�N��K����j�}q��$���s���ʂ T6� [%��I�̛�����~m�>��7Ԕ���Lڊ�6>�$�lvWǚ'�i�5��m����B���d?�KR�C�#Q�:�&��ې]�]�s�[���^$�>���	a�c�G@a���_�e��,n��@?�a|yH�
�
�
��2��O3 ��K��8%�_��]����ګ*�Y;D\��V �{��TBӷ�Ϣ*[ 橪���db��p�7��h��̖��k�ܼ��zai�N���#7.�*��)�h��̰?Dg��w���`dy�������T�4�R��xI��(@��>X��H%��s��qFd0$�e/�ŝB_1����yp8�&�[�p���}�w����A��������SזQ&�Xq^�[�A�k��gr�P�߸~
����ٴ�;�U��b���7��+{C�7әȡ�}9����r�չ����(��~L��M���T�8P.Q�aS��j�ii�vVx�P���)��ʡ�4�;E,K�(�
.q��֚r�f��Kw�",��O��!b}|�!��B���*ܙ��_` d�KOȔ�q'n:�����t^�o;+���.�9�&Qd�o2ۜ��,hiษ3M^�2z�5�̀_�������l�*�=(^-asݟ�#�\
�f|	���:>[����p��<)�{1�[����i�>�*�>���O����
X�]�qZ�K֖����<n?�+�X6�{�bH�y�$�ڙ�����m�p��u�ُ񱡕�i�1:h���- E4-�k4t��ΰm�H�~�?����R��&4[���iJ�H�Z�.\��Go�le�	�����Rm���
�Ȯf^��ނ@~!#(���ɮ:nl�i7X�hfd�)�
l��C���z����#[�!E��q�b'7��m�A�a^�Tt��i�'l8�>^@�a3���[�L��U��Q��i��wʫLw ��fѐ�Wl�Yٹ��^�T��ie�t��d���q�/qCs�2vv~��2�
:𓊃�#�����'m}���5V&ب5���9�k�J�|�+���3��MT��)�I�R%U�MN�R�c�Yt��[^�3ޡ]�O˶�֔�WD>s���� �]?sآ�� ���9C}�~�C^�ҀS�����)0��p2�k-߾Қ&Ёh���-Da;J���A��4��у5�%�"�yu��9�皍@m������v�D^ѩb��j��'Z��O�VV���+�$hvr�����ǈ�,+�
�����͑�uÜ��"���s��B��T�K�N���uEt�槞�� (������I�����(���f�����Ib�h�:����PAX(C�;'�͹����E���oן(A��cXr ���ß�-F��o_�o�[��%U1�G�Pו�����C�~g����#I���Y�@��h��NS/�"����Oe�-��L��	���>�h�/����p�%]�j~�n�{m��yK���D���9� #|����͗�4+$nbȬuA�����\)rޫ���Q�m��\V��&��l���9*�����_p����f���Qi}�p��]��!䝨���
���v�������N��_C��n�V��"㹘�^!姸�kq{�m��w��$/��0��6��=N��_��;�?@�mP�S�d��y8��俅H�Q�ܫ�Y��\�՜�� �ґQ9�>��vG�t��` �u�SR��Gz$1���Zz��7� )��վ�����^�ڼ/m�g�����d�fK���=�}A�ܳc{3�-J�����F�DSp+J����՞�����
d���\i�6�^��/U�4M����_!��6H<f��%�~�џ`�4��~l=d�Y��aũ��4������F��Qͽ�ap��Z��'���Ŀ-�O�}�Y�*P���6"�3G����z8��2+�{w�3�؎���zG�S���|M��$W㩤�=�O^>B!�S�o�j��A!
�Z:Y�2�9��~���1���C�:���j���yr��6���Yo~́7�	������k���6abU�k��ʀp��1q��q�q$�tR�g�*�{�N�^A�]���!�J_�;M������ybu�X�mD����	�u��=CKтY��C��ɗ�@6c#��Ebn��?���_�ưu�b�"�7z�!̭k���v͎��y9l���=ƚ{�3�����L�2���p���Z��R�����Q���7�b	>Beǳ%>�7d*4v�#��<��G)2+I�J���a�L���!�F�G$�4tb����/uED�������c]�Ut���Q���M�����.�T����i�[/Z�F�TIpn�U��
WlUyƊ���N�b��&2�X���Ϧ�W��9S���NGs�Td�1��![�+'�vɦ�B��MWt�m�x��{��cB>�٨�X��x>��%8=������g90?Y�����^-"�\���tW�`��ܣ��� $~�,-���M_����OA?�Ӟ�+q��əTٙ�C\G6hb�o�Vj �ML�H�N�`�h�Ou�r��?����L�__��pt���o/� r��j���~"W�?C'v���K�#Ww��㍡���9�^Ҏ6�D�
�e>��	~��IZϮZ�F�c�{4�4�AMx'�-�G,c#�\s+eV��1�����g��!>��ِ�P��a�bV�&�*��Y�(����bY�$@+�8�Y{�+����%,NZ{%Ծ���E:��#�D۪9¬I])�mM���XoD��A�0���R�xgK��s�"�.M߰6���r'��=��loA���OH��W��|��x��������lr�́�5�YZ
S{����O_�;�zH��Fw?W�X��m���{@��!��@CU�	˚�����!{�l�]=�����5���^`I_�� ��9�.\�Ӷ���S	]����*�\�O�R4�7CtRQ�!�Yp���S�^�PL5��*1	�LNh�45��)�V�_�G��mQ���p%"i	=e��A� wN,%ڸ�-A��(�.A�Ϭ��6�I&I=ǐFr�r=��12�>jWt�==����}��;^^���̦Cő}i�(-�s��'S��[�ηHp��"#A��N�:�Nh���B�\�œ�����r���2���R`4� �$�Â���e��?2"kA'毰BD�^ղ�����:�B=�����:��Ц;i����@<�Eo��͒�Q�3/���1�Q-d�6ӖA%5x��?!��S�����O�L���ѩ��irx�z���~-Hf��JƙA�ɤ�q�q��|2qMlxj��Ɗ�����r�syOc�3�5zRj�@m�Z�4Y���#$P8��8ڿ�h���h�˘f�����dK��>l��%�&A+q�8`�寢�g�vW��V���Α���?��?�3�Ǩ�A����=?��7����0�3��_g�?F��d�ș��%8����_��-�����t�7�L}p>tF�fc�s���O0r+M������U��.���$+O���׻�s@�@�T�F�eS�'@�j7��p^��<~�����t5~u�їm��� A����g��U=�<�m���r��1ad�
%gc�:��;�B%��c$��Ib��\��\�O��b���Lr�4��Q@��>�9��/2�i��x�dD��tÜ��>�/[$Vb>�����P��T{��O��O��L��E�d��A����(�Eg�?4��ʨ�:	g�(<�*h�q�����HI=N���[�3A� �3�>#�O�3�� J���,��mϻך^a���y�"lښ�c���I���~�p�J F�����u@!+ʢ
dh��W=�n�^�K���k(����ip��یlN�ȩ�].x�G���p�bZ�('�.�x��f(���"�6P��|#uZ�aW��)(9*�O�C�U����X�&z���.�� ,O�]�g��aEP���?ĮAL�Ca>���ܻY1�W��*Ż7O�՘/�2�G@Ԯ���xv� an���m�z��f�����ݪ�żc���Y���}��-�d03g���:����%,�wx���N� yo��4�Ĉ�mY���s����"��l@�����'�ZMA	dUM�����V�g��7�=9T'��~'�dNŜQ ���{��2�R���:�k{q�P|Rk��6ͪ-�{����4ܵ�k�2[1���1@v�a!���w_ c/�6���-���8�L���'͢M=i�������)��Ai>����P?�y߃P����<w���c�Kr6���Z���=C�"���Uķyg��-��K9��� K�峹B�N!m�G��<!���Jm�w�����j��r(�5�UR�fv�_��3�&����
�6U4��3
����#*ͧ�yǁ"�8!��`'���u�:ƏC>4��ݻl�;��S�[�С���
0M��P\GK��KMs�=�a��uL�Pm�"T+��ծ�R�J��@�A�����vs�\�g�9B6S�AG'҂��V)�n��$�Ԫ|ie2R0�hV�u�G�M��o�y��~=������U�i�i��s�BT�~����ʒfŞ�<�_����� �C�J���dQ(�S��͍[�`�0�+g��*~8��"o��[�-50�"4G�Y���+W�Z��Y�jk1h�iR�d0�ێQASh1x��
#K ���{��=�U|(���c^����.��W��/w�%�-�*o .�<w�'�,��ѻgd��XA䡢��''v -�eX�+$���rp,�5ᥴq� G�eA]E�/��D'�)��nY ��ʶ����	ɵ��A2��6%�7��c�� ⾫�#[/���rMk?�+H�ŵG�N3�;�/F��:R	frX���n��
�������{�W��t(M�鹀�.r1�O�����R�"@�	��y�EE�/�)�mGQ�!��j�Kj�a�#�97��LE"@q���#�7[fi���ǅ�(�|8`���R��x��C�� }��O��t�d��o�O��x����ftp�m~�~%8Sa���:b����ӱ�bfg=,~q�gh��D�Fr�_��� C����s��T��g�)�q\����:F�+�AB^O8� �0�c��h�5�R�R���5w�ι(@����1![:��w��{-J���d����z��c_�F;�����垒Es���g���_1}��pΗð�S�3�	@�����*�����l65�u�*�}�2B��U9���={o�<�?��&7�,c���8�Ka�s�p���'!��r0B����(r��\ʰ�!~/n��C�:?s���rk+�A���S�i���쁹��C�WGt��Ç[[XŅm̙�R(봘K�ȔY��p�&NV�ۥ�++ǅ�̻���퇷ȣ�q������ Ì�rX�=rT�a{��W2,P�숂(^M-��c�s�fFD{Z�h���	�Y�V~�{��}��� i��1� �����ͭ��N��:�)�dg�ֺ:��9(��'K'�4h�-�ޱ�w�5�s�"��c�H����U����N��B@p�YMW qC�&:�Uف
�bJ+-��.T�i�J�E'6��e�����d�kmVO�tW�-Ӄ{f����I�v�a##&�iJ�.��O�JA�kA��*s�zM@����	/I��^O���\�k�}�%��cZ�>%����G���k3;H�>6�#0"��*�� �)�P���䆭tG��^����A���k��m�tĹ��{���k�Y2��ۤ+�5��d��B�KɾƔ[��+�꿟�~����ߨ�>��cŞ ��D�v���P����4E_��x��+��V��z���v�*�v�/���J���m	���<j�����b@��J�3;��Q�c[ƃ�i�9�9m;��:|�>�\��x��&#=�k�&�����6��LL���T��ddX��ڂ ��.�7�m�"�;-x?�.Dt�l���J�<ڴt�G�$���0A0Β�F�͛P[]����EA�*h�3�k��gל�rs�;gO@���oEE�ىt�������aO��swpt����y&��탍tk�sG��JL�#�*�&���g����KOS���5����|�ׂҌ�RR�L�+;�R\<�^C��j���U��6g�����3����[Y��\�ͷ���T$}��3 ���)���N(k���u)�|��������L 7R����#�I��[�D�¹f�g:���m)7�!MCw�ߔ^�_���Q?jRTǟ��VU��΢"�e(�,c^��֡gy��,©9~�[V�pܕ��k�|	��Z�xhX9�����B��B�Fl_���;�sw���	a���sx�v��1�BI+�kb�����KR{��_u�I�J �&�_ڸ��%�B�u)mD9bZE��4�|/�IV>��Jx��/�sr���da���}s�/���E�Q{w��?uܳɎ8�;� [Ai6RG�:�Vv�?e�������Z� 岎�Ӊ������.bKx�~i|(�5��.�>+2���_f� &��KH)�@ę��cE����:��o�c�[h+{�0�,���@���0X��b0���C�r��}};m\e�V!�V)J�'�u�p�0�vzPcC#B���Y��I��Ĩ���D�%:	E^a!wX�n�6����-uE?�лQ^ѭG_��&_;%��=5g7��}v��ɧ�:S֗�������4�
{��32k��u���l����ߵA��6�Y�җ��:��6=�����0c5(���B
�iEO���QW�s��( ~����Vj@f.E0���9�ݧP]�� 'ĥ��:�ؐ�;���}�N�,RclҦ�van��Y>W��f�����Wh,��J���7�@��YX�1uJ����|A?1T�a���B]g�+o���$L	�2�L�z^��/�.�\t���n0W�V��MNQ�+dz���fW�e��K�Sa!�HG[%,"���:ER�L��[h�r��~��ذ������e��GRc�çB�C�(��}H��HfxF��oi�=��L�A2JXK��
��,���)/�D�g06f�]�=�����xh�d'����n6��-�� t��S¦�Pq�#�����Q2}�����-dF��0�`����Ӳ}���{��B}G�� Gkv���|�����dhD���n��"[<��9�����*{����}[�����
3��ǖ
-��"L�v�I�5;�'�\*�.�%/�����d��ZɾR%P9%3��?F2"�����M��?&�8ش�����W}���RѩU�<�f��S!�Y������h����t¬�����9���]�h|7�����T�Q܌�
&��k]����)�'M�m6[x���A<߅�3����m� �PD���lh�E�B��י��f+�%�On��0ZZ��ZP��/�֞әA�SRvB��|
�B:jNJ���-�=�霐��t�~@�@�A��N��o�(#^�XaM�;�BW��/.z�N��F­H��q���#}���,���g��IR�_������^,�f�����⫄u�cYv�K�X��@U�8��𺯀�k׬oY"r&}�i��lг�6�`�*�D��i��e&�����4�����P��O�r1h�:���u�Ϝ 	�1&�@�����0��C��2F�B|~�Ro��1�lK�A�:�p[&�ڔqL'-0p̖EF�Kl`��v���z�;�!O�����E+�Q�W"I`�p��Ba�A�4wy����6�n�m�ă���_�	��q�@��| ���@޻�EG]��jIՉѪr������ҕ-����؇Q{���q�B���r%d�@�o	��H��.���S����&ȹ��PED��))�r�h�ͳ�K,h����w��D�7`(a��wETw����W#86�4�G�Ғs﷜��������7����x;�)�F�\�:6��;k��D�ugh�� ������C�����╞dO.R�y��*]
�I��%+�Z?Q�x� /�ǵ�7/�3�ֈL�xA����L�E�.,��z�����r��BY�DD�E�$�P�K�f��	J\��y=[�E�����E�mҽ��7���������Q���J^�+�8B�n1HUX����6�9��93	����yHy�o� ����h�z����4 *��\SA�zB���@�F��{k�38nL�;:������5�����[~�v����%�֥�TD��$�ҤQW_\��Q<!�rǳ%�}�
��`��9�g�k�z�}֩]Q66m
���$Ay��wwW�ή,Lz&ź��n��R����,���}���`q��G&�64K+���i��C��a�ثDW�G�M^�0s���D�W0�t���9�r�sOq�tz��"Z�b��{?�ѭ^$��������Q���e<N���������j;������i6�q�.D?.R���e5�W����#`�?�gl��dv��#�
I_�f%c\}�T�9�]�(���8���/~���Qj�,	���g{9�a� �Nxk��+.��9ڧ���B��P{����]�'d�3�;�/�� hT��Z�|/]K��i�^�b�y��Kꧾ�Ȝ����X�\��������`��;�QE���E�s���/,�ރ��<�,9��3�����4��{��Z��89#z� � ���h����J���~�b~C���R��*��5�9E��V;��DpQ���.u�r��U�_��8W3,Ƈ�����+>��!�W�ɸ�Y	�XB���{+���͏,:��S�E��FyU9��w����<>~��Ԃ�ˋ���-ݭΚ'7�lJ�|��>����X8���X�dr�5u�;�䘓0p�ƥ_wk�Ёg�'��{j�Jc�mէ�,�XaO�\��mן�(�q�{ڕz�45�z|xf5t�8@+,�B.f
dYb��iy��F	��������c��e�p��������N��*i�� &�s��O�<����"5����eOՌ_��E�`q0��o����C| �!�9�v�G�e�{���E�f/u߳I_��x*�/����m�✛��}�P����C�������lM���XFrv�1��^H�kU���RJ�5z��GК�����^��L�2(H��X
I"�0�)>T��i58�O�2��HPO�(�~�v�/ӿ���?��I��jN6R˩0�7̉lg�I�R��8�|]瓿_���b��<-$q+�rf>����N�0�#'j�3%��L�{�:�`��[�&��nt����~p�t<8�FN�uu����V��<k�zj���n �P??TT�pU� ����o��´H����:���.O~�=A�y9^��5��;�K�i2k�: j�F2��*Z1�=��˔+�l���1��*��O�1�{�<q�N~��1^���AKL1�R����nA���S���*_͔V+����5����|!�Ġ%��]�AF~��K�b��dR/��eTn��!z��Z�|7 ��GT䶻��&��.��]�Ǘ}ے$a�o�/e�`Q^����)vJ]o��?2��!W���
���m
}O�v>,��9x��O4�ο����Y��aʧ<�C\�i�q��=���B�UJ�d�L�HT�O��%��[�� ��I*�������#��2�$?I���gr��K'��i� �.c���OD���Y��`9����|󅻝�̅Y�>�< $ΚYB�iACe>��_�:]�n6�J����1���%7rxcB�����]S���t��%Ͽ��X����-;���:c�/�CK5o����#<�x3��9ߎ�a��y&Q8 <�vA���I]�7�VZ���̕�K�����Ӓ��_I -q��\�5�}s��R�2��g|0���?6@m2;����������Lk^ ��!�"�k2:��:ܠ��� #i��s�l�-e0�a&壬�hS�s����:�E<��k���q�ˬ�K5w���z�*8�l�"�mL��j�-�q���bv��$zoc�Dܘ_WR�G��X�� ��� �s�"<|)����� �8�Wu��\�^�j\��n�����6�*I����B�q� ײX3�"j�=��g��BB��z�_}r^�T,���L�k��j����M��WG�;Ys�|A��!��+�N�P�����v�����U�Y���#�J`���D6Z�w_�A�H�)x+��z{��|p5(�N�xvZ|nw���9A(U}E�����0ȩ�U�٢����Ț��.��S�UC4 L�D�53M�����7����B�T�W�5��d��C%qP�dh�rc1�9�@�?W��Xy*Rߕ|V��wEy�M�Q�v�  �m�P83���D�H42�?�F�Z�� �+�'^��xfiL��'t��^KON,��Xh��p=%o5�y�2$Y��U�D�?rr�i�s��k���do4s&1��%��@��KW���R�S6b��b,���W�$��B�&J���{�������t�K ���iWQ $��D�+����2j)�����p!�2H���_%�剦ht�i�ZYQ<�HatK\�Yr��_�2�ĕ�õ�L䑏OԘ�*�[��)�3�8�
e2�_���F�<������~>�;+~��[�+�/��mpf\~.�L�5On� 8A7t�
�ߔSuƍ�;ѳaϊz?�܉)ӓ6�Y~Oj�y��u�F������MЎQ�mTz����OU5q٭��c�FU�G�-2�K�?&��]#�ʧ/���=�QN^��h��3^���\�V�Ε6 ���N��C���sV�}�B'��ڻ�A%m�V�$y�EY�2����ҝ��u��#�z�^�¤I���d���U*����I2mP7m�觪��VrA����ٶE�[�$�bQ��^�px��.K�w�T���|���N��*2�P�d}ܑY��hR�O�p�=�����
�#&���1W�x?d	��%�ƈ4�l� ���~I؎;j�v{�vU%��U�n�u���hE|G�aZq��K��b5JN������p���ڠo8�k��աc�'��D��r��pYt?A<�����!�^�ՙ�dJgK/��sG��\K�o:\k'8��me�~�������s��������eU��kŎ�<��6���}G
�R�% ��a�c��`/�y^�\!�@����Y0
Q�T	�Bf(h���ьZ7ݎ�;3I��������3�D�mȵ+O��G����ѝ6��j̹�i@}C?�$�F����k��(�VDgaa��q�(�;Uj��#ڠ4v�,MKht�^~����#{�80(�lV��Y��q��Ү����i�$G�i���9>Cr��?VY�@�3��{���4���u���8>��m|\y���'��tli�?e��ͼ�/��6����f��B�1
��H�V|s�wA��F>!���,G��Z��e?@r�DQ8���"a�f����h�͊]�p[�eVW�hSv��5��h�w�d\��ӱ�S�@���g�0��5����Rq���#�c�,�w��j���\��)�5�h]1��OB���U�4�	Ō���+}OTdB��J(T�a>���H�(�}"���I3B���O���M��L���ޖFr���.N�C��[w(Y�t�!S8�D8i�_��;X0�<��4]kf5`*��2:s6A'���X��y�)�L=�U���`�5��;�Ŭ��Z�6Y}� �(���<p/P`��
͜�anG�y2վҏ��~.hʧ`�N��A9�{PSݰ�2!]ls5�����膷�@1>Ռ�I���w��'Jx�
�m$�yhQr�}mL�]B��~�^���2O�㸓x_μ�\,*�j��Rk��zh6_�ǹ~N]����/�?%b7�'���2�}�TQ�<h"�{V�V��Ϊ�'F[����ϼֽ2��m'8b�Mf�(IϋP��c�b�UjI����EyQ`����ee=�"}cW�0?�([���v�#Bp�!����Y�x`FX�ш7qjhdF_K�L݅��A�PE�C��@"��8���X�z�R�^�4�E0������ɛ�3\i;�1�3���(��x�G'W v\��?���c�J���S��W��J�&�!�g\Yh?h��A�>�S����/UD�� R	��.'��"���*���8���gf�0�K�l�~�mg�6���m��ެ�.G�|�rA%BU�����x6רE������-f�	k�����K����<�HY}2�d�Mӷ���RN������k���JC'e�S�J� Ы�Юӥ��2y�6��2�',��r���-�ܦs=�`������¾�l��BW�5�΋p��=
ж�J����~U���������oC����݆4k0\sh <�\%\>�������%�%��L]���F�3O�H�%v1j�dM�=%��S~
��K��8mR7��q	g�.�ܒ�<{\u�C�j$����Y����0.!BgQ0ˑ��g&��Y�ͨ����g?��H�h�Y�b�/�\Ʌڏ9��X�D?q+C��'h���}Q/p\�]?�*�)ȸ�w������x���qU͜�(�t�ij oX/���C�]�"��_�?4ӃHJޒ/��s�����s�@�\����0aR�9��zx�����x������m�͉���`�ʗ�;hZ�?%���$-|z�F�)�{~�@Ӆ�����g�S_h��0�l�C��: �̸�e�N�J(��l�IZ��`#�� �̂�������Z{v��o�_����zʏ�f�I�5AL�N`�սcNo�C]���ϯ���<H|e�"���W[Bj!S5l���� Ys!�DFc�������a�mڧ��B�@ ԍ)�܁I��iaȘ6K����|�/F�S5��>��o�^�I��W����|��r�4j*
<����wU`��Q�C�qWܳ���#�p�Ǿ}�=�.�Xqc 4ݒ�f5��&\ӵ$Y��!�'a�)ח���=����l-h�*�^��F�������ϡam�DIWn<"ػ�U�,���B$� UVD��1��}ޣW-߱�i�#�ٟݖ�O.�T���wʭ�Q�ta�b�����Ky����HUuT����Sc�y�� ��,.���p�����R���h�Uw+�q�X�?�?@��6��%�"�'r���eO��g��Sl"�ޛ$0�R�2$G1X�I�{��4��W��O��iʱ�Ɂ#r��c���d.)q����� cv�iI,Vŭ�����4�io����\ӌp�}�hgOt=[S��w}z:@���~��Ƣ�ڟ����p�������T�̴��)��{�¨@DQ��(\iBIt7v;+���I�ݽN+����d��������Of}Ξܼ��%L!���Ě<}vq���-X� @�S��,�Uk�i�I��l�Y�^H�G�W�q|�<����z9c.�'������ۭ�pQ�7Uo�O<��{���>����i�%Dx��p�%�)X6���ÕrR�[XB�_�-h��*g\���S\���ʔծs�0Դ&��;�M���J�p[�.Ă�ϳ�*>[h4�"��P��v�ԏ	T�A���T���w92��4�>)��/���&�J��� ���a4��y���p-�-�I����~���&� F�|\1B����#����m��h.����V�=,'����!��e�HO��/�#D����	!�P!q��7�P2�tt�k)s��B�~�e�\��4j�wUE+^�>ؚ{�+#�5ع ��]�/1�uA�H��E���<ŧ�#��%�"|���n�m��#�K�x8���Lܟ��#`U�ۡ%��O{^k��L?��&h��NE��s3�u���SR:��p��0+��4 �!9���\�k�퍼���h�0������;D��x��ׂ��c?��TLFl�*91��i[k���*EƜ.6� �=ʝ�+"k�����O�ZaT.�)��0�C���G��'ء#8��D�'�g0Ce���Ь�<����Ж�S����x}tB�ڌ�@@���Z>F��F�� � �oGW�X��_e���tE�ΣP��
�#a���5:m.Kt�\1�q1,�]�q��-w�w�[�$�cn�̵����K	_�jWY��ƨ���ҿ���P+i_a���|�-F#�e �Lv�S�͸F}HH�L�rO3�1- FCVǼxD��� Rw93�&Y��:<BFBxM-��t��6�mߟy������Q�F[!�$rϡ
�n��I>Z3ƺ�-���>�Y������9 �t�˷�jSnT�@fϪ�OQ�Je=u�[k��=�%���������_��/0��]�XMi�B�_e�C{�~�li���uG��d)�:���Sp��=te���͆�n��Im�`~@�ɏ�QD�/=��P����̹��:�ѵ�?~���'�-������w�e}����êj�l�����Y�����:�y>x�Prջ6C�]�`����)z�/Ҫ
k�O�����I�+!+Q	V<c�R�o�i��8��t��Z	���?h�I�шOJ
"��~�GJ��s83��6�x=���/޾p඲i;j$�/Ⱦ�n�
���E�[K`vn�a��{��rc/�ݤ�z�	�$��b���?}�r��ŧnΖ��>1W^\NE�:/}��Wc�w"J`����t�ʼIi0yHA97x�6!R
���C�*�?�����5�'��X_���T^�e5"��h�i�$"C��!�7ɧ��?��'�
�����C(C���2낭4]j��8;��9{�pfݜlaC�L<J8
�;�Z�G�k]�$]H�%Á-{E�/ gW�gx����!^�NDo�l����T���7c�2v�_P����m�]��`0�D�}��i��Z]��C���A2��l�+4Hs�O��S����	:�F!�Ӊm��_��,8��fM�3*��U�W��7��d��.�HYl��q��������J�����u��X�Gl�z��Mx��-�p�6��:�f+��j� gZ�&���`�} �"Hǌ��K��:�i��e�B04�H����PL�Q<x�1�9Q>/���Z���;s	a�+�\G�ȼ����П
z��e}�Ԋ��|s����rҍ�-T"!
īI1�l�j�d�L�����әt�hI�����P�	<����v/�^��B�|����D�<H��ev�m	���0L��n)'g����Z�˭���M�h�֕�"zQ9/c4��m� e3��W:yq�wc�2���X���I�SA�B3���Jv#d�o�~�1�V�Ö��'+x`�]E�`z��N�

�1O�+�"��5o��Anӹ`�x�f�J�8=XR�yN�a[Q`ʕT�S���3[�t*�'����JZ�N�D�L��Q�<O9�1!AM&F#�����"�GTI�j.9�[b���iZ/aN�+�rb"�mi����A�s��7ކ��n����ʫ6�C�&n���d����E�����eO�s}�@ȶS]���C� i)(�1���".�6��0�mdqe,m�����'Ӱ|e>���A�[L���o<h��d~�k/SVF@�?�	��C��h"\�
�*�Ȟ�K�Ƭ���NN��Q����9ʯ�Mq��Zj�dS�L�T�uOk�\�MQ�:BT�%9TX��eS��Z�q��	��u)q�Jq,�\;��^K�*���y���¾�],�� 6�`��0F����	�
~v�:�i�G΀� ���|H�/IYR��J<���~8|ۍ��<�	8��{��Z`��ͪ�`��==����Ҁ���p� ��Ȍj��O.�9����H[!���1�Ě{�zʧ��S%�g���I2��e�F���8��B��M�~d�{[��+�=G
W�����=ap�n��<'1CE�v2M�\IZ�D����9�
��g��ŵ�ohF�4�c��(J|���K�i�$as�F?���W86{�G���82�+!�M�펝������
��'�j.��̽jd�P��O�� &�����,���� n�K�	د�{4TU�3�5�8z���I�S�O��}��]\��?��k"��y��!ɡt�k�}fa%Jk����̤P`o"����f��Q�Lee���|v�%�t��z��5f��d���v�mJ'xZ���ۑ�Z��5!59ʮk���-�S@�N6Պ����bĚR�%�-0�b�����=�G�ՠD��u* 7Aic0�~�!������n8�.���ƀ�˨Ƙ��Rg�h U޷Svs���q�6.*vʱ�g�=�������Ʊ��;�sxo�Ͻ�h�1��p2�9w��aS��D6tyEf�0��M�����v��^ӭ�l��\ڇ::(�³�C�F{j�#P [����X�,H��*6��v���/v�|���"���=R�̠5�Nw����A�y��Q�h��dm
����w��i?[�s�uư�ŕm��p҅�����IW�{jI���f�d�|G�i����$��H�Ae��<5&������r�*m������Z5D���ig�0<�P�]	l,��'e�ث
���6l���Jo�%�}�����xU��4��6��f~�oO�i)�Fm�����8�h|�ɠҝ����Y���)(0�Z"��@���,Ad����M^��e^����Q;L�$���&�F5���$�[�n�#������#^��nHǅ9�u�q������FrPx��۷H4����yTޖ5D;ǹ,'�6(TY�	tt�U�ޔ���6��ܲ�ʳ�h��2��^���H�t��EN�q��?�8r5����Z��>}�;q��͗���+3r��>�G�:N�� ����],(��s�nо�E�x ��v9]����;�.��A���"J��.ð���!;���� ��c8��%���-�=���߫�i�� �&rC`--��^�5����X�PI
���kWf(�Q8���HD���4�oо��96�X�H���~0Ph��R@S�}17LIHhF�n�"y��h�1kC޽.7���P�ZS5O�j��΍j
ʤ�M�%k�R�[X�[����֪�P{T-�TL�_4���y�Sƹ͙�!��i���x�U�w�_��VҠ�?�����ǭf�6��O+�.y,a}L��Dȼ��gD�)e횪��N���$����d��:���xE�=��9*�7f����HA=i�δ=rp��O��n�ٵd���\R��G���`T�C'�(��^�xH��@׏l�O!�j#�i�f.����	�/�嬳�@�m���}X&�U9Z)`�Z�5����X�Q�Hܻ��3���u�ͺ�%h�Uh<�^�z�,c��)!�U8r�bC�$��GH뚘h �����h<�S4Y��ï�NV2�u��|ٮ0�p9�c�aƖ����SOR0����~k=�}����=�;B�i��߃�iϔ���Q����1�q&@��8Z�qxE��bv�@�_�|���eH����b���4�NȎ�R�P!�q؍�󇘮d�zע�|��J��
�mn-����l��߁q�m�{����gC�y�폭J��G`h���y�!���8!��Ph,��q&��t_'/)6��l���w�����R�~0 �c\��S;}Yڒ�r�m�34�G鱵�H�
}�\2�54>�͛�3�F�ɵ*䙅����.i�F~�&>/j�䪌"�O+�� 3>!�;�x�ܞ����&\Wߗ��h��`M��9F�l�'Az���G����b��8@�k���C���+k.r�q���ɖ#?���X�fi�=g��VÖ!V?C���������Jo��Iw�B��n�P9���t���{�K�=)+�y<]���_�F�1�Eӛ�ѐ�Meʵ���x�w����p6pV�7&�r��(�U�YEd���m�� H���ɚCu8��X�C��Kw�I����}+�E�?�������˥.���uݫ��sn�!��a��\��9���>���*��1OHN�*�"��^��J�Ͳ������*�!]�yN4T�D�� !/�����[���#��VJ��p7�`����o��W������\?h��ӭ��uq�@�n�=�ܖ������ǹ��$*�5��Ȏ����d֨�L�g�|6�P�X̐X�X}��F���O��/5��~e/x)�M����r�]�B�C���H`�;�%Zj�c�7��=j�t%�vh����M���ݚ��{�y��I��+�Be�\5�j}�@��j�w�ҮT�cb�q<O:ល�E{�f|���1}��Yu��0pf��ݠ�פ,Qt���	I�*��҃lK���'�W=vO���`�9�}�ELH���_]q�٪�d�X�[h�����5j��R[� {Wݲ8�1�'h�S��V��a��݃b1��gߊ>j��*1�%L��Ȼ�iu�Y��d:���|t���vX��񗴽�pqY���I����Y�3U����Έ�(:Nl��O6X�;�݄Ӡl�[��%C���I��4 �0@^�֌��M��W��O����
��r�j�Bi�29ы�Q9)>9��	�Zp)�u��[���??�Kx�J�$�gBBC���W�N��tǸž��J9[[B�`۲~�����m��=���N,�_н�������"��8in+	�ie؛n��&U��;�@JnD��(����+Te8���-�{���x���I����V��!�f��]+lMr�T�����A�!YK꺂$�k$(��W�[xZ�2���j�tv��4ˑx�8��:��Y��jl����>�z�s����P��M���D�R�OP�A�Tt��mv��h#?*����j��Y_:�&�R�Ex�w��&��B�!<�u�YY�5�L�0�/�!��B�u�F�����Ú��M�]�����M���̄���x������0���˔XjZ1R���e�+��q�U5	l̄m1OŐ���FD��2��n��SN��$��Yj�j撕X�nhr˭4XBq�j���[7�ljH��� +��/��� S{�u���nV��B���z|�9��R_���s��ܫ��zz�\��Ηk�L�Z���[l ��5e����.�6�4Y.�G�2���i<��@h�2�Z/����= K��\j�"6��l�頱�ή�FH�F�N�ҙ-ҭ)w�,���R�+>o�-���e�Xk���]|��q1t���FH�T�;�f �ͥ�q�����]0X��/J�6��� r	�@��
�t\�|�y���3wa���ۭ���E�ݗBI�VὩ|���x���\cL`w�O��gx]5��\��%����.��.e��G�%�8�I
)}j�I�8lx�xF��� �rhm)�
|�/ϫ���X"�y������R�O�Z916�����S���+e�W$���mCR]Y[�j/]�Uy��+�&����M��V`i���(��n���Լ�����3Ң�.��(�\�u��N٧9<duۭ<�ېݡUD��)�ڡ�V�*��B².>iƙm�v��we��S�[��wCuL_ŏO�C�".�Ҵ!�%���\�T� ��"�ƧSz	�:��N2�wt���ne�e�6m�t70m}�o���0$�4��Sl��=�:��ʮFt�Ɉ7ل2��xqQ��)P������1��Æ�k�/T��h0���vP9,!)���w��2Ҷr%^����������'���F�q����y��X78�4=��ϖp���/�t�;^���4��bI$��آ�9!�<?T����w�%T�;7�,@�n�a��2]�z�}m:ؤ$m���!��Ǭm4�*���>�R��R�.�[��]��2a�A���gYc�e�PD}���N�^ o�\�<mX����w�{�;���� �����hڻ\�,�/���q�:
ȕAo<k6��b5c�\�J}���<���t'_�R�W�|��s,	�6���� ����������-!�I.Ex������\6[d�+o3�����	3Z�#?*��֬��m�X����27]��uV_�T���\��ڨ��8�$��}3xЌiV/>�?Ec��>!����'cP3���p�Y�.�('��p6+-�*��:��I�(���P�VX�g�]*���H���]؆ <��i�M���O<����R��6!���Ǽ����j\M����p	���@���^}�����]k0ZK$�[S�^�O�����1�,�2��{>���CO�a%�wI\&�����dY�2^�\�痛�7�Xe5,^{��ka�Q���=��_.������/��:���.1��Y�3����:ܖ��y�A*O-~��DC::�V�wh��5�öF�����N��%wi����	A��)yg��qJ�D�[ڴs^�(��NI^�� E$�X�w�4��QGP<1�H��Y��2��,�Ӌ2X� �F,tc���I&�I�3�c�~B�YC�#k�g�Ұ[d,�3�!���"��I�:�����P��D� ���Y��a*n�zѩb�@�A��&x�0� ��w$s���<O��>�wC��X�����Lyt.�1U�������!�NCoⶑ���I
��E��?s0ǱS�3���];'_H0����8�lr�����3{3I�]�Xǂ��s���L��ޟQv���VV�ya���y�A����4G�R���O��^�.�;��tة:����o?d���0��~��P��U�n�|�_Ժ���ʟ~4]�V�$���a]!4�d_^T��~x>]c6�'�VR���zjX�kN={�5�;�xW�@�a�
��z�4���)P�ĸ����z=c<j��Q)!����>Ԟ;���j�̋fƶjţã��_ ��O�7� �-��z��%0��/��b�722H歜�.șN	���J4/���H_U��?�KoU�	����Zq����.���W�8)�6���?��u��q�����^���?rRK'�˽���"ñCk
aL�s�\Hq�[���, �0��H�x�?��9����Z�*����Rs�i$}@�k,Rz�dgS2�d��C;��S�a3�*U��o�w/���^�l������@ب ���Y�6��*�ᦰ�"��"��w�)G����~2�2�����[O�k�+�)W<�O�΄�t>�|=�Xg:MgG��m.)*���6�W�/��[�E��� �#�.�s��~Ύg|��e�� �l���|��}\ �ओ�<p�17�_�$�8�O!����j$��ۇ<P^
f�%�W�5���T��N��b� Y�Bs�1U4K�m:K��b�9��%16ٮ��;�*��R4�Le�q�?�C];�9�lI^��pi}�2�Q�A�1�_X�/
�f$�Չ��.0�%����"W�v�!h)�j����JR]�re�j(���du8��M.�i�C�I��^ĜʤV_h�Z�Чdt�R:����%?����j�Y�} ��x�b��P+��i=�Ќt�i�셅�����Rl��{�1�,��<���[�*z���4E��i�v��t9.�
H�"�q
�5@z(�\�|�R�3%�sB�Wg��ï�n:�پL͸`����L8����n��OBn澤�AJJ�)�'M���Y+R*�,w.1b OH�w�	�8�e"��O�>=mp]�ɲpǕ��y�g3	iS��/��sF����H�P���k[)��o�
�a��%�6��~�cb-`�E�'��etݹ�����	��� M{F���.��2�v���"̙-r:'���'��9�L�༜3D��_������7���*%���i���@;��L��3�y�t��W�2�M�p[���-��V��~�<6��z��<�p���<��ϋ�s���'U�	�v�R�8@xj0b�)e��o�/�����D�A~�@��:!�˸�ņXz��2
��s����b�p��ERɱ���){��6-�Ɛ?*����'��1� t���=��������S�R�"ԥ+�&O	(�ͥ����p,)�<��}
_�-(���W�4�j.$���8�3��D7�(?���0s�zjE�G��2�,��B		lXhx%p�_�7���K�<���6�-�8�i�|�U�S��yk���t�dt{��׈�5#l��k�,JEݹa�yؤ �?t�ݸ�4]�`�Ն��3"W2
�Ä�6�L�fE+PI�T�Y���,�IƑP��h�W1�
���&��ċ���`��bw��A�b�C�y=u�=�\>Q�>���)
��[�k���&�cM��Be\�D��=�l��o�~z+�I)�X�oÕW��Ғ�Hr����х�18��p���{�N�{_�Zq�T��!qƠ���%�����2����/n�����ѧ��(��� ����xF��N��ZCy���b���s0�_�0�Lן������K� �d�՟`_����".��b2%�*�pW����fw�M�E��H��/xxK�'X�J����G%���NOV:g��WLPz��b����ү��'(e�*Uj�9ޜ]1�r���ޣ�#k��f���7eٶ�[h�bxx�#��ʑ��0���8ޤ嚿�eH�G� J���72�� �!ho�����dWXD'SD�g�w\�(c��2�(��E	o�2K�ʩ�����I����,R_q9I�^��R��\�/:�?��q�����b}�䅰lfS���dK	������r��(�ڥz�������p��`�n���W-L�Ò.F�������R� ��ki[M�8�ۆ/��ܙ��z��_���`��-�;0�*�/zPJ/�6��qt�Zڇ2L�V�]�+Hn�A�Nِ
���d:\ŗ�c��!ר���;��jZ�u�O6���c���5xq�*��7ʃ�T���'���a�dƴ�vD�$�����$��o��.-���y���q�u���ב��0�`�/�O�f��۬5.�1O���p�N�iY���v�C���o'KAI*h��߬��ujP~�c5t��>��V����]g�&,����x~O��^���j�W�'Kj����8e�Ӹ�ߊ�v7hS�r������V��9�o���ѸVW_�p�u�1fr� m�`���[�cWfbN-E��P�� �������3N)�-����o����c݀@�<��]�,�(�:߈�NM��־�@�s��@獨�Cb�y�����\@�~I����~T���W�Gy�e���PR&m�����j�r������J|�[n�u}�����F��T�
�"��Q��P3k��qEs�����u�=y�k�5��!gQ�ӵ�2��l ϶1��a�~�QԱ�b��'�s{x�ih+Xl#G��t�Z�2�ؤvRe��B09��]�Ȓ���3��<&��cf�Z��4��>2��{�&�!	�a�B:]	 �Z���KB�ƿl���^�����2�-2�aM?���mv����FDs�cg�wв�:���b�.A���/�(��u	)���e��ǧ�9gw��9|���&$L��DV�Q�v��'[�.m�#W~F�.�m����ít?���~ye�;1���1�]��urZ��k��%=�D3��C�@�wC+S��h[�A�� �Z�U�!nl��Zv+�@�s�-�]��Ѐ%�}��F(��.�,l>�0R��1#��B�Ȃ���<�'���<#S�j��l�if�	����۾+P��ѹ�NZ��+�2���M1�)���هC���J�6��.�-�q����� ���j������k��:���P��
��������n��I,��'����F�1��k���OD���TO�}P�!FynC��)���wKP��pA�b,fn_3��0�i�Oے&fb�h�PV:�ڡ<�5�$��\�&`�2��b �2��D�b'綬
T�������F�l;:��B-�5w�m�Bws���z�*o��z����p�.7�xs�d���m��6��.ݏ��P��'�A/���'�O֯��8�'I����;e��N<D
_�je���x)��oW��0�۩B�dHX6BJ|���%�/��B�`��'�n�_�v��>�E�^N�J!/ ���=�&�if�5Bj��͂P�i껈/eݳ<�ke��kW��������������x�����WN�W<���/�_���,�I�,�$���|Q�_