��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0]��?l
�4�!�ߦ����"�p8"	~��kB�J)��NbM�L��\jO��#y��r�3wA�y�}�S�{�����X�.m�lM(��R�g������B�*�NV�X-?����$��$�3�s�`;��y�@�u�ߗA�R�|�Ԝ�+�)]f��������҅i[^�"[��t��00��6�ĔR�*[�]�V�t���9�c%kz�Q��*N�| ea�z ��@������mU���h�$}���~�k��'C ��� Z���>J����ׯ,�'��3@akCc�U�U��?��a	6S��K󊀧uh���Z��&���9�+�)�b�В���ɀ�t�]z[��z�/`� !g�!*��P�����I�<V�� /o"�����@�g柅˳���.���5����9�i��)�!Ҏ���f8�vh�3�Z��ZC�:3Ϲ@�+��&�Ư���	��������Ϋ< �����"�����!b�'G����Z�!�R�l��Ã���3�����y���H�>����/{���?R%|��n6���gJ�2!b/ΧW�}�/FM��%����� ǜBk{�.�-�ّWz�*J`����'29�05�J�NYŪԚ��N�F2���������q��y�-Y�	����D�0���7��%��,�-.�O,P�y�w	�	�JT6'�Z�Ҟ���4��\��י����Ə��g��y��E��q�"�ӊ��N���H��`����=l�r�Ed�tP\��� �c�G�����/�('�'˷5����+��3]ʸ�:xõ|D,"���V�d�@��^Nm�D�dK�+l����E�ȟ��_��O�՟	����ȢM�6��������U�²��;偐&r�+����q���_j/�/3Ew�?'�Y���7ϓ,4���W�X�`]���eop�B����nIN�_K�����+�-�J��^��8��c�.)��+eR\_�-�/��?���}��@�|�VBp�zq�4���tsT������wPφ�(�,/��3�3~����]4�_x}����M��t,�Wv,�,�t����#���ιXz�^U��#|n���q��LlW�'_�@aQ�Ѽ��Սu�7�q��"�u$��NɌ'�Ϸ��z�q{$����o��9��*���t��T�=��|\�y��;��rMfV���_�fx5d��Dj�?	�V������ñ,�ʥ�Zy�rZ�W�l��3��b̉�8]k� ����L^��j��s�(6Ew�:)Ko� 2�\�|{��O&ɇ㏇=dr�7.�)�|��9�l�~
��*�
�a*�}�Ug��@����C��Ox��f�-h�H��G�wuV:lg���?��i�����k�DXܟ6*����jX�k�%F�+z���ù9(41-��*�Fd:ܚs�[.���J��":wԱ�ӷ��oQ^�@���,i��l���G����Q��"Sp�x�&r�.��J�qQtf�X���,�+�x�i��t�%#�ןc�f���[���
2�<�� P�3�+�3�8�H,R�K�p\|iT;��L�"�ގA[��`�.i���X��9U�����oҦ��lRx�_��1��E�;�a�i@��C]��D"Ũ-� d$��B��Џ��K7�S��<~��WIr�їBWȫ�er��/Q�0|��k{|`{9���uq���L�ݣ�=�K�&�mP�t��K����U�2��&�"wJ1*��n�������c|�����62�R�>�V{���AL��@��Z���hd>��)Mp��W��uqQ�N�˭�[���~��J�4u�i�i�#0�'.�t�6���t�\\8Z���!�q���r9�D�#�:ñ�0~��dZ�-g2�s0�6����ҷ�aǩ6�].�,bwwJ����
	�yq�Um�Sٓ/�t8��a`��kr+��@��|��v6����B���j��w�w�b�2���BE�)-S`�R�WlL��9��b$;mg�r ��*>lI�,ߓ����Ђ�E�}� t�����i��V�e�kA�{F����*������C[d;=�$gi;�z�P�p��`�r-g�l�D���ΈZ��#QKTk��L�@N�z	J}� ?�c�	%�W��H8J�M֫�bFV���}9���E�Ԧ���ڍý}%�E�Q���?�g8^I.���r��:dwn	��AJ����쫁�1:#),+��#�ׅ��_��:B�{i�u*e�K�+y�p��y�
\P�'����#`4<���TT�	ѡqm�%�*~�^�P� &X�85�a.G��=ݿ�Y\"Q���&��e�В�j#�ʞK�.�XT!QPTZ���{���������,6�J�T���`4�Pɲ�>�^#ﺺ ҆M"����e��7uF�L;�j