��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܫk�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α���N-�`��6����ݾ�FF��eF4��_}<�ےA�[,�|{�?r+-��]n?���A'xin�XO�v⨺��sZA�R4��g�psXdm"�d��Q� N���%>a���k�:_�2���Yn�2�VX�TGgz�)׮QC=�u].?�W�
�T���3\Ƅ֭�.�	��)k�{"3G���z�&bH��A'�'��:��r��0z*C36q��3��$�6�Ț`�����i��I��:	�ϐ�-���ʒ���,+�I���x#c'3�Y�~�����8D@���?QY��?;���`�ˇ���'.?�م�"����{��d�i�8�~	FW������Z�w�;��_Du��[v`C3C���i���{�F�K�K,��F��E�FOC���:)�����?��|_{R���<�ޏ��	x��˘�#w�qQ$[�d�L(x��^�(x����Xvv�w�v�H���[K:�).�`��������	kk:������UىK��C� $uF���$�X�W��~7٧���*�UC?=���
�iT*G4�
�8�ImYE_���\�I��4Vn�uHH��jfT��o���ЙA���"���d�u�L.�D� 4���u:�� ��S�eFO�Cz;�a�na�*v��H�� �|5���"�xA�5J���5�B��zQVt)y��{���T�.�̃w>P��<�}����Zg����m��X����Q8�!���h�!�x�܉ӹ�}k��&�6N��g &��oį��0����?ز�R��f��x�Y�0�|z�(�@Oö��H��E����d!���i��R���Ty�H�a�c_��S9E@ZO�u6 q<�\�����3O��U~�)E7wTA�O#�b�'n�������R�U�H�a������v���� ��������*Z�	8l����MH2��)����D�Vb��TfuT�b5J�D����S�ؖ�����Gx�Ԋ�SEr�47��`�J��:��f�֭���4����2�Υ�����)r���i����|�:���wP�~�F1´B�pc)H�T�v�*�rt��r��HD�6��K�|�d���C*��~���Y0]�i��+H� �J+�1���u)o\+�#��!ȶ�
1*o�|�vPtI����Y�&��r�"I�������IT�^yc��'	�Q�XC �+�W�c�E9���(�ҳ!�36�h��W�A���>���׋��Yaa��Z�%�R�'��d��Q{�M�;�U�s[��)�)�~����JF����(���� �iUa��ϢP������W���r
X��%'��U������>�@��YԘ��V���ZQ0 ���u�7�A{Q�(L���v�k��DL���ͳ��4$�n?@��)�I"3i�%g*��,K��9���"��]�6���L��T�Q59���P$��4��ĢUS�AA�1��وv�8�pr/0#8|dC�ɺ�j��p��>
5s0���%Fj����NXQl`xn3A@q�#d�͞��#U�:���z���ӱg�Y��[2֑����]���-�����t����B�P�b�.L�Fl��z�A�~�)�G<`,�n
Y��܊�N����t!T�)����%��@p��kY�R�ߦ�߽�7��W��o*
F�ч:������`