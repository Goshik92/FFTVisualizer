��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�2>P�~��H�d<#���,5��b�i���-�u�1��GNY����떯NZ�qJ�`�b������^Tc��V�9�_۟�?���m��`2��U2e�� ��_-O�k E�+9�x��=A�׍U�?�S~��t��@�t�_w�ɽ���|/��bR)�c���|��6�ҁ5V�eS�����=2��5W��!�������7�Ɠ���{���n�������4웝��H����m���) �:	�oD3���:���ArrPM�UT+�PXg|A�)Hh�iIT&���k�<qRZ0L�ĉ�m�yl��Z��ґ���|L�k�:�����2RU�}Hg�(}���T���יwB`pq9:��l���q��sNci)F�Bm֠�� ����||Ö$�l\�}�֬]��LI�v����bm�xOR��8���)OHY���h���Q����fc秚+ߡ�+��J���Ʀ��M/�J���y�����>T���E�����ЧM�S�Ȗ�ZR�d�}G������x��jNwZ�
�k#K���c�#���L`�Q݌AI�NZ�ŃU!ۤ"�]?P� 	����/��n��9oS�s��b����ڕ�1S�A1��GʁȗvO"6�ܚ�tZ<���L�sXa�t�CQ���&?�ލ�&`�Zcc�!O|s���K��kMt�M�B�d�lH�p����m;(��~�'�G�Eߺa�&f�5@~/�`N<8�?��3�)���s��곭ە��ٶK���<'+�-���mD��(�Z�Wxx;�tð�]��w4��-Y�)��{H,�����v�����b�r�c�;�T�F�v�ñ��oJ�R � ��gl�@��뵹���A6��&l���z��m�1�!�,<�5XDҩ��Iu���:��+��%^YȒ��AK�!|�j��\QC6X��"���T$�w��� Ӄ		<pSA����9S�8���"�8����&5P-��r>7Jn�&�׀��a�����c,�a��S8�類V���;�<�c`���Ӛ7Ի���ʺ�&��"����#�HfP��7�����m��
��ML�;�
P��Dc���;To�o�1�A�s�4r���D�	U� ������[b��5-6Z1�Wf�^�_�CQ�#:X�ZJ�B��A�]�G�$#�A�AzOU���Ĝ��c(V�CkT�'O�,�k�ajD<Tu�+�J�q����g��25|���C��3thjq4�Ǟֱ	�qž]�r(B���C�:�`}5j�y�=�gܚ*]Z91��� ͞qn��0�#��D�ЛM�4�uj�T#.�u$`A(�Z����'uMy�b�W\� ��ĸ/��F]�U�m��8V�Pk6����z%����$y�I`�զ+��ϭ"ܖ�[Vop�s����B9�GNG�tr���"!^,�^��)�l����(ߚ��VdQ��mI$��>��#3�Z�� $�?%���j�w�Ty���ؽ2�ݮU�uB6*�-;}r�Ǥ��3�lM�+���߷�u��0T���?�kx���k��+}|[�3T�����9^Vy5���<��ۮOѫ���$D��*I�j|�5.)�Qu�t�a�oxȜ1~�*�X�6$�IhP���z�T���]u�6L�y�3�7F�5#�1�#��=E_��cλZ�M,�P��}�/�.A���絸I���u�Q�^r��)�Q���e����f�O�H��,�O�� �!aŊ�rS�/�����H��	G{cT����*;�����)X��D�>��n�;���l�N�Ys���$#���fT��X����ќ�D*�[�4X���%$� �S����P�S����,E%��׉X�z��t�)����.�Oò���_5����rw� [�*�/`���7ǻ�_21t`������F`���k6LY
%n;�F��Sl��@��7ӝ���h|r:��̸+����D{�)z��@�!�"!��
-H���ǷޟI�z<���@��k��qA!^ K�Ž�{~��A�Æ���a���ʝ�n�ۃ���cޘN��6�9{���щU��eE�[7��P�.{>Y��:qD��p�C�^1�ų�w.��c�K0q{8� ��>����:)l��l8��IvD[�)H	�d��W%�1m����O�L#R[��\�� N�C���҂�ր��BIðm� ���?�l\.�c��l����p�<�)j�'�~�{CY���L9o��]2s2�/Ԁ�0������$#�I������vb&�а'�T��w�vh:�N'� ��YuН���"���xE�F].G���O���)
8�:Evf
�x�/�a�,�=r
�g<ov�Ě?X��R�y��?n�dK�?���w���[���s����t(��<���6ϖ�H:��� �%�M�
��X�^�n�P�I����A#� ������r�I�f��9��덅g���s
��&�x����Ld���Ĺ��$�Oj�l�X�\��Ӕ-���^Bh�m��B�x��'p�	 ��+.������T���T>(�Z�b�%M;otQOuO.Y �H��+i�gn!��
�Rr'Q��2�˕��V��X8�m�3X9o�sc�.~�딶Ag�3����H��LƘ��^t�2��r��g���1ۘ�BВ6w���h�>���]Շ���v���#��y.��ݭ��Cx.�Ʀ��Ŝ���o�~Ź{��L���a��XH�nbV��:T7`��N�v;t� �3E�QӤ%�UE���)<?:��&%۾�Mcv.E.����$�؆h��*�zǆU��!�i�!7��D�v�`;D�^��G Q�ڿ�u}?sdI�HQI���!k�p�@�ơ�R
$�x�?��Y�����y��㏘��Ab�Wxfl��@
Ga?>! T�^|�&���Q��KZ�w]�}��\�]	
��D8!:TR��i}G��vw!	f&��z!H����w'�w�*S�:�đQ�?7�W7E�۰�eR'7����R�/�������G�}����C�&wH}��Q:���H���C�	�p�ӄ�q,+�1'c�kv˻�,� -|�eY$�7==�o�y%AN��W���ʪd�Dh�h��?�s���ă����&�k� �n�a$o��m������&y�nw��4���u�x�V����ǭ�;��o(	�
yэ�!ɦM��?������m�Y��瘿�����*����cE߽l������y�f�7��?�oLBTq�J�~&�ń"0�?��#֢�I���8��Yb�c3�	��{�[�5T���fJ�e�G�����}����s"��+�!ֹ�!�X�)jV-��a�א��}y����"�ŏ(���#EL]>��B٥��� F�qu�j�/S�0��$���y�L�͝�ƻ���6�똺��A��!�/�iI�q�1�Aê'��Wi�����0�B6L/�D q"P�~xb��$FVx"|���~�����j��e��Td�+��U�d
 ���eʄ ��I������d�ԅق��D�\b �6B�)�L;<�
���E�������)��)#�ـ�#����f'�X�٥hP²6���ξ�(m�)�G0<�jA53�u��tb�Ҭ65�9���"|c�ۃ�"ͬ`#ɲ��t�$�����JG���9�C�Bx����%pOq�jǡ���6<w�� }�P��6��'��zu�
%�S����u��-�/;�#!���(����&%5K�"#���Xw��s�� &u�l�M�In3Յ�p١"$Y�!� Zzݡ�=Ky�Ec��~�y���re�C[8�^�`.�ϊ����h7���g	����׈$�q�+f'���~��z�\��ןS�I1&w�Vz����>�--[f0W5�i����:�!�f���e�-rX�`<��\v� }�y�Y���E3�gn(�F+?�.�$Y pF��]E��=�\No�<_ ���#�����׎05�����Y����ZCی���b��f��!��x�
,]*+trz����0'qe.wɵ��D<
6�bC����xְ4��O������7�s����{ʲ^E*����9`���N��bﺔ��8���Z���xn�&�6�G��G��C�a�0zs�_!��Pޕ�{q,>\�x�7�~\˿�֙��$C�ՍX���z�S����j�=0ƫ��I�R=_M�k��s(�I��q"�:l�C���G�A89�g�\|{GUZT�@��J06��_�� 8څ����ǧ ^���egѨ���d�o��ˌ�����R����-a�pa9���4U׼�s ���(ylA��>�����m�i����z��Ǧw�
����^�Tw�J��6�\����a�a�_�a8ԟ�9����Zי�k�u[�Au����^p��n&���N���' ˺=��Q�(:�li�	��~�#�tf���A��绱(�}ʳ�F섅iG���I�{��V���ҽjަVd��t�D������#,�B��|$�i�cI�w��w~��t������xj)W���s��ӃHCۗ��v��w)�J���U��A!Z�$��V���r����mY������Қ��e��z}h���|<���	7�O����u%���[i^���Q���{�zf!����$�SV�B�9Dϱ�B�4�l ٭ޛ�h܃����]E77��v�8���#tNH'-A��=�&�ɯߔX4����<2O�ϻ���|T�ɜ�\�5�#a7��xU�I(1�	/�;���R:��b�k+��;I�E������	X��\����8���GO���m0���נ)���ugQv(ϸ�SF�k�nj�� � Yn���uʲ��@��ֲ]������`�p��%���S�%w��_[�����
p���Z:�4d��!���
B�"����EN����$���y(�X��Ja)��"wd[7��Ki0Ma�ʸA���\��_m�5�(�d^���?b����gs���z�d�Z^��&�G�\�܆ѳ!�-�J��$�Yݞ�Σ��H�CJ�<T�'�#��I,�Ԉ2f��Y���<���OB6z��_DģJ4��R����m��:/~ڃ~
����!R<TP��(�����C��X���9�du]�?3t�c��
�]������U]C���}��=������������a�����[��X�	�f�I�N	�Ku���N7}�w�{�P�x�����:�S0H�q6t|�����5�}	��*���s��<@�t���N�̀��-:3�_Tqe���辙YBD�#:��7�
Jy��d�XPN�ė%q�U@$�YT�K*��Ã�b6�I|�u�ݴ�;mO��^8F^{��U�U0�@�+�=aQ�Hc>c��mT������ZR�����.$��b?稴�n(���"�]7`�&8�{(��M�$.+��Q�a�`&�W�3�H���Iڳ���&�y�fs�q[�|B��or�ެ��ERs7�&�P^mJ��S_�:�z��"G���3a�������-�mA��} <�VN��)��������/!�}�;C�J� ����^�u1�('�|_���b]���O�����\�l����4�/Jۨbyb{�]�.s�"�w:	���J���3�6.X��؍�>�=FaG�[�K�w�ܑ��h�uM~�5���4�1;A�R�p~*7��yP���`ty���\�eύ��7�k�qL_'~H_�4��;�M4��^�k���Vk�k��r+��v횒��GN�<�"��
�CUډrv;�y�-�n����c��ע؁/�ː��5��,o�V���� �"�§4y�G��т�|sYI��քO��!s=$�>HrXc�זG�kg?�U� 2�Eaw�ˋ�SV�_�h�o;^�5��Paj���0D)�c�K~~��Oؼ:�c ���#Qd{El{�C]n�L��ߦ�q�fsD-͊v,4�sU��z/�i)c��ӥ)��y���1�����Fuh��k_-X�2��Cs�f��Q��{s\yr�-���Nra~=J]*�n\'#h�4;�a���¡O�&2�K#�1���%Kn2�y�A4�ˑmze������Pi({=4q��"����BF��}J�� ?���!8��B�`�"����nH9w���s�HD28A��!�����TUW�� pa�Hr���-rfV�iυA�����ݳb�}&�Rrj���u0F>�V�«��<B��j���`�h��,��
ma�d�-T�J_��^#���{PQ�ѫS��^��������sD*�E�(�	XB�-	�i���VD<��*��
���>-�@�C�*�C�<q�����wl�9V&�~�;�5l#ئ-�I֏��5�� [kK�{�p�Z���OK ���L("NcKj��kfy/��p	�$�ӝ�!-��2oW�y �4d*�s4���\��`��	��t������oQ��=k%,V��պ���7ޣ�H~<�>$���4�k���,��iCb�>S�Q];M�v��ÿ��!�$x�d�o9Ө^�)���ߗR�]��"�E��U�.�(��J.���4�F1)I�7��r��\�<$��(#�p�e*����6�~�*r��z��Ѓ~�������t5?v9�/0K@�ĕ;��&���%mr��T�tn��`61�S���g֘��02����v�/�<���ul``�;���n�N���q�&1���?����`����b_�[0 P���f���r	D$�������q�v�0��>�/�c��jޯ����x�ɦ���A��7V����D���z�^��=��i��	�JKy x�7?ʤ_7����s�' ��9h�P鱪��}���j��"w����}�������V���ʸ���
?OC�Y���6��YB�P��X`�`i�Z�(����7��tPc�yX7�*�z��Q�!U��y����r�yU���W܏}O�@��h4����g�:V6Փ-�L�tja�.��rm�X�I�����hl����+�`֌+�!}�B-�\��z�c�cRs��ѲcJl6�'�lC�--��a*��v���2o2�F��_=k�#��,�����@����ZK�'r)�����^�%�.(��rp�� ��=I����^�i�\�`݉�bב�9(�R����b<��(�	r�Ì,�Eh�
3~��P��t��I�8�.����\6��5��`�1.�9<���O��O����C�np��p����Gq\���1':���
%0~?$�����~
ٸَ1{�ګ��C�5�|d����a�ǾH=|�_p�w�&_s���Uػ^4�q&���#eH�4��Q@]&�L ��L�|���e��x�Gd6q
)Ǡ� ����	��ҍ]چcF��<��r�E
�F��(u��+T]���a��@���Z��et��).���q)h,���s��H}m�p%r����Je�AU�/��Hfۯ���f��rQ�hץ�%zB��.��"X&"��p��m�,e&���]�sˏ?D 5�j�I�����c`� ��(���^��"��(�����}G�<` k��K�Rh{� �%�u�!*pǙ�WlҏcjѬ��Ű-�WI0�c�Ⱦ�8ϐR�a�]��y��㸙j�ؠ�s�#&٥1 P�fέ�Z��45%��;��̻��	�N��αI��Oߌ%�!w1��ꚙ����l���g"M��9��y��8�	lWT̏����_�� 20q4)5�z������_��uN#����+6��Z��<���$���n({ЧƄ�a���6����� �'�һ!g���y��1�y��!HkJp�����HN!�8\���� ��Γ{�`jW�����UPFwO�/NL�*r�8��R�R Z�F�E�/��� D��>��?�K���P;�Fj��N�sJ�Dhǒ�Dӆ�):��u���v� H�6�3;�_�oP��J~8b��R������Ы��F�%�|Bc�6���¸��w�er�Q��fq�R�㦍�6��!&�=���C���8!<��kI�3����{�
�M�iV�b�z��A�j����x#�jC i���0�oΕ��J�����n���Ɠ�
鴺(Z���D�wgܜTc8LM1�E����`@y(<�G7,I��֠�|d�u�vnp W�d�DQ�k����/�ћ�U��q.�ʸ�U�1 ,���^��is?���ǁ�'�ߘ�2�.��rn�V�+ �Z	�gRo:ZoC�γ����zr��{w:���՗�,(��Ǒ�����WD��9{:a;�����W1�v��N{�8������xr~�$�o�l���w���*j�%��<w^aS1�8#n6�}��k�;JF]YA6�ӊe�F�H:��^����{�;]�1 T���L�{��р"G���@��'�ݐ�����=	u�)�4ï�X���+�s�s ~�)s�-g�:��]����d��jU)�v2��� ��j�sǞ�Nx3�Uf{����;&Hq���@�A���;������8��o�4U~7�ժ������9^��bU�q�t�ߦ�l��}�������Q}C�:��xm9!�(8�H#�:��M�~�)F���������K^�D�*F��<5�cIQX���5U���e�`��U�t��%f��l�ή��y�-����ޞ`W]�h�4[;6���yg�,���?~5g %���=y�8�I"a�����q7	�^�x�"�j�K�[xI��G]K�_N�;�O��Jq��ټ;-%̜�e��D���P�� ?�����E��6c���n�}����+�L~�2g���ůw�IT�;�?Z���4r</ܺV�������O�D
�(�=�ۜ���� �����JKT�d� JVh�4(�Q�9_6]��lv�!5<�����e���f��c��^L�|؟�)�E<���g2ǋ6q�ۢ"*�Ug&����5aEA�:v���;��NId?PKz�ϓ%���o�%g��1�/V�?�+��U^.�w��/�P��b��J�o_�O��>�O&:��%1���[�x�n�zh�0Ϫ��.XQ(F�ޓ��B�]�?kux8`Κ�&Y��>��aZ}����)S��3�^'qx^B'����pD� �����@��j�Kyk;�xe��j�
�҃0��7@\�T��\0<��(������uԽm���n����l٨���w��D@��ޏr���*Iu�
�U3gsƓ&�D�W��G&�H�7?<y��ZC��:�:rZ;��v|9)��fW�C<�8�e ��4��^FY�Ɣ'ӋX.zPH�N�̿1cVr�Cl��l O�t�q|rAa��Or�A14�Eu3��:9"���_h�<Z�2��b6�ͥ�C?�Vb�i>#y�ϩ��� * ����!Đ&z&*�tFU֏�y�ǫJg,��U���a������Ԫ@��I@)�j����:Ԡ����!Z�g+r;�骱����ӫӼ�vW94G��T�;,=+u[��pF�����.e}9Cǭ�|ϻ�~�&�����iK̬��XM��AKL�I�.�#B+����*����@UI����1u�Oܢ����ɔ�=g�+�w���@Ŭ��f���A���l뷖��P��L(N\��_���V��N����K�c�cZ��`/�pέ��;��R8�X�r���d��N�ήB:��2�(hK����<��U���T�e�U��������1I.���(G���E���:�$��MѢr$�}��Ł��cr���ى�=5?z�<萩ݬ��������zPf�Yց�C�+��q�ϒ���0�J�j�Y`O�.^�j��� ��&�S�A���'���-�����z���������K4ea�D	���>��P���X'�\���ݞ�/�Sg�D�J��1��_�������cu?*��~[=N���'����h��`�{K;�	��B��&�Q���9*�(6����]�O>�C���
yiޱ؀���Y���~LrT���)k���+љ�WN�Pj���:Y�8gC{�ȁ��
ph^�Wy��v��8@�V�M3h�e�:�݅��X�J��w��`��c�m;��Ε��ze3P톡:	x�%�+��+}������Ő�Cd{n��O�kC8qCb�s�X��x2z��a��6:�W�t�,5D������hƹ\'�(~�o�o�~�QO�B�'lx��<M%.�	���AǑb�Zw��>��.�{1"��ڵڄ�ډ&8uE�Ⱥ��6��dCE�S!�Ip:����@i���g�b���x��Cy��%S�cNl�o|�8_>&/��-����!� [Fx��keVA����kA�ր�qOp.�w�⣘c$r�waͬ�Z�B�G���.��=�����`������Y�&f�V�����"u!
�ø���_%B����ݝp�}�m}�M�ٔ�v�H��̠e��o�?p�ϐ�#�¥~�Jz���i��+?5�����������9D��4�.�_����`:_\Gs{��T���ʷu�O��i��!g��{#>�|Z��?��Z�ə�E�p�Ҫ�S+�e�����e��tݼ\d�"��P�8K�
��b�AB8�0%9�@�>ʒ��A�MK��E���юփ��%���l��ԉ��$z;]"�f��mR��F�c�̳Ӳ	(mi/��*.o�r<�����WfU� u�{���:�jߓ�����Y�]ud���#�1J��t#�yQ�d�?�_-���T�_�^1��cF�����s#�lL�0��J��?�*k}6�-�(��A"S�ux^�_�[�-sN��/�b������sќ�"�}��n��/�*`KQ���L���7�g�k}|�զ�r���\�{�:��S����+}�K�wޫyR�(��ҳ��جn֟(�� *�,\�| ���ғ۩a��uN3���xa�U�?h��5��ln��o��L#h�hM�������^���u������#���NoL�u��?">w���2�o�3u"����n��~� �e��܃�g"��w5}�<
����Ph�2�FF�	Iv��`"}]͞�W�ܙ��x���u1���V��uD�%۟,	�jV�RL�3D2�dOeYa[{}���F�����g˿��{� 8�Y�^r�2�4;6CAY��ֶ���=?��R�ن^������{��K��/��W¶�B��������^~@�l+�d�X��6��%ݿj�ý0ty��	9�%`(!�v��37�X�M�3�=h��p�p��lC�DU52��a L��#Oa�쁯;�Lyˠ�ދ��lC g�5��/�(O�N�?e��$ߺ��o�*��-O���Ps�N����I�ε3 �DQ��CzAzF#�z��o����((�s��O�f�Z�E��i�>/��55�J�vz�!fY�7�/�t���<p+�å��߁,G��_�l.��L�C��?�������!�^Cl����8�s O�}6�� i��c���5
^���!}�؛P2o&��iUD/���g�F+���*!g�SO�t�̳5Pn팒����!��2G>da�*��dkڣb��D���)UŔ�Vuu���S�n�5�T�� ��6S�Px!��4�R\�}�j���}�H�t�֕B�~�������@��1u���Q��sP��ԛy؎��/��d��ه4�gBc9�N6�oo���%�׿'E��f�j�uզ���Sޖ�e��A��:A|[BEp�Z�^҈��o����x9�M����ʯ��iפEZE}h�@hx��]�����^�=`	*�rT��阸����A�����	h?#��!pYjD�Q"� �J�`�~�Ɛ		)�E�"�w�
UxSx��E���x���ʇJ���DFR�ʐQ�����P(3g�������M�:~Gy�v1����Ri���q�3�e��v;�N�rņ���Q"U�s���*����1fe�؇"���;�<�?&.�эF�35KL�[t���8O��.1��ć5��oa��̺>���F��ZގO�S�f�=+7�<͐�s{�s����+F7�t�M�R������+$w�o�;�Đ���m3���ҋĖ�O13�+[����vQA��|2Ê^�N�u�g��T���������E����ZmSa���S�������f�^e��d���X�a�u�O�i��d���I��K5r��z������5��3�4ڧDك`�iؒÎ��u�U��3@�r�������f�	�
��r��kW=�9;|�B����sՆ��U�n�P�Fb
,�@��(�_u�Z�G-�O�M�\��QXж��]����/��"̫Ư�nM����۟lNL���f��*���q�V~Q�?E�d+K�2������MA}��{�0��B����0r�����K���7`��T��x�e��7�ܳ	������""siS3꺧=yd�FN��7u��*�%�7���k1@n�1�,�������'	���+�Z�M������v�N�Y�"�[�f���L��<}O���yr�JY�k�W�ܜO��ΣN�f�*{�z��[�Ω&�nW]]P��!�.��0w��Z���ȹQG{+����u��@˩�`En+Ru7$�V��tQ��/N�C
�����,d�f�P�D@r�84�M���JT?�Ӧ8zj�Z�T���Z3��������>�j-;�a���gђ57
�J�`�G�GZӣ��o@�?H�:M��gx=cV�ftM�@���Q�8I��x.<�Wߨ%�B����l:�5S�Y߬��"U�P�^�M���01�F�w����ݛ��2E3�k,�#w���Y��׈���Eũ��fZ����Ko������n���3�G&��r(?�sb'wɱމ��!l�q���=��Xt�&6}πVf�u�bc���������#n&� �di��
�lS���AT@�ͮ�SӃhF|[ďy�wK����[n���5w�E��Va�_)k�@�~y��F���+�(_I���L[w) �Q˟=+���n��ɔ��&M��������Lm�|����_o���۳!���%�T��G�,FH�jU��'��C�$.C|-w)(֨'�z�X�?��754N�V�d��x��%�9�T���b!�o��\Ij�����f�vӈ�u��XH��&K����BK���D�����_�tb����p��<>��\C��4o��v�'�~�l|�e�T����k@*�U�<�p+��I�pKz@*̈�->d#XS���@1��{4�z����@�b"^~�1:���	�$��b��}ƒ|ud=@��p��v����|�?;6�@�-�.�h�]�LS�ۙD�#�x#�o�rIe�]���M%��������m ���+��*����J���/�rn_P?E���8��h���W���ˁ�|5 E��J5ږ����L���f����+����x��-l֩]>$ ��a�t�Ξ����|@v^�;9�����!\���2�}�x[��PVCk��Vq�9�`��X�\V���*�R�m�&6������?Z(Z��E�~�϶DF�ۘ�ɜ+�Yb|م�Bkl��J~|�,f7�c~~s=@�!tZ۾���2�~�P�dUA��7��Ӿ�o2���3�W�cp/�\o-[Gz8)�Z�E%O�&h�Qq�U�G݂A5���j�!v���W�F���S���,V�[�@���N�B}RC#1!B����^��W;45#������2�/o�8����>S��Y�xb�f_Oz>�1���%۳l��L�5f���˂�R���I"|��C��i�V�P^/{O��������E0 }�4�By"䶙G�Ȣ̕ C�6�UQ/�z������#��\�)�A���C4B��e$�Ҧd�䯳�(1��0���|�n���peF�YA��~��(�S��U#D���W�4���ǘ[xh�\��Ķ��hsW�s�,8������*� ǃ�_5�;Q����jM?�ez��?T=҆cTt��<���/jP	����w��P�eD'�����/j\ua���������J�k�wuJO�z�?T)���Y��Q~��#�B��z1���4<�!>�|O����� N��E���փGP_��Q�8�u�o��5�n���^S�M��Z�x�~I"_A��p�ʖ�R�n�,������Y��3�$	:�jPŠ}�w�Q�����m�H������ũtS���y��br�x�p2�o��¶��G����S.��Ng�ڷ�4�#4z�_Et�	���'���`@�\��Z=���|
f����eM�W$�١�����\Z��K7�J��t��|ԟ��Я�G���i_5�$����}�gm.��j_�P�L(}�����ͪ{��� [n#ݧ��fb������r�Oh�S��1�c��%�dd��tq�n=}$���H�>���W�R�=�]�a<���W�<�t���-=�oc��>0+{!!6��ۓb�?�?�˹��*ɼ��"�E��JK%�֎8Ӵ.Ɯ��N}֪S�|"�J��4��%�����~Q<R!~p���pn̛���u55�h3|���Gt��=�baK��L��ہ�!�[d�~���hxMUZ�t��5R>�eg3E�M��|ܛ%ҿ�����C��/#3�Q�^���I���(�aa©$r��d��o~R*���G�9��fo1e%��5��l�������i	�����D�1�::hk/��x����,�5�Py�N|�2� ����Ii@/��49g
�hĭ@]1N�B4sH��Wg�DU�P�E�ڹ�g�]&hd� ��^0g��	�ž~ڳ9�q���	l�2d�������G�w4�H�1��F?:�=�+�M/�k�j���y�o�.��M�a�&��S�?�u�4o�KD&l;��;��c�p8\Җ��bcbjEx������!�aR��R��ٟ:��Z� �n�S�Գ�Y��l�[�pi��؀qAu��MVM��9�������)ԑ��|����'�o(����ҍ�{�����T�_�{m{l������a�h�' ������% �v|�ٌC�fg'�os4���K�4xp�n9÷��,Т�G�=��83�`��_~�q	��t�Fx�	�Ⱥ�#���)��*W�ms�cU�[����=o���jR�������3�`&��%e��H[�=I�n=�ǉNv�zw$��/=�}����Z�O�5���6��V��=D��K�����f[�z壜a�Sը���ދ�'� �^V�-s!�%�0o��U#>�q�
�}M��7#g�b?K�6.A@������m|���om롭���%Op?�Hx�������ﰮ��S^;�k���� >X�٬9�h�T���E��?h�N%���pX�y��g��KII��p��������>O��,��Eǈ�S�S$Xh~dS	��P�����J��g��m�%�^�/���k?���Di$s��0���?Pik���sR���z4����>K#�ԙ&zu�\��FY��8n΁n��Z5�+]g���;P����B��hl}���~R�'K�|K�ҋ�: l�_e�Žd��,Oy�g3_�kTU�ؗ�:H�Q��S���r�!<:F�]��w�V���v����}N���eA�A\{�����?]���E4�U��gqnD�?�c)������QX�"]�❉����Χ��X�����C�H��h�f�3�ٗ��a�8�ش�����t�G�L-�4�Ķ���s�R%x9P��ϥ���v���-J>���g˾�z����X�����o�48x2���Qa��}���ݑ��^h�x����{�q1�t�c����4D��݂���L̫�_)�)�Y���/1���I����n���l����g�#uTy��|˖v8* \�IQMh����մ���xD����6!���G76R�n5>��uj�B�ޙ�r�ZJ���٤Q����S/x�M!-ك(u�Ćw���s6W�	GU��w<~�����Ⱥc`ov�j���pB����@�4!�O4�RD�ԨE6}(Mܢ����9�ǈ�?	q�Wr��-�ylf�9>��o|v��%o��5TE'��z@�:�cT�[K|���U�e���,̾�U� 0r��r��|�!�նF�[Wl��T)�%4x�\d�#Q���a�iǌj����\�u	3Ľn��!CX�t�ov6����Ӑ� ���Y@��B�[S�ՑID_�����IZ���R�ak�6k¦�K@�?�z��r,�D�\`�*�\�)Fu�-��7&h��\ڀ����$�٪)�U��|_�Fɵ�Ɩ�7����F���{�6����*͊�6�H�"-	&NȽ�1{�z�}4f��P���r��/P�aWXi*��R!"&M�̽)��7��:�:Bx�]�(�����ĸ�duC>Ye�it����6�y:�?��=n��%f[���Y�9���1��m#[��M2rF/C��r�
����b5༢)�A�%�n���Yo�Ӕd�BS����Gm"�9T0��̞,���8�R�������kl�K�B�F����G/�3�aW�|7f)�}�L�糖��P�q@E����a�YNF�L
Jb���K2�ͅf�5�>u�����k0�P\��)�o��H����2�����7�Lo@����G՗߽��O�6�hh0�R���Ȉ�L5m��vb��9���&���+������Y;������&BU5��;0�:b�������=9�צ�
��X]����T�j�Ib��H���Ïby��L�dW=�^Av�c�5x&竏k���t������W,�u֥mH��	J�S�
����0�`���[n�W.%����\ȁ` ��7A���e�'])˗�T�`}-yE�{���r!�C���g>z���Y�D���aRƼW3j��y�i�n��l��BzL&���s�����;�x���x�Bj����TcB�&�wB�Ո��G�9�
?��>Lg1gkc���G����������
y[�>ϖfm�b��r��1����<?�(�J��)��#X.o)T���s<.p��4Y}G�u��5:��'�4��C�n3� ���^�o*m�"�0�SP��
�/�+��G�P[�����eN�ڸQ�K�5�<����Q9�U�E�O���zx�K�E����`ía�uH��E^�t��{'����v|&���t���/��TU��h�C/�˱�O��8&�1-�ހ$����P�;n�(�O���<{>:�B���Kr���F7�
��E6|�7�H�-N�E��J��� �}�R�W4+�f�( *�Ғksj�7��2J^g܉��&���xjE^+޴W㥫�����3�)�k$my:�:-o~���U����Wg����"װ�@����qDB����9�u���M����NY�|I��W�e�"���F�r��=�y|�x>��ڗ9���ui�'�{틦ζ=T!R�\�h5x����DJ��]�	7v ��y9DG+	q��	v���֎[9·���G�7k��U�H'�� �rO���j����٣~�}��l$!���w�o�Q�nQ<S�L�ҿ��1F^jʙ�4s��'��nbp)���u�I�d�Dy0�M3A3����#��=�,���g��V%}��� !���|w �T]�A����?�g2H~	��R�8%3I_0��>�h���UԒbz�ܦ�T�$|J2�{Q���V�����}�">���|DN<�톬�Z5�Y��bs̚
da)֫B. ��k�zHd�5jj��Gj��
��]�a
A0-���@xc&t���J�7�'m�!�TH�<�I���� w>|2�d���o�0���xA�c��6:�f��B�P�?��s�	�w�~�Μ�Ўi�V�����z�T��Յ����������U�~N尝+� O�t��e��ZǠV9j�V�c�pKWᇧ�0s'�!�K�@|��0���+�?��"���e�f;{���ϻ��Y���������5žc�_�v�^�/��I�΢q�2�5�i��<o�&&\|��ٕa�t��W'�I�Z@o��k�ʡZ�}?D,m&�����9Jw�=��$tƅ��@3�>�}��3�|���#�޳~s�)x�=F`��~
�`ʖ`w����6����0c�⿏DK@2�)�.)_cQ����ՠ���J��`b��݄��sp�l�4�I�+�sN�|Q*E�}�{�[��s	#��W��I��ņW{�֮�J���K��bL��>P�FJT�c�F�a��uB����� ����hɵ*ii�&�{O����ێ���|L�#���K�w_@��Eݳ�v�S=���q�	��N����&;릿��������b��[hb?ƕ-W�$�G�ezj�X�e�{��~��	�ya�%���ŝ�>jC�$��a�Y��Yn�s�����3*�Cw �E���>k�6��R*�5%���_9�4��68�f��p�ߣw�L��c����Y/�3�D����Y�s�`ح�O�^��]�fj��U�τ:e�?�R)i����E*�J�G̣S�9��1绒�?���T�\�e��c�pP�%֤�L�g���)C�)�0`q�a����}|�7��L�A|��
�̷nϧr"���2���Ǯ�TT3~}�L�.�@��G_�3XJ��]��he:��^Ё,�ؐ�;ஙb���q+�M��b�T�:,j�"���8C���4�`���~2T��S�DK�������c�׷��ܫ���^��E��9m��ߛ{��п�ާH �1�ːd��/#�Q�1B���ɤ�F�dL"z�n.e���`��l���r�sX �E����_�^�M%�U�������T{|Ip0;c=u���ϰp+��� ��b��WhjXYL��Eh4>/����S��c�n�|�qU�O߻�iwOm�XF�x@�u"X{g�H��v�������B�O{R9|i��[��!�޸�h�xo�� �cJ16���B��Ve�����ԉ���J�c5��F���=~yG��|3���CzZ�ܳW��B�:�?�XȨ�$�-*hz`*�}f|$r��;8p�)ft����7�N#%�E���܋.��D�Cuy���*���<���W�-A��hʴ݀��_Q������'��Ijnۦ���}ŉI:���k�>[��0n�L몙@=S���&�R���n90�c�h��n���䧢
I��3���;+��T@nS@-�pZa�-�f�^*0���Z9=~�%>�
��.�i!�7�t���K˒X�?K l!Wy��V��{��2��/����n�b8�8}����<_}�㪏����F4��"v�;͑P��q��[���n��29Nsi�r�C���tt��]	_p��V� l�.C��e:��Z��P	������s30���W��#�����/o��Fs�eB�����
e-�;�0����.Ő��f����IC ��{�|O;���kW5h�����]�J.D��[?�c��WȬ��A+P��5�
�����rA�pUvţD+�f��<Q��n�a-�hsU���>|������hu�-栅�$�o�z�%��ͨ�ߓ�|v|R���6ʨ�u,��� ���3�'�$�ĩx����?����'�V�Þ�s+*�e�0�K��g~�Ѹ�2��L�k�GW�Iv���X=?��j���O�?���{��ʪ� `>���C[�U��U��}�o1�{�#�U�w/�����u@�7d7��kY����r/�Va	�B������X_T�/cշ[�	��<C�}6��"PL�T׫�!�\KM�@�����OA��L36�Ⱦp���FΌ�iF��<�{�u-_���țruOc�.�Iz!���Ѳ�W�9g_�r�o��T��l����7X�B�8c�B�6�cd^@��Z�gt���w����0�U,#���t&J��l�Ǫ��u���ON=65Q��	
���W�u���Vf���E�V�{�Y1��/|�<4�er��_؄��i*��}�sDB-�"�[�4;6�T%_���L91��zQ�w� ��A��w�,��-�x'���x7��ϣ�MYh�$�Z����tT�J��5|���-Y��4�,�8������}4A��!�"w��O�E:z���I���9�ʕ;�/�^N��҄T	9ߒ��W�p�(ԃ�bK�u|��ɢ��4`6�����G��y)�\�X��++>�B����0�?1n1���ep.$�X=�'�=�Z�65�Pd��r/$�������;�2UTaS����^��r��;�=�7��A� n�y��ͭ�� ��qMLz�Q���������C��]*�ފs��j������H��J~��W�+2��*�*��0p���#_"�\��/-��Iv̉e6}'(~#K�=�B;]i덩D� �y�hC%nYJ���O�-M4WU�?	�G��9�Q-��%�|U�����
{�U2���?����j�@��S�/z����]�/{Fq���A(J^���=�G��XS����M(6G�2)��A5���1��( �O���|���a�W%��$���i>�7$R�����cڠE�T�΍)�7��'��LV���釵0������s=�9��&�̕˹�x=�@q���K��O�m�b���]�A�v���ZH�%м!���t�R�Ig��6�B����8�'\��RZ�v(Ȋ�[���I�Hs#E}v�0��ƚ>��+<��7ߞ���2�E>W�uc�0���)>���~<0&C��t8�|e��h�ʃ��1�bH||��C`��`������۷ˑ����W�━��Bs��N��&.&�k���@E0ѵI,�V���z�ud���b<�7{M�"�����NԒ`��@���|�}8�v��'����c������ẙ.^�y��_=�dq6�[6ԥ�2�]V�Q|h�q�xLT/�*Q�Dr���������C"e��
$T��?���a	I��jz��NFƓ�K��o�5��F��A�@������9\���D��o!�Vm���z������?��*8P+�%����@����@7�V���(�%�J+�*�)��P��4[�ʺg�%3�V�Xl����Y#�OmwЇ4;�yCbV���*I}]�ê�5uc}�����5���2����/��G� � sF0�����>��P�sl�)ITΫfE��O<e	y.���Z7�5[��J�0�6�z}�m��x���>�u2�x+���S^y�ei ֞9Ѯ��`���j�-�4�Τ���a�.�~�ip`\'UJ!�E¼rc=�>xD|]�&�7<.q~�i�Vl<\�P�a	�=��*�9T��?��ݬ��/��f�
K����LK�S�aˠ=4��X3�O��x�uN}�1�ZEB���h�)�~%��g�݊<��ɢ
X�L+�Y~RÂa�Mt�|�]��\��3L�J��5���OQ�� K��Oo�9��2q���ᠡm;�Jy��h�p_���m\��g�t&a��G�$�����8h��+o]�>�$zD���ݒ�sw�4q�K�,g$zd�i`C�F�O�K�rmc��j	���m2�f�n��Jٶ���7��r��h�^*��
�>uQ��"���ۧx,��Hmx��yx�-�4�n�`kܵ�88Z� s31���a��R)���
���^��A�Q0�-(gs+ܮ�<ʖFQ��;���?�פ.X��	5��*����\f���ϲ�(@�h��l;�C��l3±���8r�#�L4�w3����2so1��E�!){薽A[\�Yhx��
w�KtY~]��vmkQ�ۧ��@�q�63ڠ�>v�q0���f�sA��{ى��Ҙ����ʦ)�N�;c����{�hژ��?Y���T��C��cS
�`r^���8A5c�q��Wc ���
��}}v�h�\ƚe��߸GwQ��./�.E.���+��5�6��?Ҫ�v�T�m��/MW얲[��ٽ��!{���ݘ�֣���e7�H
���[ID���
��_[�Tx	��Ų����R��o�m�$W3[n�M���a&�Fi�Ёv!���|YI_^ZuxX�L�*�A�� ��Eo��o�{Y�����I�'�T���t�EM�H<Y+P�d�!:�I�4N��o˲.� �8H�q�0�ihԷ�Z�p��y��{qq�7|+ݑ������m9'`�Y_[�	MGc��Id�Q��;aC޵�ӧ��`p��|jS�'�r��ZeTU;S���~�l��-/��k0%� ̮�I�����f�@�-��Ў�1�x��J�?���\ܷ��óRtCڏz1
��;O�[�UnX։���٢�����I�\;�%<faI@�T��䥱6D��5m��� EIB�z��S�8�D�=MQC�3�6%[Ka��`�L�7��?�B�=�s촅i��0U'bK^7���\̴��
�C�����������Ep8R��-���	��Y��Ѐc(�q��(��C�C|�Ť���ڀ�?2���o�2W����tH�L0�azz�(�o��� @���\٧3ԳJ �y����] �:.���ߡw�:��yWyԚ�F��.��S���X���R���udc�K!q>!wP����=v-�Z�s1���ec�K�9x�9�+���F�؅�ub��6v�}p�Ҧ��s�]���su3����������!Kؠ��*i2�dd}i����k:�
VĿwZ������D���@R�6vjn�E�,�`�ғ��KnCzK��gC{�\�3�?ulji�$�����)@F��}�$�c�5��:�D�Bȶ�ڞ�zߎ�~;��OG�|���� �\�>�����2SO����OlN*�U/�U�k��v�6ˉ˯����w�:�}z���m�~��"�ȱgXI
Jn�	��b�Pn�i)��H�4*%� h���0�pp�gOl���t̓�����a�,<;q9zDH3v�N�c�"%���'1#�b*��󡶾���:�Ĭ�7H;�2��`�D~���+0��=�ď����)���̅��2?S�����'$�d��U�za��a�y(љe+�������f��FU�t��|�u��=�9o�3���l��m�qF2��-��]���w�W���Gc��;B�<o�8��Nx� X7�~§��W�b�~˽A���l��F~4+����_A��u�MQ��Jp�:�v*O5��t�9�R�U��cj�\hxӊ��3�"�[�7���׆s#a�@5�?�x�L������kE~$R�uS7��*���Ӓ�{�tP\�j��u&߃�7~B�4+=�:��L#M,��"��JA��4�J5�"���Z��rТj��f�ca'��:-ɓqh�	'm�#= 8ԕ�V�Z������$XK75)��� ��v$A�wǴēd�Swg	��j���7�����*"[{|y{��y�N���1"5��]Xo��-N��)s�W�q�;�Q���6���Lh"[2
��@O�0�i5v�����:Q�P�Zh�6������~�9�e6
�Ȧ�7�DM���{^��u��E������:�3��7� ǀ�+�!�P����=|����i3�C�;3�}�24��,f��>��°��X~G�GV�M6��}R����a@Q���S�|KxOvÛ�0�f��/|I�9��0�-�e�X�J�,O�>iM����y�n��r�<5��l���q�ٜa&�2��}onb|	�mPRwu��u�-w�
�䮑�9�B�A�F�GW���8b$X�]Ǟu#����R^fћ}��QN�Q������3k��>r�:x�Csn'P���꒐WV�;�|�*���X���|����-����ن�o�,9��~��z�
�NЖ݃�b�U!z���]>A;يcb}�r*`���4�!�6��ӆ���Zz��%L�<s�]����ʶ�y�`�������nłI���/��Y':kH@�HD�Pb�PD^<"4#R;��S�W��k�^X���w�	h�ܤ��.�8	ܓ�<?}Dc�j6����Nx��tcc��yœ頍d�nM�7�e��k	�lWR�:�f��"C�(��_�:��@�^O�����R�;�fB}Ѯ
��M{��Z���G�J�:`���8���tP�lw?��2@r}>�VM�L����D�;�S]������J#��lA����!R_tg5+Yk�-glФx�>^p��r[И7�4��#JPGx<>.,L�޳� Aj=���p�^5�O�����ϒy��T@=_����8�ٕ7�&����lR�"���V���t9�=e'#o��,h��T/.0  �u{	�^��al�=�Ϲ�i7j���R�C��eѷ�|0hۺl�e�����9������HW1}�5����͎0�z$�^K���=�!��j}�-�sb�YY�[�\>^���?��䏽��B3�k������X��"߼I�LZ�ƈ�G Z��߅�]�s��]�߻��D̗��2A�W����@���\�i���'��Ee_k@��D�%e�ɥH9�Ԅ�:2�ݣ�{\�;<fj�j1����!��)����S���Q
�l���!Ƴ�m`G�k�p�����9D,��|�U��x���=��PSO8�ݢ���W��Mh�n@z�/�,�@�l�	=R�@F�AU9�Ȏz���$l��z3y��FC�d��o�x�܌q�f#'��{�0���l)u9
�]�WdZ�A�:'�c�r��.>v�<|$���%�iCA��K]����ι�����g�K��jӔ*�e�쿽��lI��XNo@����<ܳ�7Zp[q�b�Φ3�ߚ�.U��-0�IhqEC�n��\��d˄���&�{�[���+VT�������d�U� �O�8�"�.���~��x�v��R��(J:UOJ�T�㋪<�,�8VV��4�
5u�L���V�Vǝ���[J��<�d	��K��������  ֨>m�k,� �̚/V����Y���`>:��bs��Tj@pۅ�w�<�Yrq��sA8���z� 7H�����y��}��}��,�K �;��k)�+�%�A��R���"���T6D��)��U?�4P̄K�d�c~�E�^:7;� �?�����U���c�NDɢ�F���o
��bް��o"�^���@1��L����D*�|�֗�,/�t���A�((�T��Tq��;�,{	6#�Jq��Xb\���֟�"H��E�%eYP��*���.ߞ�M��g�X�1��	�E2=�&_�I���(���vo��Y�����Z�����m�3l4�U[W@yW�u�b�H������:�b��nM�d&+j���H� _��<�q�u��F4i��
qö�����i�b�}����q�$��p�NL����WIP���ӱ�+ˁ��	D��QנikF`�|�%+F��* 	���l̳�jڬ�?�XgiP��?Wx�Q�hC؏N� �8������:�$1>�!���ey=B~CKX�����8gs��rг�]�����cH�C����2��	G�X'k��៥}_�p^.�fiw(���� ̅%ʳ����vQ�vS�?K�ʗ�\j�8D�ݚ�/׉~@e���xm�;�����,t�Dd�Cr��k4��WH{�ӜQG=���5Z'������iϚ�fH��V����kk�g�DW�lQږ�݃/�`��Z�9X@�j#�\k>�uz�C憎$ �tPI[��:2:-N�D�6�D�)Na��O����5 ��l�X�*��'p���i�W�/�,�T������RG���GZܙ ����K}88A2ߥ�4B�A/�&������G���=#�3��ng`��F�M�T.7�d����H�t��p8�\5�T~*1�gj+"2���������C�Y���w)��0ls�x�E��>�U�H�Rǭh�`�8��Wd��w�LX!��o�f�R��_�ؑS��mn�}ҮYu:���#d��FU?k��,�N7�ڭƓ��?op��jH�r��RG5�*��Pl&�&��Yb��.65�Ko�*'p3q��3y�Ľ��H���������9��{r���m�Q�%Z�~�v$�P,i���͘��� �_�\ȜIt���nǚE��Q��?X��i),�Z�Y�S*���GgrjـZvM�/CJ��IU�D�b��Ql�G:#u~Xr�u�;)#�z�#�*�l��IV��_���!��+ԗ}ɴ]�~1G���ց�.x���y�!��"�w�w$���� �h��t-�H*�Z&}��:�P�YI=�C��T��_�TH�?1�Œ'���dJ�S�qO��8 JF���(��N��C�����θOm����2������Y�vJ��l$�j�X϶��7Q,a��������=�#�|��;�]G�h��Tŏ:��fb������B�.yF��x�=r��jpKn�yQ%#��'��f�����O�-��TS;OD$�}�{n����8(���|�š�P��cU�F��Qg�ܴ�&��u1�'�"*\gp	�X?����Qb?HC�M���!�3�;� ��������k�١�<̓z���#l ���f���y�����IQ���I)Ĕѓ��:�6v��6����x�i�V���ػ�`�O��/�p�����t}逶SS���U"�Uz�waf�9�Õ�Rnlߩ�h�$�Th�����R*e��Rr	r�ȋ��Ӎs	��Wi%{�RL��_��#o=Z����5w��ƦgL� [�
�{�J�����4�;Z��6�����<�Tyly�؍�.̤;�Û�w��
�J:X���p�> }�*n�6&x�~&e|}��`�<��&��o�l�Hn<�GE���+[䫹�am�^ћ�hٷ�M�C�}������	͗��M��F�W䃗���K�(j+��������x����Q0�H���|/7c���k����0���V���Pd�0��\��?�KA��6v�)���B����h�X*��_1#p�=P~0D7�m����OHW��&���J�@&��D<U��]m�-I�5o�(F,��r��̔������Lد��CRu� M������_�#6��ُ�]v�I��C��XV�g�����Y��*�T�r�0�����k���;���dtvhR{iB�ۺ:�r���ؚ�y�W)^�xK�;�0�Tʩ�QN�1�2���E1��*|Y�gn��U��PΎ���(�ڴ�����z� c�� J���k������O��������'�MǿtU�?%B��T�S�c�<l)X�%$�H����(ԃ���ϱg���U`��Ed9߻���=8Ჾ^}���^��KF��ۗ�q�Wy0<vej �x��6���3Q�mV'�zFvgZ�c�J�ǫd3g,�e?����!�_�vU$�o�|��lSSLB�v"�D�"!�P���G�&���E@�Xϴ��RN)����C��+cZj����`��8�	���r���	�,�ݵ����`5p��X)8��!E�HIod���`�9�v�@��]1���srGg�`��~�U��E�OX��N�HZ�ܪV���6���{d��:*Hլ��A�d�o���oh`��Rk���K�<q�5����)�!i���T9�b7������Nt��h�7��V�5�g��f7���/qpr���Db��롇N5#U�JLX'�_��(�-3◲�w��f�Ϸo�p)d޽/G�1$[q>�arBk'D��mQ��.�S���R5A����Z�|��r*+�Nٜ�lMϵ��eo8o��AQi(�l�t��:W1�P����"�d��0_�&��֒�_�V��Π��%]��;��@��/�_�WɎ��.��Z?�"����|g�2�Ι.
��c
��G|��I�-Eљ�7j�
�Yp�7h�%��J�Ú'�6C�y|ᔣџ�M9=��u��1Nu�����4z6�|��yԫ�=���{����78����/�q�ɱ�U��煉4��_��:i��E�{.�i�
�C���EHE�1��F�V �f�w��&I1o����4�E��I�@Ɍs�FqZk�E��R���F��1��e|^�<:�I�;�50��0jU�� �j�C�����-��Ix�p�PAuC��ZG�=�T�VGJ<���$�Z�RC��5T��Un�Q��ʭF�RY�Cn��[���I��gD0���f�F��^0�3@�DF ;�� �F�r���F�'!8���fO8"�eO�Xu�7�Rs-=�6�%W{�ûL5vY��K�x,VuȺ���o��D���8�d6�1h���]��Cf�V��{M��o�S\�������n�,�Ͷe���y�u����󽀽m�<(,b���z�=#�)R��c���:(�*8.���!gf�-� �G��A�rƬ�	��������K�e���蔟#��_�������y�y�O��2Y0�J��Eps����Y�`}�ny���z�P��<��WL��A�
�@��M��q�BL�J+"2ń�5��8��F��($�p�M§��~�\w%�`���X�xz��O��%^ǩ'O��nԕ�U�6x�t�3�̴���A���>S����_M҂)��RܓC೼	���So,ۏڑ0\M�⿸<�T���� �N l���@�M�]��K˺v��E1V��~1oZ��w��/�Y;T�S5���9ZD��H���~�FWѤ���Z��>�?�ńܗ��JS���=�����-{��K�UB֭�	w�4��`ђ ���S_F禃��>�l��{D����{Q��_+*=�@�i��0 ��U�-{�[r0��X�,Z��g��\Kw9@����r9����7Q�=d����>kW�X:y��Ȗf;2=�GF�5�%,>a8��g�О~�����4C��فo��H ]5�P- ZM�Mt-�^�SX�+&�ԣ	+D�Qm���w|�UzAq �.ff�[YE4�h&�GŢqh�G�@��0>��X�
m��B�1�FR]�t�X穵)��������BvweOUr[�z��B�9����u�4Q���k��~Ķ����̍i3�h�!v] ��M�'J������m4C�����4T�7��I&���'��}�`R\�ۤX�!L���F[b��\'Rrr�}n<�¿��� ��&I�P��օ��h�øN�&]�����H�{�����`Z������=��h���{����+?����|��t���dn�nU 
_a� �I���0L����x��Qլ�Z@�(�	��׶m;��"��_M_;%h��۪�y*��f��L�PYlNc��4��ǩR{�t[(e�@�&zY�؛}���?�IE8����w�.���>�R/��"�xm���l
_�nVwW�_�fB��%�bK.�⁕�A}�����⻑:\���\�	ؾVc�M�j�	�OX�r5�CɦV��F
�-�Ď&�-��L�2�(�Ź�&Fg��0�wD�a���l��v��i*����N����p�{� �������Ioq!6q�9̟��	r*'�iAm� 3�3p�j �^�+�qe��q���X��B$?4���x�*ݨ��C{�<�����X��~�O�c�և']8�-�I�����Dz�iB(���f���ċp��]�~�"ۆvI<0
��)<�Kp`a��}}z�k��Q�|�\t���=��s�°k&�MB��&Y�=uT�׭m��+;zm�m�
�;�,p����ϧ����Z݂u����TZ�gT�>��cꑢ6�: �g�1�4ޅ��
HMF���)j5Wf5*��c�5��3f��C#�g;�%��#M�2�[+�+�BU�k�+9�	��=�V�ՐTJF��ƕ4�mGIc�AՊ�a�[R:m/��Q� ��i	ǫ^�둖W�)E(#G��9zC%Q�2 ��M���:���v` <�F��>�\1t�)��e�Mt��쐑M�:�aq�Z�T2xCkU����>>�2��^{���_0�j���}�(��RT\_n2�D���e��|��8�9ƟKو�qw�I�q��{�����z&�{���|mGia��x�wԩ\IF�%}����l�����u`5�HaX7�*�Ia�퟾�������$f�=��w�S�gBK}��3/�4����w�8�l���T�`Y���q��o���c���HW���8�(ϒ��JP+�daw\{�{R�f����9�Y��y��TT����U�aT���U
�B��x�����X|Ϗ�|R�{m�4��|ſ�u!8Z%y61�l+1T8 -�D�����44K�վ"~ŸA��'o�DtY�Ą۝&W���i����:hS߫,b|(^���zV���g٦�O���g�.wM�����
P��l�.h��F3�f��\°��	��*�5��1rG怬�P�E����eiT���ě~f�-�~�}��F����gĂ����K�� ���)�9n�&�5T��ȏz<B���	���4ڞw|�}3�s֬+&��;3�K�G)�A	�[u}?0�+��?��I7b��^eJ+�K�?V"��9ɪ��I`i�_𻝞�糇��׬�΃��0N�R4�45�}����2b���C��������pFϟ�0��A&0�F%M�,��{�4b��nK��kJ������}�o��9��\�y�q�E�H8ƛ5]XC�2�<�)#[��{�s����>��C�m��d��z*����"~
�����?ïUAr�̶́4d���r �w�Ғ9[��� 6�6�'�?�	��rPP�;�F�(v\�~����m�D�E�}�N��a�r�pmlwߔ5��YV��sP������7�峈��f�v|a+�)X�5:{Q�Ձq�S�O1�%�N�eh_�\7�g�Bf�i��֕6dv�Q��rE�]�8�s!�5���@V��Kyg"�,�>+�5�QR5GҖ����j��p`;�,|7�3���B�K�W#��W���(�홤B�[J�(5�R�깠�399��h��L-�>���� ��ֺ�
�e�ë��K�~��s$�)(�o��v|�Eu&#D"ɽwp��p�@��$< {V{�1�~�ݔ���5<F��	��ꏀ��ᬔ@�~�՝> 9 �E;S}���!c{�Gr���ش��[E?�$(6=(/� "&Bz��^�h�g���NP/��0�a�-DsxO�����c*>6�"�D�&��щ��P%����L׈^�)�|��:<���nC�!�eSפ�ׅ����r�Am�_������oP��s�$	ue.�K����?��%���Li[�N���6ޙ� 3?h
[ ��Rn�_�C#�|��2E�s=�3�
3;l�D�Q��]���A�~02NX~l'͒��=��U�v(E���J��s�1f��u� �g
B�|C]�X��?ꍾ�	�,K_��RN�)�*�z%�/=K��g�
��&�y��Щuf�t�X��1i�bHU�	���w��HSij&����fRuzJO+��.�A�Z"#/�S,���+Z�`+9�V.��|5?�9G�o�s��M�&��R��B�������q��l�r0������?�ӝ�e1���,�#� �o�Kq��DS]��Yr��M<~I$	z�Jz����O[Ka��� W� �u� �U8�d��f\a��pUh(����z��A���%�����#�>�o��\�X�\�J'��3�#����8�_����X\2г�l��'l�Ē��q�.���d\�%3����ϝPO��*y������`�8;�s���o��^qZ�j���W����M.��$�y砭�ڞ��~��O�.�����Q�x���|$��&i< "���}f���|����s�s�~!���~'�	K$���u���Gܹ�.������/��~�B�`թPಬљ+�b���c����N㷕��L�f8���A�2��v.��pGv\DtA�>��""�'u�a�����Cc�8'(��va�������=�@>�g;���J��,�ü|��ʖNlA��d���t�e	U%�添�lx�mK�5R�+"����K�o�u$��h��$^~|��]���Vߓ���M���Ħ4�;XSBCc]��a��?K�øw�۳7���N!ᚤQa��S���>yn;E2��>����q1���.�hITf�U����^}��Z�����!�?��v�tXBj�
A1���C	*Z�Ω�S����Z[G��W���e7���L5rH*��Rm#�g��a5�������s�F�s/a:dn��C�'qĮf���n%�-Xg���y{��R� �_��H��� 1�WFO���27�îm��ޗ:6WC��U��k�8mwu�ĩ�X%����\{�A�q<��0a����ip9�ʩ�,����n��	F8C^�gc)��{�ę;>y{�˵ ��� K) �MښA�ߤ5R�߳f�j}X2MAQ}n��p/b��/���/xuP>��mkY��T��<v%�	[E+�d!�@�Qe��;�Q�e�%O��X	�i ��2�m�%�U�)����_H@�ߊ%�zeq��0RR�M/��L��Е0��9#>����U7SZ�{w$ԧ5�}�hV\b���I�b*hM+;:Јj��8�
�&����`:5��a�#�M=�*@���٘f�pҟ�>�Z�s�r�b���u��8j��|A_����P1׵��:�����[�١g�͑6�~"z�]�Nj�l�hQ�%,���D�i�C8��0�/����K�E��?��O~\|h���'��m��"�P[��L�,�6yK�h����_ �\® ��5ޥ��%89����Oԧ^��f��e�D�o>���IGS&�Q�7E�ϲǀ,�M���E�d�L�,*(�0La�i��^ۘ���Ŵ�e�o�FB�h��F��.��e�� �ӑ�C&��8�)��fV�W��$��L蔣��o��C��~�:Čt'���l|�mGVK���6֎-w����L�#PoݣC�V%ViӼ�S��e���O�� ������ޜ�E�̣Z�{!�U�b
�):	����gժ/��m�m'֔�_4�
n`��z��d�)1��C�����t�:R��>V��ک`L�0�ڙ�$Jc��M�m��?�0���#��{Pq/���1A9��ד��U�ǹ����h)Nך��'�i�_�_��[�_w;��O>���T?�0��V�AH�d�+�yݮ��٪�bA�R
o>.p��N�Xi�]{90S4��X�a��)�5>P�U�9z�T���}��t\ƃ���f\zg��7.:�J���e~}ƣ������eZ�%^
֭�*�%�:"�n���m���jv�f�Ő=�-��E���X����jm<}g������MC�q",����h���9�-��L���ʍ9��K��?}!��$mU��a���ʎ6̑���?'|>�1+�m�W����x��Z��J�*r\�S���Y!�_R`�����K���Z>=g�!\CYg �M�2�F�<�A")_��nç��ŴdUG���0D����
!ȑ�x������ �d�;�C ����]��Q�h��FP��5�l��\�McsC>��<�E�p�N�
g�%���(hw1��7�#C�Cӝ�G�ެT{U�hh�h���,����`��e�{A]޾�$S���xNT������Sc�m�Q����H[l�Y�&:�e��M�Ni�T�J_>Y��dU�¶�ǯ���R�c�(SZ�Gm5=2e����#<E�Ym�V�!G>!Z7���p��f��L��2\0�*-K�������q@�⭊���V	���ԗ���<����y�ٵ��`�J�Z�A��OkG����e�a<���2��(YQJ�ں�lT*��R�'Ρ� �fp�q�]�� jWE~0������K��o$�0��A��& �^���
��
������",�=á�O�&{� շ��
HF�]jU��4
7�`x�fgܗ�YK�<�9��ٱ�K�R�>_��&����ف�g�Qo�4竿7X�Q������2����l�\�<$.驒�N50Ũ��غkb@�U�Ќ�U;w�Ǳ�����E&��vJ��y1=d���ߐG�UX�a>\�9Yf���"5��K���u���-���P��f�砞n����A��"�Sx�o�t�Fbvd���DH�4��|������n���Q�%SoK�����:4�cu�C����{Y<iǗ�L��̅�:�H�,^*�
��x�-.p�$���ϕ���٠���P^U�d}�H8,lb���;�aNEZߋ��74;JJ�L����U�U�*?�bW�O1���V�M�@E¿��MCUz:�V�S���5������k��S����Oq�fxm6Y;���P׿d������8I�g͈t�5XĐ\��\��њ��œ��un��V��~w�H����v�*P+��Iг��R�����ݍ�6�!�+j�rq�<q�CPƈnwC&�*ryY|	���^U�v%����~>��jB���`� R����S+m��Fb{�.{FM��/�n���2ë^��s�������0�+O��.�&Β:uЉ���_h��(!�ə�f#h�X�����)��������+r�`v>��g�v��1�<�`��p�R��g�&{��Qp�_����5?��z� ����o3bS���%�"����b>)W8�l�� �������ԙ�Q���0b����X_���ߢ�����]��B�>i&�1�SD��t:��k���\Y��| I_�0��$�c�%;,��n@?�Q�%߃���w����/A�,c͹W+q���=b;S�e�����-dɥ�(��	?E�=�gp�q�hJϬ�h�8�ںT� �*\F�{癱��RSm%"�Oەw����.��E7'�ct�f�#�|��f(���7�� ���I��f���/���b�'��T��0�ʝ�R��H���r��1�l<ށv�=�=�F��}j������@��i���t4��M��?p3�P.v�=*e�ѝ1���5��k'�O5>���	<� hX�0�8��>�\*���D#�M���d���\��.X,���<ͮ��[�\��z�!y>�.�{$`�*���/��V��6���
���b�p�ϓ�g@x���"4y��V B?��U��k@?�;��3�f5�ǜ!�W#^S��Ij��`C����0`ƞ�~l=�j.��� H��ґϔJb�۳�6|������ i>L�Ɇ����RF�}A��]i���#|<qEt�����\�%ý�W�Ҡ�~��ϡ)�F?�`U���
j���6�ǩ�e�f�[m%��'y�hi�I�L��2����7N5��9����������#�{Di�UBH������p��O�s 
J�=E��j��
�y�7mVGm|�E$��+�1�U1�ׄ�H����M>zw��3ԇ��k��v�ȞjT�I` 	�U�>/��Q=���h�~UQrjm��wN��;L�-va�������̓""P@�����9�*�^�w�����AU���Te�+�w��.���x��<�vV�X�~C 9ۡ3�`V�����H��Gbt%A�.�T��D���kQW����)�ч�)�͝�*�fqi}`��|F9�e�U���t�P��Ԟ֩� �F���1J��I���a�$?i_<�V+�P�
�Rg(�Z�h���^h�~߽��*��G�YSkvi";�f�b2�.1���}�%2�'(�)G�h�U>�)���$.��T��z<J���*�0;�H ��a����]��&��e��d��k�Cs�3&�18��-�_a�¡���0�'#��� �p�oGOX��`[Z�$*�k��k4f��2������_����^��a�����s(�/������`��Jw���o��V캆ro۫k������2�O�DI�K���&7/|�{2����#4�2���|���J����S��![49�O�KRx� )�O�P}�o$wY0�R$�{w��Y�L�q�����V����>+��Y`+oyaMƊ>�y�U�)�4��Pm�%�<�71�����H^M�	S6ŉ�-���*,����#k�	��-�~���\z�m�t(,���t�d��M�����B�b��P"��,�"*
�T$x��1|1ql9��w.15Ҭ�{wV��tn	T(��V�K���U����[�{SO���>�-N��5��l[�J��	�!;��>�P���M�D�s�t�Kt��S*�����ǀ-�N´f�UWD��W���+# �$ZBp���`�u~��Z�[thR��Z�|�^q�����ȩ4��3������#?P�X���4(l�v����),*��=�Go�c�3�z_������!��N�8i��L\��-����]�pQk�3�oS��f�k�c _5��=}XU|!�ƪ^`��Cv�ާ�̀�g<J�����(�n�0;��g��5@U�o:{W7yy>at�k�����;�;o2IS���7j`z|�0V��k9�_�A�j`?����H[0-��T5j҉
T���1�<��ڗ�ОjaڒC0���ũϊ`tx�颶�y�@Oe�Nc۰&��9����Y�w��/��S[�!PɱR	��2� +��L7��ӕԵ�-�y@�����0OR1��Ρӽ|;ՠ�>��KQ�+��;���;r'�Ps�V���arRR�aNz�4x�w2l�{�譵�FK�6��wrG�'���>�Mq�g��o�Hw�K�p��{MWxl
���Xig�*X���Q�4&���Z�X���v��z�ã�㲆Oo��2,��B��M���Q2�7�ܯ�^co��MO'O���	1�B��8�.Qjf3B�����9�-�C����դ�¹̕.�G���4�i��a���\Q��,��!W�k![�,����O���횎ߍ�6�;/��yL'qgl��rq_}__lҴ�)�U�G+ ����4ރ}R!$�}]��%����;y��)rT�[�ߣ3	i�`7-�y�젛~���4u��L�k�!"5'4t#�t�3m�����4r:��z��5�U�@{��
��&�-�-�0����9�+=�ђ�+��%��D�yK��-�P&{����u[�׭��㳏�~��!,�S _�;l�Hʵ��1<�h=�G�Iz]o�HȒ�<t���S0�V\�?o���)�K#��!b�V#�"��UV-����� /RH�������O��#'򒔞��w��� !��F���\�Y���7+ Cp��U�/MFWg�UeM�_r|ŉf��
�#Rm"�@0��4R�5�=��X�(`h�G{�U��4��σ��z$;��d@uq��H7�щ0�j�K?�m������E�s�^���W*w9����H��q�L���0���5i٥�tFb�Bn�y�ޒ��謔k��?Z6����4�zw��ic��⩃'�-�~�!���]rT@!��bn��dE���]�Ԡ��/2&<�=���&���Sh�5�*��-p K��/���["cx|[���n���%S��i���q���-�D���"�;f��O����)��s��W��=���+V^��U�4Vg]�c�N���>�kq�
��m���W;�K�ѯ�ȹH�2�,Y�_ã���1�vs��،����
$�h�u�u��`�_x���I4og�)=n
�é���z|^X���$&�ǉ��E�0�Y[����z�L���U�x�m'A�k������$1�Nj�j�z*����������~��-�e��L@	pF]Cu[��T��3Uٙ�@����[��2��I%{��ǭ`���Vti|{� >"�yky�)�����Z4)��c�6j����'�ʊ�#, ���ӌZ��	�ۺ�S������W��/�����ۡF�:���r���Ok����\�R�Լ� րn����x'0�V�WɍB]���� ;V�A*���궐OJN�g��l2� �"�|R�}�շ4wA�_T��
R�PU-���n�ߑN�9y�5�(��H�`�Е���4NcA�}"� ���=�ħ%a%�+������ �73�ߎJ
rMpങ�#;j�@K;�����r%b����N	�`a�2:�LW@6%\eҤS���]lP9=��4�J�N��`�~�Q��W8�
m�"Mw"'���#D;!M7����1���Q0C�so|���\�%�47�Y�W"��4����M\}oo���
���D+_��kt�_"��>�L�*���r���=�C�3T�J�3�z���I�9�>��7�~�4��M�T��eQ:PD�E`~K��a8h�$�u�/W�2���租O����a��e�mE'(��,��b;5O1t��O��FIa�lٓM��z�j��D�	��գ���]K�i�hKK�� ���~N$�zZ1;�Rm�PĆ��r�"T���Cw]���Ͷ.X���׍G�Ծ�	U��'뾬e��;��mI�x��7��%�X�#��F#2[�ͪ	�8�����O�0ղ���Di�1��sgg�&Ě"JK�����.'�o�2�z��e���� �׌FQ�ᬇ9PbF��Z8�6��0s n���D��0���Vd�3����L��t�C�Pk���E}��>�k��z��l8 i��Q���t���`ȷ5IF.z���aJh�i;W������m��i�h夿0Y<Fq[�h���ќ�D�_h�*�+`O���Q���i �F񡣣x�K�c�tXoڼ�Z�%J/�[�V����xK-���$X4�J�+��{'UW�W+�)��+tuae��i�jBm���~�O��hn�VP_uڬ�-�B/RK��do �Q�+��.U��kb���1K_�\3+��ɱ�U(�n$�>cv�f��ct�a}�Ծ�M�Sck*��c����?o��p�Τp�M44֊2C��cY/�RշJ���٧��ˍ��r�����lL�����|j2!��	���-�A��U,;���B�0����`zjv�%!p�j��:�t���x�����BN}���C6�	$\��1>6�X�tu�\>������wT$|.(���}]W����ܚZ&c>X��0I��a�gy��4�$pI��� ����38�_O�� aF\�k(�E����\�|/�9�?
7��\�+yP�����ݠ��E.�?6�i���f��@
�ȍ�n��%/�:�d��l���ӜHJ���	5N�H�h��Ì�vQ����E��0�D�v�#��	��x'�������^�k�I�"�� �U?@��Nw X�O�Gky��݈�)���}q����h�.�t�)�ZG"p��p��]ݍ��V����2��L���W�1g1�̪��O�K'[#3NIw�'���{���BN�5$&�<4���7ٶ�r�t�6F�ۓfR�ش�l�͊MX~� A���&"�.)ͮ���Z�ޮe�L�/?$�[;�|u^rH��"J�"�%����*-����=�½���Fp��?R>�Y&H9hm�&*�c1����#�eOL'd';��� sD��2X�\]�_�>ǛB�,��U&��X�Z�J�)�%�qpO��,J�r���G������U�'��;Z��ض��8;V^����a״��;�r��&��AU��MyTa<���i���-�	��~_V���ҜP�-���<����7m�ڶ��p���S7,�Ak9ݡ������J�=BFP��������IfY��Z�-�=����J�����;r`w������Q�L^�x1o!��(�yHk'�NN:�#�??'������Dk��I�V�	,b?�E�2�B�f�����`�M��/�I_FmMX��U�,�$�J�	�Px���)��#b���P8v>����d�@|��?d��Y	�Zs��5V�9���'/����5�8��%'g~��N��=NS��S��u��������u��7@մ� ��d�VZ~Γ&6�]�Uz{�����B����0������ȑ��Ճ��n��n
��A8a(���,ɸ���n�.�rB-���1��mmԋ���έ��8i�af�
�j!��mX^͓%��!�r������P*[Hw]tk�>����$��y��ŀX�4�N��Kf����D:{J�g�XSv�
(�
�������7:Qm��_�ʈ�#&�߳�w�~vG̓�ZW& �WN��8_��Ґ�4������M��pؕs��\��&�XFwUI����������� ܴ�u�E��2����߸
+���t�T�u�o[�^����T훋Y@x�����j������C����X#���J��h�u,SG�/m�뙃N�0n�F��  ��~8Y29EԧiI�}�ʐ5�hR2���B ?�9I(0����_g���~�[��U��sPn4N`�s�;h!��u�zX�q�]���H�=�ޝ�!��/��x�l��H��`�|Vgs!��<�H����h�����"��5`�����\��3*�|P�� V��c���{��

n3#��At<���2��^�����@����jc_��-2�O턃.R���N��"��8"vR���C��X�>�X�rՐ����<dÊ�ݠ��Tē=I��A����_z3q�YJ�s�P�Av����� �B}؆�S�� �W���^�e�*� |J9�;���Ή��_�QO�������̎Rj����Q�d;~�q���4�A2�y�S�PБ�1
݀��I���O��Y�B�v����ޖ_��U�x�-���~@�C�baNt6L�^����G�eЛ؎}�ԇ�����U��[��5�A^
�⾞-��K�vƃ@2L�z傥(��:)�R�'V��c�!��c|�G�:�Q-�r=H�y@A�r~ 72eS	e�����y|�,�j�ksV�Tk%�y����Vi��b3^.���r��W�ya� �%[A�GB革�u���q�4A�,:�owp$N'�fT@��R�P���Td�,kQa%5�NM�C5��+SPkS�	p�eMW�8�#�}���[=�U����l�V��-A�]�$5���Һ��q�\w�{T��q2	�~x�M� �l�0J�����h�[�l��tN���q�	��x�`I�'�x㣴�?3��:g��N�=�rλ���^^w��B/X�/���a�����d�7�lzc!��Jr�1���<��F�bx6��\E�/�ތ	��ޖm�ݏ�e5��FJIb�����1("�.ލ�?��Q�U1�9䲰����L�@t~Q8L�2A���e�� ���� #�?�������'��Z��k��a�@/���A������l��W��;?}"z�?�LJ�d��
����&PLj�VJ*�"�ۺ�HL"{�<D�H	�<��٢���X(�\�MX	5�I��,��� ��|�%����cI�)�Y{ p��V�E}��3IG.�X�($$#�$bx-�j��P�.!�u(z�=�F�.��(������Bjj�P�P��{���JYm[	�=j���,9�[��0sW��T��bս�Ն�/U_�Z��VQ�ɗ�pO�A�w�9����9�Q���558 �OD-~N� �X����ifӻ��U�eg�$�d�g� <V?��g��-���v~���D�ml��rݗ���N��Q���&�"Q�b�`e0���Z��T����|�<������L˽�S0���^��iA�a��7N
��j��i�WҖWM��ʯ�[o)���
ES�Y�>*�pˈ`a 
���A��/�\W��Kh�}Sy��"�z�����(��}鳆�CD��U�I���ޒ��0/���谢��{�0t�G��K��^�C�Q^�	�ma�m�џ�H�1�*�)Z���A�q�z�.95����o�i_�o���~���X�..#kn���~0�lԇyp��&�Z�Ii�2������e�HI�Q)|�dTI}�"�E?zA��SE�tQ"HZL6@$ފk�cA�۬�i���	�`M:�/��	�s����Q�oz��(nFx	�6�K�쾛Jl�+��u��O�f�'�Ή��"�T6�^���g?:j�$V7������Ǿ�L�`���m,��C�'�k�2R~�̍h��65qqN�7g����B�V��Z0�u����.��偸<��0����YH�4�I5J� ��9�M�V�jRm�]G���*�~fG��y�� 	�U�y:�i��Di3`�����{e��C̏�d?a����ӿ~���� �/��w��G_K��l p�[9�~7�3$�@��3)�9��9 �p�T�顑���Y�$OY��Z�CV�h��	�Pl���;G,>:����+;���zSt����X��g�}-ީf�;v�9�g�wFJ�w3�x�F�^��DS�Z� ��J��!�H(=�� ½�P}<_�\/&�|	�;A�\O�m�i��e��. ����@��E����~u�_A/��R���l�A��
y�@��*�Z���)�^~�[�垪���8�L�ʏ{�0�d2Xw����+5B��Ҙ��3�MÍǏ����-<Qo����^�7��3��ӓN���!/�Ώ�p.�g�ո2<9���J\�xl�S:���^!�w��H��d+�l�QQQ��)	�:zRǴ�H�E^i@��(���u��g��cVD�M�T��G��y6&Lp��h_��֪�� J���߫ICA��-��x�k͞d�O  �F������m��u6��~��oj�9�3϶f��m�`f��_Q�d.�M�)>�N筩�e*~�r&Xu��zV� �u�TǨ�<��Ҟ�je�*�>��UO/*� 5S�f�Fw�P85%dH�Ծ�<2���A9 Ų�+��.E�W�2��|!}���A��`�Sn#�<�:׮��w�`�+7/�2�V�.:�H[����+`��Y���/DR,�GJ�tG�N��G�$��u?�Ȕ�=���Nz���%�3��H�TO$9z�����e@�|nBM�O�$Wуñn<���b���<u�oX����/jݮϫ\����0�=5�ynMPK���&���~Bk��)I���e�!T��X'�Ywn19�7�'G����}���b��&��[{ƺ���9y�Ǯ/��T*._��~���*�Uջ�\�$H�T���oK����,��p��2r�#[�ċ9���8��/�8�!"@fSZ�'͵]��-^��I�=�]Qh?sDK�����	�(�!դ	��C���G�X!XH��du�L��^V��	��:�x��<���mKU��nRʽ�E,���x�c���f�NP�o\q���sd=p�Q�ҽKE�ZI�
���#�а1�{�ɺ��5ۭ�5�W�X���[s�x�*������؋Z��$����Ƕ��oO�\)�����6H�b:�������E��2���-�T�ø�Y�c�q�M`�bu�v:����G*eD�& �9�F�5�W��y��x~{�Ը�0�r������xcVf��Z���_s�3�?���(s=�z'R�S`Qgf��-�,�x.נ�UVԄ@�*�o�YKz���� Ɇ�z���Q~�Գ�o:���;~�
�+N���tK���<)�T�3��/�u1�ϵLԛl��@d�����C�0�dT�D�B��}.��5��-$ˤ-��t�2p�NU�L��|8hְ��H�i�W�x�9��K��>�����d�����O�-��V����Em(��A?dl�4��d��h2%;~Z�-4G��)a�Q�~Q���S���e�,Y��m�L��
)w� ��7��x�s��� �q��sZ瑡�!V�/6uB�Z�D����gdN�P�	 u�(�nʪC�[�
rV}6�[��b\�Cs-���9x2J?R�`�
96����q�lf�=7˟���|�lC[�2�;�@T��B.���+gymS��5"A]�,#S�7L#����w���d�}۟��XiW�A�ޝҡ
��Zm�c��m�����LJ�)��j�u�61�����|Ux�9���袿��>�F�U�IG\���R���a��*�b����f)�!�ȳ
?>vۡL��IT�3ڗ)Q�1m�6��|\�X8���p	�)&��`o9�{aωK�~��t���0}�<>�)<�����]�-��6�G���o��9�Y�6 [���\htTu�]�����d�:�J�� ���]aHY�(��60R��#�����a�+��FO��>m��l�_�Nk�{���� jbLP��zݶ~�J_/���S�0�$��$(�ck;)�1"��P��Rm!0%����C�[gB���go{a�$ڠ���Q6iP�Ďn�BU�Ao��_tP1y���T,�O|����)��̪bH}��U�({��aq�PI�4n9��޲��<�՚ �`
b���f��gw���9ƻ���
)���3�C�$A�k��
���O�W5���V�m�+��,9����n�{��s�#B�	Z$�W�p��`Y�C.zI�`��ƈ���T��l��ho�,�ԣ!�nj�j�~.*QKf��E�\���Z?���Zs��tB�Y�3K�����7�R�W�e�?|�h;��fn1<�l�t��`Ms���[^�忄�l&'�{�,	�d����C��q<��px�}q��m«Z8�ZTE^[rV�Oe���� !w~�?_�^z����@{q~Yًx=�% U���i	�����)��t(�pN�_o��4B<*����J׎"!��pz��O)s{�N�5����K�<ޒ��B�WOj�r�y���	�,�J,�uW.��(=�9�s'��R$*�U��K�H��������9�jR��5����!��!K�4K���	�����hJQ���A���
_/
 �F&��=����1s�o��7�仆���H�J��'��Ӑ�M��Y�J�x��n�[WDY�w��8ǥR��9�Mr�F�e�w�b�sX��Rl���R�
o��;ED/8�d�� aO���1=��.�Ѕ�|�� �����g�+zM�:��A#�Ol"$߯>9�n�ngE��N������h�[H��`���H䤝���8p#ڢ1R�dq)
6���}�����J"��D�ĺ@M�+4�6|�ľ�e-�$^���j��Y{�����kJ�8��(�W������%�����f<_V�x�{'Ŭl�<*�oҜ���	�R2��ʁ=�C��O�A�Wu����9z.b[D�;
�w�s�	{Gu���|���8NGU~���<b���Kŏ���hC?�4�9�dpĮ���A���W0$�:Yt#@;$�؄�ߦ걝Tiۍ���|;�h���Y ���>����C�4U�V����N����]KH��Cܡ�+|���CѨ�r�,���x{�=>mcEMY_�@���s��o��P�U�Y���-��Σ�LM�������)ۛ��-Rt�7��&ƫ�%�mrZ�3���6�vr6鷩/�x�m�q��������p~f8uq�]Ⱥ�j؊�Tvh�����`�����I�tz�i�C�x�YA͟!"_Y�)�kh�P*cW���� �q�X�tf	��ȚJ�# b��A'���~��g9)!!�5��*3�e\!��R�j�"I��4L�ڷ �Lcchgm;�v����҂��N�P{�n"�,�[-��t�X7���w������{)w��e:~�}u�@��ឺ�	� �
��o90LKDTUS�&����u6�I��m�_"W�f�iH�c5�[q��}��05�ba�����B�w�e��ƭ����\�d����a���e�=ף��S?�g;q_�A�mc0�e�k��t�8?����1�X�9*{�o���h���3��zغS�u��uz��l~� �R��N.D'U㬲�Z͆;Ry�wts�B����j�y���	G�ڞѿ��~�$��ӢWw����!�G����kq��g�.d�Q����<G�N:ĳ}�W�hG�"�R��Q~+���Ѵ�$*�#((�f��u��*�,H���AK�T�Mv�)��"g�+���&y�
e6��21�J�ç1����?OCn�{�N3���4�����Ι�ޥ�g���K���e��5��[y���E�ÚO�u����D��L]��;$�'k{�[�%�+F"��h�|?}�9�n(�r��2Q(�¿g������Bc�?nR�[[�b=�
 aN���G)��PZd� ���W'��źK�+E[��4Y�ɡ���O.⟎Ka�2o����ς����9�g��B�F< ��S{!#!EB��%K
GƖ`��-���X��������(�`�X6�I�8�9�0Ji���^N�����u��%��|v�N�����|0����9�|r��Q��M�j.Ӌ�DO^'��P��|����Ǌ7���j�h��B���Lӄ��3)8kų�yɞX�i��/H��e�J�rC[_s��u�Y_
H���� ;�z� V���NZX�ǧ������w�oRfe�$Dd�/�_�Ӛ���:�5�1��=�#B�L��	)�Јvf�2֗�{��I7��r���0q�� ��6�)�fǒ���_�qb�ۋhQQ|%�%�H�q$������tEi5ˀ;;uN�%��:��X��o��9�j}�"أo�J��n��u�H�����w:�>����(��%�39�k��N��/L��<������/�����B/lN�C�W��u�=h�iO9��%S�ځl9�vv�Ϫ � PF�3� �=�0q�\m����:`p*����,ښs��lYO/� �&۫;�����/�
n�Y\��,��D\�Gp�(��H�f��f��Em����i��y��m���n<�X�I�04?�v�KD��y/�^@���g2D�H����Wk����h_r��&c[l�*աnE�@���~��5x�bTt���-���A�f	{,H��x|=�Dp�7�,m�bD��`�z4DΘ��dB��o7x�S����q��JQYs��4��p.��O8�o/��� �ؕFn���M����]D�����,������Zz�����?[�Ai�h�M�|{$�-��u��@S^'|��	qmʮ�t���no<�/�����]��Ӂ�
��?>-��W��G�N�z��
-G��Qa��b��-�7���=X���qJ]i�<̦J��/vdq�bo�q��L�ebN0�I����bn��A�����L� �^��$��0�"8Z}c�^�q��On�	_�]׆�Ch�"x+��-'Z)���%���D�@GqB��,��U�����՝�d��8�񅯈�I����r���`��<fhI��hc�9HS>���V�a�A�K�/ ��j�4 !6�S1 a^�-���*�� A ��R�g>c�]����d��q"Q��Y,
&�r~�E_��Z%�/�"�A�D)��h�5�6M���Wy+b.j��!!�
���E�Зe.:L"OH��|W;��&����;-z���zLty	��C����*��vْ�`���;C,F�M�ۚ|S�9!���%��^�7��a��y�t�\x���%���!�k��,���)j�k.@]��p*]�n��6�O�Ɓ���Z��b
�
e�>qBvT��/�&���䂂ob���}E�f�¥�)�`�"��j�5婈~"�v�%
���Z��l.k�#�]�T
p}Z������X�T���!��	8�z�iW4�P�����7<�O4�Z�l[�#��Rb"�^we3�����r�@����OI~����ȴ����4D�ː�,�R���$�� ��W�Tm�ŰT��Qi��%�N&)��9um������?�]��	b4>�@a���BI�ҠR$���$����}�Ϙ`���V�t�r��m9�Q�d�E�\f�	E�WP�n}E�����^A,�^7o�ekS�&��c�N�K@[拻]�֟,��� ^��P��{�֭���������@Wďկ���<o�k3��PM=��%v0���Z��׈ ��V���7 �9���Q����+7i���t3�'W!!�-zIm�~ዏ�
,I�(lB&������h뙪"��N�闊����0i�_�\c��x�1Ŕ�&f�ʌ��D����mۍK�%�^��4�)���u��Q�T��T�X��U�8fy�����D���`-
�q����BLbW���A���0��@�� �!��:S�G�[2��~2��l��^�X����?7�j-�P�1����L��&]�ם�t~M\���pF�b%Y�ĸ,*���sGvY��ɳl4�o�we�}7��'�#Lm�7 �eلjb��Fm;AјlB������F�blZ�-�u|Ajz4��fC�]{A�����J�;,��#2��3�5�j�J��zVL`�?x��\"��As���/�V��'�|�.J� 6| �� jd"q��a�}�d�m�l�����2��v޸�p�:���8���bK�=h���Sq����8Y�&��=��z���7f����|q�t�/�v���<�Y�,v����q~��%ҳɬ�K�[M.��AZ�1�`�R�����9����>B3�8�`����s̟4ȫ���V(,5�w�G�m��H撥�˲��#�ݖ|D���f�)���w���]��R0��%
J([U͌�v�����e���}����U�����O��0�!i!�6v�����?v� rL�n�r��Q�\����G�5��[	��I����X$[ M�Jf�Q׳���D��F^v6�7�N�V}�$��KM&���`�I{W]r�IUA�ִ�ӑT�7l�XCwb����H苫QX��j�1nBN�k�.e�	���ϱ���	,gq9��b��jd�Sj�i T�,���c�I�\'7�4��̒���`����Уm)I�g���i6�1S9���O�X�e�V���:����2���\��;S�������y��2hy�?9��-h��d���⥅�uG��Ź���4��6Xz��4jP���f���B�F���yE��N[��G}^up�9U��I�I��3��t ��R$�SN"����&�� 3}#�s!�%�rm+Vs����4��w��܃�`��5�#�^�!(t(,�(�U�)b�cz�gD�����Y��fνz@��?&�/���*�<?s�;(ڐk9��H`rI;y�tn{e7�F�<� �@�^+��zV�V�̆�i�Է�dd d7t�9�l�� Ģ`^���l�]�i��T]����D��t�F����$��2m�k��i�X�rdA:�L�;si$.�17�f��O���^b�@���Li�`��V�� �9(�	¹nXB0�Q��Wթ;��P���@��1]�
���ڭ`B"��5���xT<�7�v�2J��Rm��|uYCV� Ч���;O�0��;4�E�l�J��]aX�������ԑ�1���S^~��>�LX�N�rF����u������#ә�|�sWOXH<I��I�1�ؑ����n;�9����j��V;��(�����@�u�7�.^�f,%�(��,.������OB��3<[�ybdh' ~Yؐ�4��HO�em����a"ct�(�+�y�S��Tղ�^!*m��࿣�1�-�pn�7-v�|�N�s��p$���Ba{�k�����rQ���r!�c������}ơ��M��˳"�c�6�AMϝ���?�}3;(2җI#䔄�mRRw|�He��M�2{ccd�I�4�m��x��U*5f�äe� ����x+U�j�_�g��ވ�o:����>��[��f#գh�m��p���y����C��-�����Þ*9C���kјz���!4v��D���ZTR�����V�w1��\��B��F�I�]���)��0F}f(Zp��T�GDNS���{6e�Z:DHG��@{X�h�1�Rf.��(*�_8%% �-V��j��8&��Y1���Y~�<:��-�V�ͻ=Dc���^��f�CFO��@�#8Y�P� n3�a*�����,��ę��f��ҫ~'t��	��������G8��ɝc�����}�
5����4l?�t'�c�b��YC�'9�,Y�7��6��t^F���"�����JH͊�7��X�G��|����K�g��C� ��F2^�ny�at����U߿���Э����s�|�j=Y۰�ܿ�H+��lӐ���[˩ó}c�%abg�Mb�,��K
�^ƦN*TI\���E�0vg,M�h����T+Y�ۚq1�h3l=@n�䠦 �B:/ZH��?1�1�����_G~IxEr��5�!jz&w�DRʉ��G�����f���8F��"����*F��Щ��l�q�/i}S7�rr���ť�[IE(��J�N�I��hb��ul��F"W4f惈z����G�|�^�+�(�A�m+�Ƭ�Srl��C�T����J~��v��+�V�Lv�ݘ�	~�E���\ I�{7ڒ=jk�o��5��2�G�����g���i]�?�"k<.zn��k���1��j�ֿ����%~x�����ZS���'tG@� X#f^������^M��q��=���2��-P��d�Ox��W��:�[���-�{�ת-�=^Y=�-�Ⱥce=��Ue��(�LE��M���%2�!䷅ي]�h�fP��_�����)	kg�G?��NQQJD��4H�SM�E���l��N�.]-��R� �A��,���4']��W�w��K��n�%*��>��U"VV��K|�E�UD��:uV�%�fnSd����>L��1��u�CX�����Ժ�H���x^LD�
�;8��T��u�ŃM�P�_m���P|��Uqҍ#>uk]���?u)���/�۵�Ε����QE����(��~�$<숷̔���KV����ڌ�b��/�r�#Nq�����ҝ��yV��"kt����^�e�Q��R�%RS�=H3��#t��ԕD����p���ݳ�1�8�DĿh���"36~M:���U�ĉC��q�Y��}���v~���G�-NK�����LM�&�G����M�2��%��ʺ�6N��2�[T,5��-�0������k���lǂ�>�邽+�D��4c�پ�t>��&��?{��\4D����Yģ�d2�o�0?_�?��F�I�0�W��C����93���w$";�Q������h�3��}��3|����$Vo�����b>;�_y�ج[�}ׄ�3/�{�z8r!"��z{u��\t3&�T��_[Kr!�u�.|��ڔ#��Y�/�fr�s�Q,^Q;�{=����SbF��w3eR���O�V� �v;�����-��t~{��"qZ��o������㶕�o�~�S.�d&(�m~ [l�XO@-�3{�=��ޔ���E�f�m�\'��� x��Q�Po��58h��
����Ņ_m�GU�V�lՙR���v��g�5R�[��qd�?��=V�q��j�^���L���1�@_�ݢ�Nb�W�v`��uqv��ض�ܟ,����$ c�!}kY���k�A�P^�{��
{�t��y��r�t�6{��YV�(
}��8i|ܖ�lP��|h�+�����35�z�:��z����-�DN�l~�J�17T`f��j$�B�5>H�8��_k�6&�5x��qDn�6�>3��?����O'�j�jۀ�H����y���Jp@5$ڼخи��H'3[��͈&@�@%]"�|����l�	A<�=
�̜���
L�-�ޫ�zMt�Ė�e�i(�-@t���lYI<3�go *�:��.�1� �� 9u�b����+�#숓!�O�yv�CIE�!\�/����` ��^�~����q����?��'����Z	nb�ib����[�c������D�Kq֮�M��)r|��|�S6�q��>0��÷��NN8��v	oQ):s�u�9��Ǯ�}Hv��>�!�	��;��3� �^4�eN���V&�D����V���%d�4�;�%�
�<�\�y������Vgu�W���$�<˺�}/��݌���xiq���!��L����w8�~��Eن>!Ǽ�!����H(�� �xm�����-���1�>�b}�z�0	��B㇣y��
{?ׁc�ѩ�;�!{Ia�&��Y
��4 �:Z�4Z�\ X-��ZA���Y���3
η����o�\��P���䴀{�I'��Fr��D�:ݸU�i���������x����ឝmTA�ed���=\����R�;s�6LeL+q3�p��^�[E �޵(��ٿ�Zx:��VѤ��t�����y���O���,7j�݌+c���v��{�����)if�V՚�ҼL����k($	w��58�l`�yp��R!��K���[i�B�w^ͫ(�#̗O���a���~`� ,#O$����u�.���u��[6#�e�V�]�	_Hː���~��FgL�o�&�����v�v�2�+�5\[�ŷ.� ��$�.�Y*@�|RT�e;.p8 ���ʗ�t�NYRyg$|�fz}��CN7z�V�5�����}�{�5���yc���93j�w:�Z0m��A��|�c����b�/�۹��	�����Js��a����=��^��i[�x�C�1�ϗ(iSK&6a!2�q
��S�V
h��h���9���C�F�2��cH��B��4���`�s1��o��$m!�ٷB,�z����H-�!�Iߊ��q�&���+�o�;I��@{���=�CbLZc������w��e�W6MѨˏ!���$ϓ��>C��u>ڠ��n���5�rg19��16�P��\����A�k(��څ/��"�a���d��B����w,f�Z��+��1R�w:D��n����S���߄�h�6ʏ+>��&{`l.3����fp��k`X�S�["èQ0MIp��A0�8W��䑒r������$1���A�˳_݇���z���K�
O
M��@� M�@��xKK��y�Wƕz�`�g�[-���4�|��Af�]�YT�����ke̫�D�L̶���S�ˇJ�PU�::�Q�
G��$J���,9����|�zH�VEٶ?)��h��Kis�'+����14�2�eҹ�R^��K�w	ῆoec�����Y�sQ|RR~�˻�vkJ��r���c�k��L8�Z�z�p�yXE���`��i�7N����5hfi���m(Rdy�ZĦ�7,���w�E�����*����	�x苳�_��´�{Ptʢ7�]lYy��g���d��rV��DE�� ���?������ z	b���l�bx<�k��ތ��TB�MQ�m�d/��`8�*�ԙV��Am��/��`��B^�7Kt84�(U���ۍ��w�Ĺ���X[��P,k;PY����j˥������T���i�5��ue�V>�&�$&���D�k_:�>�/�~�4%��49�v�k��/�9S��K��UQ&����_��U��@�M��B�m�7�4��;�~��J�l��b�\*I#�����nS�Ff�˰�b3�y���N�LBhg��Œ��x7��>� o�ʤ48yń�DC�l�d4|�	L+)o�.��#&�`G2�� �����h/J��LK�^�i,�w�S6�d����N��P�Z['l�^>�������ʣ�GK���$���,&�����f�s2v����v?��d`�i�������Z���]�Lv�;����T�"#3�`ǫQ��wp;�v���$��������/��"J���V�_�Yȅ�I�Ć�k,ό.���oZu~]n�*�-�ck�޸� ���#J�M��Ts�����LM�*:�6(v�-�Gժ��M�D�L� Y���X sԦ�,�6��"Oes�N�c\/O
"�N�`�z�D@-w�}�Ï�4j�ϫ�,ӂ�V˦�솟��'�����Z�m�� �|;�J�l������t���c<��eP^(�"�*a��-�Ķ�]�t��RD�NxB�ޅ,�OP��@	�YC�	-D����G;+|r�)�<:c����'�
s�P͡sw�"�z/�/}'���)8�FG��1�F���Bю�J~� ����G��և��W�K,��~��!�{�E�V�(o�%?��AA!�¼3I�Ž�L��k�cG�
ώ�{g�Keny0o��?Y��M�
I�2��t�@N[\��H(4�_'��=���`�=M�	��c����7R�U~n�{w��}�d|��B�_+�\`�Z����",��2;o�Z��+)�OZU���J���7c�J��Ыk����ʴ{���1�T~��5뉠����,Z0
:@]t���ϩ� �����iQv�6�A,����Mvmr��9�/M�O��>���<�E��P��q�x�T �W�H�둃 �^��Q�>���UW�g-�]�¸<g�6�x�C���Q����o��I�X�&_�l�A�e@8��5��u�Y$��d��W��r��3vb]4�z�ml�^*�f� �v�8�α���mfjp�p�,�r�b�raPf�\�b�������;/k��?-�@�O��iyh./g{U�&�-I8Ɛ5)��!vȿC�ԑ�
S<�����d��w�U����`^`��x��}`/H��*G"�;�&:�&qi��<0�~��-��U��Ёً�O�W��1(f��6a�Y�UX�cR=L"!^�$$\%ױNO�9���S�-�����.��@�f�j��g�p��/6w|��Ҍ���|!^�&��������-��)��ߌ��s�b��'m��g�0P�-::��_�c_�E<��͘$B�k"6�dW,��&�.��]\eyR�u;�����?.�hP��n3O��XV����;f��}��� e�T�.s�dɚ�LM��U�1�����U�ޡhQ���<i%th%���*��^`�kT����g ���$Й
v�Herv�q ���rU�g���0�����	���C��y�'�{�Z� L��P��,��
���� (ŧ5,���A�6A5��?tgN�W���:3�JY��/��2h�v�>J��r��\߇�|vD5�s+�v�}�*������[�"��C7�9�1�_��Ή\U����>����A`�o=���� h��u����s�nL�M�/�P%���&9�٧�3v�����-[p����l���$�9ْ���(i,H.�"�:�Ӊ���kK�O��x�a5'�@|������5E��
e���_T�3�~e���^��i����>Pt�3�/�?j��_�ꜟ�D(�y qDE�d���ux�)�� *Jŗ���d�^5a���{���m�K� .�h]�笢�@s�H�m�{�O�l�C��.����D���!��5������"�S��̾�Š_`��\a�à�!���F�z8���۹�>�`�Z��)�����b��F��n����g{��sE��Ɇ/�h��/<2n{�		̓���H�Si�GY���ns���]Y0!��Q�X[�х1�<��
{ّ��y&N���$b�Q�Z�w���8@�P�+��nI|��L�`4ܦ*fV���w�ӹ{㿼�N�Bw�D�!O|_�D�rȭOY_�z�"�r�\|�����]��tI��b4q�X5���I���"X��\"�y:���>!>w�k=�!�ŞG �W�H�=#]���z	� �u����S�L������S����B�����'>��_��P!/G��D��
��jLU�/2��������~�_��/W%�Fc�$0��t7�v����6�p�����>��$���#=��p3.&�t����&�^*�hx������b!x��0r�h����	\�5Xg6s�%Gh�W����#�K�!��p�31�1-�NM!9�L�[���m�_R�p�<ӕ�:��g�2B��
�V����XIP��� p��*�_�B�P���E�E����CzR�<����=���Y�q1��
|���xU��
���ȣFC��Z� `Ӷ��/����׫�I���6�0���w�6�讠�T��c��y��#0�o�"�ʢ���^)v�ڜ���a�;\k��8�T)Q��'�����'�%�����9$�㼺核����H�S�-�����V�a�|�D1��O��3��\*d�ò'2$�g�U�j�&�S�w-�����7twNm�N�����Hw�0��` z�z��t�}Cm��Ƒ	�,�ɔ�6�B�w��(��n�o����<�@�З�K���x�&�����I�V��t&y�Ĳ�Qa����\5�{�c�a���u�<��Q��cF�]�?~#����f�������#{c��n� �l������7kj����bc������*Z�=�k��~ݠ3W*.6�&l�>���4����GH�9�����!��%���c+�ʃ_Z�u���o���
;k*��������9�busȘ��'V�����N�b�~��܇ݢ�����H�l���z���m�*���;Y���y��h��;@tU��0�]��6�6��,>�z;��s��p�u�H�/�s�ɛ3��u��/u%')�ƝP�^hILʇ0ʟ������8�����%���6 �vv9:TP�Ѱb�>]�
*��Xk�GuD+�͓A��r#B�-%0�b���	�}Rh�r�v�^�[�1�<�pm�iӟ����&'z$���]%����s�>������2�P+�d�E��[�-�3����ZYq��f�M(��u_0���ۮ��*zʆ/xq��Z�ɪGH����4����ҙQ�N|�2}#����b��z����Q�zE�ify1!���M�	m�a���Ѕ_(l�R��C4�ߟwrѭ�J����.Ȃ3����L��b7$��Ʈ���%+y���e���� �x0@��۝ �=,M���-˨[�v�i�U9��.|�����|T����U��'�V2'�k)�!0���G��y���o�wܰ�Òa�&��k+�YI�5-���#�1`��<�^0^��e�G��lƁl��%��ZzöZn�Dć�LT�M���1�+qC��i�7�HZ�e�7�Y("�VE��8u�g�yzL��u��̗D�4f�P۩�qC�b�m��v�	>�#Ax�$)?32�>�?�+E�՗f/� �������6���|Q}u��V��u���c�z/��م�l�;�6�U�nsi0U�/)C]�|���P`���+&?mLY��*&&G��)z��`��SS?�>z���X����[��F�����E�U���#mG�}5�{[�����u)P#S�#r?XB���
�8 i�;��/�������� 2��܌���l��nZ��H�v�����⬢Uc�x�
�i�e:5�p;��+s��9�Y�:�+Q
��	^K�c���:A9��޿哴�
�[�ٺ3ά7{� .A����@�@B��_��v0�iwwa�\Vd`y+o��%�~�"�4�����l���#In�[��j�ށOs<�N��ybZ��[�41s�ؠ�u���H~���c�{�ICܛ�Pz�)����$m�܂��g�m8�S!R9��P����MU�D��/�X���֒�1�.[�Y+V���@>2�=�1#2�O�SNGh�������3Gd�&�m��$�Fۢ�m����,��n�(z�D�_�
�8��x��8G)����o4�,6o� F�bK�R���3�*yw���;v�"��5�Z~?�':��%��NJץ�=�u�n.,���̡��#L9 ����. j���"���*=���EM��A��F�i�������3�f~�Ũ�_)�Եi��m��F���SR�ُ7|RH��vh�K�kh՝t�ً�0�M{x��0�ǘxzG}�b��C��,���\>���[�&�z�xژF�ԂF���6���<G8�ȸF�8Dbʺ���߼�:xK����_�y�Ej8�2Yd���K���g��	v=�Z�b���9���n� �%���RI^D@���t����2���6���<�T�WX��\�X��Z9_矑 ���F?�m�	��7��-
ڄw�_�1Xh�S33L���A>��<����K4��W�� -3� ų[+a-N�ғz\�i�k1��4�Ნ��t�:]�0�ԑ����.���:�(kZu�U%���G��H����E���p�)d�jsܴGG��l�����mʚ�Bh��}�ò���|d��b�&A��[ref��(O]�f�� �{��-�	ŏ<�l��rl���T�����v�k��[����]V<l��[g���c�~q��`�Ԑ�O[�a�<�]#����Cj�a|���ͪKZ.��nM@��nؓN0YK��;C4Ss{����}qü*�vbA5��[��`���⧱W+�iy�ó�5-k��6���)���k��==�2��1#!��ىA����h	�F���Π�cHb�4rn������q!�Wlb�"qr4�W����U͚�b��T�.)2�~jY��g��a���{��%�I��7��.	�h^�\Ӽꃑlý7U���6a7D�26�,���7�b��vk���wgev�T+�n��H]���!����^�y.;8*CcJ(��PJ�(����a]�����<
E/I��E��5帖t�$���2Q�i��-C&�b�T��j(����®@�I߽n%P*KK�m��9���Mu��!v����>�cÈ!Q�p�cM��|!ύq��{Vȕ�s�Nc��<��&N�k���ɟj�dl;%�̴}t��c�� `�>�F��9���s7�9�&�)��)�+b�*ԡ�F^ �,1��[�}-J&��|�-8�v�,$`�%����RΊ���z�%�3io}�pP�$��X���U?)�@"��0'��C�S=Ӥ���k�${d��c��������K]�0���4�I���R�����j���b�3�->^g�.�����#�-l[Y��ﲘ#rj�ʧb5r �5ѝm��h�g�R3}:�ٰ�k�7jC��џ���֓�J�8�j�0,��X�p�u�o^�]e��ߦ����)$�a���sG/P�"
����ܸ� ���aW�.�VҰ�o������º���p��p��>]��o+�ѱ2��?k�$�MO������zX5�:K䀱���Xy,/�8�e���dd��<�/�X�u����S��*��eK+�|�oy�b]���@ݪݮ�u��T���QK'�w�n�=vW>�u�
���B�u�3�T��[��ή�x ���N˥	�#�]��,���9�q�Y����8�O�><^��0�#A��9?4j�s4#��mJ<�6}1�:�U����:h#v������)I1�4\�F��6��d9��V¢��א)���{���	1mF�nX��o�P��ͫ��B�lU}���(t��g�mPn&=a�[�l��#C���D'*I��L�}�˃=54�^���t���q@�\ZkA���&�n4���0�L��2P_�~���t����UY�ۥad@��t�+�����Zc��^u�s�<�U�@TVJ%�0�4��/¿�����Ɂ�r!��k�@V�ϲ���d̮dß��Yq�M��UCn��N`�5�nok�
���ɶ]��ӝ�(�C���&�T�Kl�YM+��c�Dq%S@� �,�?[��l F����:��B���n���)�#ϕED�������\N2��C���Y���v��"�_�
�E$K�h�^�εa�Z�W�A�}Ty3���|��&Uv��q*(R�h1xly�q	�.c)\�0��?^�M�ܒ㎌ރ\n�&�V6_K�t�w��m~�Å���Y��a�
���e79<��~�2>�P���ס �=�B���-�,�+�����U� >���:M�h�i4\DdK��Y�s�p�lwP��|oey��q/{m}�����vaP���x$���R�U��͹�`�C�1�8�����ٖ���G�M��[���"Jd��y��V_y۲�ZS������b�z�K���'�4���J���k�'��#�9��\ZG{i@&��/ ������T���&(��R`|iL�[�����ٸ��EK���j�n��ج�G�-c���=�?��qLCbc�l{;��������pڷôaZ�Y�/'���2�D��j�&b��I=&ٯw��(�r�^k>`mD#)$���;�1J'u�wK��Q���S��Ur���_���¤������8��"Y���\� �N���Vuc4@�]�٭X�uhP_.!����0C��Q�x��ͺ1z��R�!�(��i·{�j�^��ޘ���&����z�H���c@�,���:x~ǭ��|�$k��Є��:oƱvI*Ld�x��)<��T�k��rͅl�mT�Y����}Ps�ܺ��H�H�@������ue�m���"HqC6�.��]����4���
�˪�`����x���I����s)���*2M�y��{�>�W*V.?ز�<�?чK	�����)'�a��dᥞ\,-)4l9��X(B�M��
�f���~�i�T*4.�xA�)���M𻕬�=�����cQ�6à<'Ɛ���e���f鰉��pT�Ɍ,��K��gbqcl��Q$k��ˈ��4�Պ�S�d�}{�f��j���A�y 51�Q\b2�D\��a�z~��vc	7���ᜬX��-Wzt���Sd3L�^5�x Ι�%���Y��'��|.k΍�g�'JU��70P���4Ivu�o�J���N��
ʓ�]s{>k�M�1ٍ�]��na��C�����=��g��k�22{��V��}61�W�Gm��]��� ˁ��~��38	J�H���)���λy^����J�&b�Q!?�Ew �:g�ͥ3��v�}�\�e��e�ή��,�&�wӈ���F.y�������t��+��5eYCc���(Q�R~�1���3��m �����$+C��/n�_����f�C��׏J���A����>RU����;(�l����G�a�;�
8*���ۭ
�!sM�����Wq�$%�*c/�/�b�(]九I�|Ҽ����.���96��V�Yr�1�;���"�B6M����QL������1Y�D���;lx���UB��L�EzX���&:
;����S�ғ�	��kWm��K-"�l^:�>�=���^�%�K�l��w��78D�_{�Pv[l������y��8�N<[��`a��N�XU�1�BA��K��M����˂tE�<��Ų����\���!����;��]W{��XS�%��,�\�� �=E�] <m���8��RYP��.����"���fב�Њ�^���A�L������m��b���Md��SY���'�C����@�̕�'#kfC`�����^&D��ʢ)І��4&쇗��vj����'j�7�6��/<F�l�����c(���S.��Pb�N;t��#�7�,�-\d�g��lܳ�T̧�Ҭ��}��<�/���x�A_3��? o�ݲ��u�$U�A]C���~�x(�A�I�Y��#>Dy]=����z�1IK�g|m3�࢐I1H��v����e�"�%d���/>�'6� r�|8'�L�8<;��.�r˶
v��V9�h�f������
�-Z�����.��e욧~R��^���:3����p��(9��rC�?��֡ ��Z]�a��5$�{���*H�G'�@)� ����T�����)�M-�C���sY_BҲ�+��ѥc��9�q�ji]�hDj
8��i��z=O��4��ɪ!l�̅��\���㏢Ux���ȯ6o��	�/_7��dV:�?��Z�Ǖ��;>��ߣ l�-�4a��S����#�J#0.�'%�DptN�@z5��,�b�Ƴ�����-lٞ��5�ro��H4���[e���8O�Ρ��R^�| ��!mŇ����2��y�
�����$1��.���=-�x�iՙ%ɴXo����UP�5�J�JIjԾ�@��^g����0�Z�y�*!Ei�6Q�M�"}�H#B�F	�xhl5���������y��~[�R*k9�[�P�K��xím��%8S��<���&5m���*%��&����5s
*a{?�Ρ�u�fo���p�ZP@��?�7儤�A&�7	���>n�D!�m(�>H��x���2==3�����).I�T������7��M�zD��	�^\��М׼}�v��:��S�-ŧx@#��x�ݧ��4&��ٳW}N�^b�Z'\9�~��k׀��
�iY=�Q)���P��	�Uw:�p:��Ng,#]i�A����G��3xq0{��@�*g�Ol l�h���
�5Jy�f������u��beΪ��:k���4�gJ��b�����5w�J�L�Ӵ\X|�_W�2sO���Y2�o?]��O�P�\�_�P�r�.���$΀AI���N��O�R*�0���y����,S�����b��4!1&�@�c<ٛ1q�0	��N��d"��A��-U}J4 �pp4��U��Ɛ����t<�vD������V��D:�=ŷe�G������U���wK��x��U+�y��$�*��P[���-�^6�Y2=��C��|�<�2��
h?��,e���!E�o����6,����,�O�Rej���e
fmh�A��F����FtQ�_�>ed�Fˁ��c��ad,�n��+9�Z�&�{.��-��&z}�Ț����5$�.XGr�,"5���Tz ׯk�e��!	�i{ncCu^Y��C|0�9�$KX}����Ж��E��Iwbwmq��A�Y�8l���?WDa3�o�R��s�e��g+{W�|��.��1,R���X���v�2NMsk&�4<��<ͦ�<�u�9�by?f��%?��Y�d��tBw���ـ��� h��C]d���CT=쇻j�%&?ޞ,�-Ib�lh?<���K�8t�XiK�N�x1m�u��fk\���.�0G���Y!����ミ�6&�S�BQ�ͳ�(1�Z?7
��0T���?���C)���=^��]K4��T鈰�)R� �*{2!�3�(�w9J�N�s�j�=媾?�!��#�#Ҙ$ζ�l���U+�EQ�>�yn W�U!��K��Z(�]���bTu�v�=Z"�8�b�R��w�lpE�_u�f �%_z�_ݻݟ �><����x��k[?� N����%�v�[�	����;��â��4�Ք��ї�m���T��N�25+����<�	^��E,!J���XyM��)_��`{�C/��!Z2Z�2T�8���gh9��K隽��٧��p��J;M��c��/��,Q=�x:�ch����t��Y�L��Hj�@�[Hm�:��V����˟�3�`�W��l���������!�% �6r�\�e!'�~��x�¹���8���>)o�rZ	���\�����jCӡ
�P��D�d"��p;��ĝ�߰��R��$�#Mg�	�i��;X��r��e\�͉nlG�V1�J��ϧYY "GZ� �s?�տ��*15�?hԛ��0BI�UG�?U��/U,|g\UH8�^�ܺ�$=_�D�58A�
�(�W� g�~�ת9 ����l��bl��W��*'�FZ]2��}�C{epdvu�xgd�cs�Ɯ5LP򮁿⁙����)�hU� 8�H����1f�'$�V}�3N�}�T4h���'v%���t���{,���h�F�|[t@�7:��J
�k����\��� �#bH��/p�����Ț�g�tS�U���O�5�,h�r��GP�-��R�6B�M��P'7q�!�n}L�m���sݥ&(�׉��������2��<1A����P^�#}Cga���A��=��N�����\Ԫ��ImKm&��4��������?�>�=�5�cҺm��?��Љ�e��q�씥��/�^e�s�J.�)���x�/���Y���f��}	�n���E� �Ih�$�^q���_R�|���QVY�'�?����5�Z�W��4[d[���2o˜}:'�[���2C��*���c�̲���$��,͔~���$/�q��������-�"q�TP�;���+8!�c��k."�u��t��5�:ܻlt����M�|�	�O.v#̄U��|Ռ�=k��	��'�7j���.���E�A���棎���۰�[���+����"W{<��U����I�"t>�h�Dٿ�>l�րHk(���H��w���;���e��}E��H(��6���!p��e�]X������[,&���N(�m���8��e�j���)s6�Oy�� �-2�|���1�/��ls�V0%WC.�޺ز,[&�I�&i w7�.�f�����c1���>B�-5~��EG�䏴)WU2�_1A��9kWz��cu�m��I��)��1e?4 5�Ih׹�aj�8�:Tg�V���)O��JYL��^VXg[sd�a��\>u!f9�����]���QO��l�%��|Q�>�
��%�!
SB�4qM��-���l_rFg$1�ǠE+��2�>�|K���hr>��+&��1����� ��u���2\���1�2��t�Z�OG�&�f�i��՜����MQ:����2�9h}�U���NN�;�E ���u��@ubg�T�*��[ ~�ii��v,�.aɘ���co����C�G�)=������6�U���W��bg����|;'�me�儛N}�Z0o�1$[�m����
>��x�k�U ')u|K@ww�|�?P�?T
�Xa+3mtz�!z�#��zO�cy:����oDd.j�d��.%��i<����;ak5�k٩K��78���$���H/r���ؐV 8��Z������2��D�T�!��yr!��W��2���������$y
�S�m�Ĳ��%��<�f���,�	��J1�hR��?�4�<�[����\�(ןV�ͽ�����R����$�V|�*� xg2��E����g�g���}�;��lϪZs�h��,XްZ�����������+�B�YK�3�'o��{@����]
\hl�T����G���	W�?�����`�Ӎ,l�f�q�q#���В����8l�B���لBP���8�_�FzW�h��.��!;<���mJ���iq,@[�(v��{�E����jS!]Y�ʹ�(��MR[eý���ɬ M30�l�)�
F�5�g�YHa��nEf!����ɜ�5���B�
���z��|�����G���e�ǟ@��[n�"�Z�QW����*���8����H���Ih(4!>�j��m� �i�~n<����fx~�RP?ےк���Tl N񖵨�gW���BP[)���e6sP�V�.����A>��<\��	H��e����K��"sD��g���o\5Z����A[����9X�#r��vò�F�7��8Y�H���Et?`�'j�y���-�u�FY�}
G�mP��4�X���e��*<��@a���W.�:�y��ܑ.�G#$�����)IG7�u�A��BLO<Ǎ4�	�#�E�r&�e��Z~ә��^}�<r�w{(����e�5��H�a��jm����&��}a��E�+O�.Q��^`���;��):�:i���n��Ia9�˫O`�e�g ]ԗ�E�n鮳�^���`���ؗ�mTc){�\���͎|�HK��ю�r�a3���:#M�����R$o��D� ������;y.�2�/Ȍ����Sz0F��xv�R��1y�A{{��+:4(��韏��P�U?�F�t|���w��U��M����.lVMQ�(� nR����[�]��0�g޶!n6E�\���m.Xpȅ����)��u�|d�L��g�h���P�:r.�>�$o�#8�Mz����ZzA��q�7J\�[J�,#��Қ���fRa��*d��W*.�Ÿ�a���ȉ�ù~�LFa���X�F�Ա���T6�ԙ�lzi��x�S�M�8a��[2XyW,� �]���g�X�4�Vy(rR|T��P�DyO��@�N�x��!O/6�#l/&�5hq?%��Z�_�ډ_��Q�l�2��`�u�� ]��s"$E������σ=;r���Z�}Z�A��v�>Pj�c��)-�4&�"E^�|�l��(/[�H�R�O��Q�b��=�
�cCM�\�@�\.�`6à[C/nQ1������w��
�6è��㳑@����
Ϝ�c�Xc�1��\c�D-A*�l���-i���Ҡ����r�����A(���u:v𖖽⎅k��	M����o��+���M�m$�x(��&�����A���C`.���I��Ь�8��[:E��f�b}�w��l�}�Í��%��>c�M� ���g4��x�f�uL��A��:�EZ�<��B���k�`%N��$�c�[��ub��� &�c]���֑�}�9��x�]�X���B ˺����s���ͦ�XF�W[A�ҕ��*q3w����������*�S�'C��ʻna$�Q�;[������Ŀn�U�S%���ͮ�4�콙F-|;$GVOg\����7�>��K��E?�F�H���X�_p~�\}�Qw���A�6cg�/�<��s��{� �xP��G��~���w��0
m@��R�B�^���o�(Dyy��l�ҫ�������'���'��o�Mkؕ�H�H0�V�u�����o�G]�B�g��ib�1y��i����XntA��4E��5t/���T|ot&"ӳ�O#yJ�6���0o�\��P�x��nLu�8r,�l
��phK���X��SAT�IQ��E�� 5 ��kUf|Y\�u��
Q�J��'0R��h|<� Z��| *o$iqe�H��TW���7�o&����X��p~��zߥL�H򋰖�Jϰ�&�8�"y��Ch>ȉ�iY��u\�J QH>p�cc�;TO�$�X�����1��U=OIH�:��x���2�����5�x�Q�����x�x��߼p����=��?}��~,w����V��^��?F#1�lW�<� �'�|�w�<<"�g	���?�z�p�G�L��	��b�v�R0��Hơ���漗�7g5�ᳳ!��P�S~޴���#O���s{1	�֙TC0�4�i�]������T��v�AQ'a;�¨1�\�;�Gb�9Xr�qR�Zd�e]-p��M"�@!���!�i>X�X�pT�=�8+*W&x~ޞG���q:�yZX��������r�Ȏ����M�+��F�i����is��X\����p
yM�&�ć$���Di��oh�&�3�^�x?�`mJ4̺�/�"��-��^N_(���u��q6��Mm`|t#xQ�a8ENK*�V�F1s6����o@u`#jM�d�;�2���(κH#��U�,���3�h��lʪ��}����+/"�1�Y};1>�1�)��R#P �b6?-��Ef��0��l+� \`3��f�U�Mcb���
9�YۥZT(ȓ�T���:,��Vk�HZz��s�g#���v�4l��q�	�0á�~|0�J�VJIC\*$&�pz��4��S�Z��Eu�iy�b��T����|��6-�Օ����ݬL����(�}+��a����=�.G��2�|��!Q�lF:���ڀ���A��*uQ\�[o� �eZ������6��
�3��A�)J�I�|�a�+z1R�f�!k�l�=~�(�с�s���o�e3'�,A�<��w[aR�x���z}��c$�k�d�5k}�Ђ����R٢�@�Ѷ �l�����a�|�Q% �@m1�t���f�*,�J��	��N�T~"&G����kh��j����L-7��VF<$�Б��0���L��p_w�j͇�z�
�2�P1�|�%*m�<y_,�Ɖe_�y��#x��`E��2�%�h�n�k%ї����!f0e>�9C��^�^ i��ᬐ�!Re��û��+\]�D�Z��#A��zE��R�m�R�'۝k���{������W�UO@:b���<�g�gA��0ϗ�e]-wV�ԋ�\���f��@��-+;B�*°W�K�o�ڦ�=?S�� \}�
�	E6��פ�̝�͏U΂H��`�3�-S؁�t�