��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]������]��𵗚6��W��dy��Vu�*Ş�2��aK��o�/N���j���ט����4��(���W�_����2�	Ų�T�/�]-�2�AW[ OF?���
I��Xp�$%K���@!��3�tx��{f&bh���4^;tS�x���RL�O>N+S.��<=AG�/K��{���]w>����,13E�[��E)� �6�.�.	U��ZՖ�q��xRpe:�=�*@�IK@�E���9��u��,��3~�rz���4������}����qQ���[��[; ��jL�M�
b`�)���N��Щ"���3��49�9f���m�x����ӸzH��0i�U����zd�΂�UPa���ctb�����:��cX��%���,�'�r��ux��δ��U�-����z**s��~�&�Q���D�t���M�28�7���9����FR�UH���vw"x�����GRB���tm�-ᩣ��+<�^�jw�]0��(xY���i��h��`����/������;@�D�6+��<�@��_�����B���O+����I)�''S�/O���8ȰesW����p2��|�&�t����B*�=w߸�e��R�mn���`�٢]u�R��#7K�d�/E�7,�����e�p���%"ԉ���'�k�Ɏ���A��!�/���������߲��ҡt�Q���a�]D�e�xڐ�joj�����V`I�N����)��b��x;���;�O���Ù��1gU��ӟ��F^io�]K���Y�/1����/oO��_q��Sw���E�����O��A
��D�=~@�����+�����g����U�ݰ���o���*2P�8`o9�*�s
���9�ğ�m!m�"�m���0U��I�0���g��2J���nP_s:�~��Ȳݽ؊~�_!78�� �h���տ��q��b�I>9��{j"�r+L��ٝ>m�۳'N4���]xR��	���{�i�[���YѫR%�`�,N�b�h"Z_YW%T��n\2�I�x�e2�QB���C[8�m���q­��|\!�,�>L��*[i4T05hj�E��S�&
.��y-RT�;�����L�g����"���F�3���~��*R?޿K��< ��m9��CT����c�/����7���2x۷k$έ�H4 ��<���(�
# ]�r�kT�
��̏��n"��8��`֘�%�I.ѝhN0 ,T���o Q�ϼg�y�K�DY��kn�9F&q�|+�����ͤ�y
6y������Wcu84w�,��2�+jO3����td;�#��Q���Һ��$ǿe�VC��c:�?W���}�O��/��w�z-�V;m�4孴�'��(��0�}`j�Y?�Ê�,�dX�p�Q��)F�������Q۩�-���M�w���#M�����\4��(|������H/���I��F=e�N�~O��dma*u�$<�SFgt�#y�.5R�p6�����:)��r�m4��my���g��^�U��Hl����2����;!�)��i瓬��Nm�=�= �cN�?�&N똢���M{�S�a&��cާTF �!�R���!�a=�Y����_��UM�S���U-�8��L 2#}f&f
��] �����t�8�������-�]�xk�>H����<�$ �D���)Zw)Lo�;r�y�M}0��q��X$R
�+�B��MS��KQ1��XP&�*o����}�R�Snܠ���{��S���SA|�c]R��{�%gc�s�%���H$2��䘈Ä�[B�����޺j�=��˴ ̅<�M� ��ݨ�H�J)���=M�dmw�/}�/ѶJ�����%�j��q�]���ǷA���L�MA8���R�����|�P�\��B�)̓g{;UT3��^��$�ٹ2_~��=_��H�T{	��n��W��9������vq
)��m�=]��]?WQvP�.〄��Us�z�89��,i@a���'|.KH~ Ƹ�QK��`�"j�_��{��ޢ���?�h��[%Eq��j���F���G	�g�ئd@;`���߳vk�R�	�wKcA�Qq ���E�H�Յbo�����\���y�Fr� �'�i�{�o5��c���~�S��D�_��.�,��^?u����=�q�m �p����1���yIi�}�P�h����^UNUZ���AfȠ�_�g�whA
�Bπ��v�j�g��M;|	�5%cۯƣ#�p2��-+��؎�W�)x��׼��;�c6�7ػO��F��1#b��u�̠��ϲ\���eU=�%�I7o#�}�ԩ������j�I0�}���'9�� ӟ��r~�\�7�����Q�jD�d��?Nq��}$n|&J]@ѫ��]�QE7�B52��b�I��V�n������2Aĕ����Z��-�X��ǈ#�k��hI��3��|�8P^Ϩ�s�����=�|�kx�(w�� =jw���ڊ
�y�Z�Ls �O�X��2Q2�<����3�aR�i��Ѕ\mj��ڽlZ�u��"��bJ�$��viQLǠqpj�Fyh[��>�����6~Zu�e�G�a���:Op���/�qY��k�z�ì,�"T�%�4�$C1(_w�=�A��ˌ���+5?�A�{=��6�JL(�i���_+C�-޺WgF��X��ǖ�8d�f���腖иie�ִԱ�h0�� +�c���T ��~ڱ�'YW:��T4v��d�����l):�#:2UO)8��*`涗�r�YH���EԲ�8��z���C9K2ә�&����gZ������}'����6�w��\t�#���wV����!د��!��l2r*c�O��¶`Kr�xF�Bi!^�r�9��1��Ok�m91.�6OfI���ekC��M�'�7gƟܿѶ�u�5ٛ��<� ��+�����9��)p�=���_U+hYP.����쟀ہ���j;͊�*&���V��	�j����K�O�
�>WD������ s�M7��`��<��Uz��uES[Hh��d?9�����t|s�5�-�U5��}��Q%�e��)l
��)0���Օ^�	��P�Jx.���m�`��44y�a�K�E�Oe览
4�d�����5�r��t�:a�����<�?��*-��FDf�E)~V���(��9��}��ލc��=Et��y�������R�l�ܳ�T}f�~s��=���ڷ��(���ḕ���ߖ4H���:'�����	�<-�:3�Z����᰸�DN�/���$(��o���n�iP�h��,r�q�9,�3Y��u����9��Va�n��x���>@އ)IލƷjZ-�����
�S��[�UʣQ�\��.�* �'l���dL�֝U��^?���{�-]U��I�&n�a��+z��&�&U޽"�G�0>w|��\f!s��>�&�k��T��5�%\�Z�����h�sJ���5���H��`�f�{P۷����%2�9��/�#e��#\Ȉ��sbװ�_�r�+	�:��z{�� Z)��#&&$��9�k�IȖU���M��3��PhcI��atF��v` 7DFR@d�'�y}H7P`���%��4]�'[�@�x����[�МBw�6-T���c�(�/�_���u�羜;&�:9�������3~}��I������_	>�P��)��T4B_�bq^����5qla#���U��L9�RY�Oh�������ALw�H�͡��0�h��X@��ya�>��H��/���|x,��(�6��έi�
��V����5s�+�	+��u�����9�Ey6s�ˇĬ��[��
HQ-d�q�r�����v0p�k��Ns;�K���?���m�@�	+���ޗ�Q��/,(��������K�3J��u��PX�_B,.P.8�2��V�)��9Z��AC:�)���)�7���A<UmՔ<;���aL�b&$��U���H�sc�T�'^�����I�����SϬ��V# �:�!ϧ�3R�O+[����t��dh��'\-F)q�!���q9Y5����S����%bi�lR[���p�j�m��Ҍ3�u)��T��|��?��Ѱ�Bλ�i ��U��v��~�?�|���_���h]�1:�h���4j�f��$]��U��;�G����d��$rc�]��f�%�E`=��n`��}r��(��5z8�,�e� ��J���x�H$�O�9ɴ��q�h#���R��GR"�/�C��6�f���O[<bm��K���5�{΋ga�
�	S�1�i�s᳥���y 81���1�Y`&>m�_$���1��.�� ��W� �3�:1΢��~��J��]^�K�"�8��w+?}tKO�o<�Z>*��I��BO�rͪ�����+�bߛr���4tC.���341���Aވ�s��l�� �G��f��L�L�S|�Ejs�I���![�>ں}/8������W�����(!��zP�r�񁙈��_gf^g�G�Q���H�Z<�b��\`8���m��jD��Kc�hަ�<�Kp��;����8�l�z�ُ�`M,��B��~%d��Nw:N3����lh���ʣ�ù�z?6���YN�Mu�	 H�/SE}�Z����/f*��/�SG҇����o�.��Hx�u���Cl���n->Q�8�J:�G"����p��iQ�֨�m��,:��MP��2�G��ص�	������0�}�˝'q�|c�(%��)�/�� ��x�v�7�_�*p��#RX�Ą0b.�%�h���8j{��(F���g�Ia���ߒR$���i��^Ջ�_�����2u���S��H֧z�D9N��.���H9(Љ<OB���380Fa{.�e�&RѢX�.���/4
�KN��&	3T�:�����a$���:uN(p&���*ϧ��J�P��Oi�YV7Q]!h�(ef.ŦY+t��+Y�8o��0�8?K&��*et�l��$~\L2UL���[�iL��ҭ ���+K�{uq�M[���e�U�Nc���C S�O�DdLG��0b�Qq10��W����c��zvŰ�1o�) [`&� ���*�.?g�v�S�q��,?�C	��H��	���|�I�4�����G�!�R�4�Y�:���2�Ac���[/��@�����Ʉp�?���
U�	s0sK{F0�H�9�