��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf�&���>b��z�Pkk�ZK�P�18w^�9�u��0�3��i�?m�a�5�+���4���_����K�����x�}���0�$!�*WV��|xϮ�y�n��A��&�T�*�qY�q��w/������u!��$o36�7Q{"f;Or�̞��{�4�v�^��h$	��Ki4�,\��M��6m�PW�>�LCz�C���6`kH䦧�m̡wŬ,�(��ue��y+�j��?ՊĠ�o\I6lsj�S���I��#d E�O�F��A��#�@�!�#1��������--�=݌Q��*Ζ��^[q��MA���������M�����P��Lp]}ey1l��7N����-�r��C۟0*lv}C�`�]W��o�G}���.��ـ�Z��g��މ�����_��+t��`,���r���oH!�Y�pt��޼�ξ,[m[�嵎�h�N�ܽu�=�$�luX�VpD�@�z�y�l:S_�ݻ6-�н�=��3�?�p�g�r�K�nv���+�H�!)�EH9��1���[�[}Gͭʚ�����"�b|�V�N¶�Q���?�Gz����AP�S�`Ȩi�Y�7S/2�1нףK���@<���L�{f��|2VJ0��x��4�A��`�[T�t �L�)������c�ګa7��{�$��<T��/����1Z���<S��] ��USz~���T��o������%f��=���Uۂ���H��K�oxW�~�B`�T�`\VT�̴� �W�>��z6V6OԊ�R箸���ߪ;��t%��+�XW/W��\�&�&4���W��%A��oMw�]��6�֩��^<hAS�CA��"B��#c����V�o���Dߍ�5,}<����r0�B�����e�AJ�����\�f�|_$���8��]�	�L�W��N�a��bN�kT��S��
s�]�LR)�E�䜒G^,R#�$��9-�O���SI�� ����r���]�W$v;�]��mL�UL|Th.<�#kE	)�N� B{����׵w�f�]�׈v�%��/�[�_M�b���ڭˢ���p-:	��~�m�'�`�W�8�#K��@�k�a^�/'��_�P�7f���T� ]���b���;TѦ�RM=���
9ZO�.h��ʗ'����\�W�<*ULv�l2�]i��%r3���jY�󒤿�v���?��ҹ�{�	�["٘�rq@రF
L����?��1F��2s�+���j8�D��NO�Wi?Sb��hƻ���ID_���gv��B ��󭊒�A�]H�2���Iq�����^�AK�:�����
M��E�-J�nv�������s��HPI�U4x�١-4s�@@�H<,�1ԠiLԵ���Y�8B��Q�|+��N�D�g��e�J���rgŤql���	�ٴ:tf'����f"K|cuƗ�]}�-֫-�m/`_��
B.�ǰV�>�v33����:>��?�����Z��j9�$��0C��Ľqb詝��Q.�t�A���ku�iD���Z��/��s{�����B�vr���˓�(kJQ|���y!��nbr|t��=�$����m�j������v]���O���~���"	u<U�N.�TA+��vx
c��Q���{]Al�����s�Y���� }84�@���-i8ct2.��F�y'"��ɉ�uN�a�� ��V�8k���m�Zg��P?�XdU�}e�#�%����Y_�.�f9.��AyM/����1�������,���e�^W-3~R�-��F|R�c��{`~yS	Nn��	j9�$�t#��yg���@jЌ���x�8Intt���o���-�.�<�=��'!�uP�ϡ��/������&�Q�l�m���|ˬ�m��̀�(�����?+�@�e����?�w�Z����E�P�}�_�7\�h���ʀ \�V>]�Z����61�Ez���P�����b�)Rw���"Ґܮ��?7�<�U�8�GLM�yí=E�� �mʳ�o�N#c�;;����k!���)L�3�,���|])Y'6�_�&���p��k��QKy-1P���]�
�;�m�4�(?$�|�HQ9~�[9�}��ؼ�=��3�W:Z��b*�f*�Y��ӦԎ�ZhgHs�>���R����w�j�m��W��5st�z}�K�w/l)�4r	��%�z��Q�'?�Ɇn.�+U�>�	������}��z��ACRF����.�@���~s��t�f뭚J���E�X���  �>��e2�)'P.�z��"9xjK1�5���ws�!��`�#Iݱ�KM�_��1�aI]D��Le�s�p
�1cݕT��}$ݔ
��ܴ�8�!�yø�Y�y����l���#��%j^���͓Bз_c7�V.�q|�_Mo�S�x I?���J?�p�M�6y�(�/<�!}�T�@���VS�P��JI9��Q"�CSi��LXH(����	��Z8ik��
tL�/ڕ4�����a�>�� ��f�X,�����ҷ�E�y|�_�꽂x+����eu6{A��\^��u��_B)9�N[Q�6���8Súէ_;�	^vg��YS��͏fD��a�Ta���I3�Rd�};mQ�e������R������ܖ9��rE���lO-��+֒�����M4����_��6�V��|g�5J����זGEh7{���ͣ�N�sג� D�r��#.��~n��l@���g-��
o]L�6}�]�`�o>,[c���ҙ
�O�\͕Fb��M����^f/�,%U���ȍ��k�d�%�_���\m��0X�xO�r�����X�͓J��K�L��Y���S:o�KՄ^�\xʈ?��i�$N �3�c��$�����ax-+]۽���=�ZAC�߲ti�Z`P�=���ih��}�һ ���`,?�	=���Z�&�ޖq'����g�e?�����=���z)gvź����]҃ӨD�d���SL�3c�MU碖�͉A��j�e��hǼ�G��fQ�=m?�T�����]����fk���H
ºo�\m��֚n@ry�AG�)�u�5e�>�N%�E��K���o�8��g�be�6J�}���T����\݅��jP���Ji!�S��pvg��P<��wb�a�G�k��Pp�tUcD8�}/��>��A|��dG���!|6gl�����V"�I�B���
�s����dDG�>�Z��:�	_[[r����n���Fi��j���o��{b���@|4�#;Ξ�MVM��bY�;��y_�XE��_����K?�#= /�CG���ayݖ4	7�wG���ߥ V���Wd���Z��ك%� {U���P��g��l�h�Y��Q��S��@AZ�%�j��]����~2��������Mg+�ހ��B��ZJ+�d��2`�oZ�ꇄp��V#I��^y���c��vBG���vZ+�T����k��_.l�r~�b�)U�+��j��n1�q��Px�ECk��R�GP;�'Y�o?���y���Ug��[��Z�GS.��l)���診�	��|X���:Lj���x��݄�&^ Q�&��'�r[����B��W~�tJ��c���>vx��
طS��gX*~zJ}�L�T�{���zy(��܅�F�W�	=��N[�\�$>n|��z�d�q��v��)�6
���\X=����c�1�%��=�6�Tꩇ#�u��^�8��Ep��Tr��Q0���0Yi6�c���L��@�5�g�*�YPzW���N���kS�m�鱆z��:���'Cd�\������N�<9�-=Q;����ӟu`��P���V/�ؙ��?>�6�I�t�%����p�k�ɸ�+����Z��� ó�)�y�>���Dj#�r'�皿L��{۪s>|D"�]���藭#�����c�Lrk��~0S�2� ��ngQA��X�j�yPM����'E�{Z-��bhCy0�G{-�TL�l��EM����o�׻F�U�~@�3�3bΛ�����l	$�����)��2�*�v�0<�8e�b: �ZP�OAi\�%j���"&R|�b��~d��Op!E��oF�Bv
�)�����!W�������.خ )��%�����hgV����p�Jjg3�v��׏	JN*=�cJ󴹗g�g��檢�s�$�4|����"Sk~�S�ם?�%�P�eGK/�&jz�<j����A�o����K�u�(� ]��}nsz�2c���^�_��߸�u\8�+�\|�LcN���%�Dn���`n<qU��p�g"(d��������A'��t���^/.w�;�x~�:�w_0`�J���S�m8"�k_O�4D�r���h ���xH�V�����Ϙb������o��OkG,S>G!A�y���Ԝ�����R�Z�2:\�v��W�H[�ˑHw|���.� ��{��"�SDw?}<=nh���F3F�� ��$�����|J�>�r��Jś���l�i&���C.���VN��9]�Y�����O��i
/�$M���V`�'m��5��J��	��uX���{'g�����❐t��9�=T�Ƹ� �#���wP}�~mk.-����貽��+{�g�,�� e<�Z��ݥRbbUI�'y���^�gh7Jy�P���(�b)��$A�d;��t�5���֐,M��T|Ø|J�s�1avռ��v뻂����e9hRE�h��Q�� ��*,�w .��g���dr��+PF������2>nu$�:q?�hc��1��|���	���e+��Ȳ�����g^`D��/��`SM�����u�CC�F㤋��2�O_�<{S�v�S+[/�X�et������n5��=X�+m�[��L�%2�UD��~E��T"��F:W���7d�2�q�Ň��䥘�����j.K��o���z�-��ɕz��z��N-AlE �aA?]�l*u����LS����פQ�3��	�qo�6�;����-�@�+b�M"�S�P0�s��������%���n#�=ɦ�	��ZÒ���r;�I���[ i=�jv��QB����q2�}�"W���2߾�I2�A���w�#�f ��o�uO43\� �̔z��B K����lf4�C�&�p[*�0�9���#U�4���dr��/.߽��b:��3(R_n\�nq{��J�+��po�RIB}��/D:�]:�E�?���R|����^�������T2װJ[%���^+9���%'e�\�19�����m�T¦8�����J�� .�+���xN�?E���W� ��P`�~�F~�bʧ'��2P�[{F�o|��"]���k�ǛΚ�*xv�o"x�$�~�E�J�����0����S�\k�A�<��k�굶���&%�b�,\�7�"�o"�%EX�JХ�N�=,���n�2�&L�{zg���]X<�JGg���\�R��W�&LL��<}F=�{���ӓ (�uS�u�����J~)*�rW�\��j|pѢ�2�0<A��=H������X������V�܊7��`�Q�K�����7�(��&:.�dd�@�F��z�oL7'X�_an�R��E�^�auM/����R�٠(`��
��`�gQNK?��s4�����l
�CiKA�#a�"ds6Ǫc:a@єh�Gq 4Q$�����,��E�Ea�NhܼO��m�u�=e�����~�uيf]w��`t�v�n���WHz=��'�6߃t?���g<R�Rs�~1���Ӳ�f�n�Li2��^bbN(XLz�x$ҍ��U�WC8��{1?=Es�@�yr��h'�%s��k�R,�UkĄGbj�V���bxb�l\�����X3�xyN0M_���dj��<2I���e�&9�g��*�+&�ĝ�#���3o�b����B�CG�
hO*�f/:R�%��F����o�q��/���w���E4t��^}���o��}	q���}��R��
'��N�D����=D-�b�Pk����P�^S*����X��[�jL3`N����Ma�'�U���{�����-Y��)��@�"�E��WG��P������M�7��v� �%8�Q�wg�wS�Egǹ��`��d
xp�ڵ�0f>5S�n���wmO�"� r"��n��#Grۍ�w���4D��=�#�u��Mg�D��r�d�R2)��f�	1Ǫ�`zd;���ifwh�(�{3��#/j��������wb5oH{J��:�� �>v��>�[)��RvlPo�]|��2r����X�E���i>�J}�_�ۇ�˟�8���Kb�(Q(����@ѕa�q��������l�F�3&EQ��ؗ�����r,�7���x�|@,'��,�95M��<�