��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�^���x`�n�ɢ]�426���}�x�7��b���o�3�K��NK�z>�(<e�J���O���I,���ǵ��|ܫ��j��;�Яm���n�
�*/��s�l�O��wa��/�g9�	ܝJ��VZ�����k�$��y�����'�٘f��Q�h�\^�6�vk ?^"��P�_F����ٍ&��j=k�g̑��*��i���l��5���aD4��Q8~��[o4<}=K�Jٵ6~�V� в'\�QǬ��l�ʖ֤h�� ;�&�F��Xf���3�ֱYc� H�`�UPu� ���Ә����k�׫Am�xJқ�� A^jIi0��e�d� 9]Y��N�"��\�gd1�_r�K��ו:{y�@�ԅa���`^�(H��Ia����U����=���h�Vukܻ����4K7��s���(�z�vor��O?�b��n.bi	W�"�<�b��u$�2�e��n��������5F���{�Y&�^A�5�hYQ�?zO��RM0��/�c��J���_�q�O��n0#������:�Z�8td����?@��{@c�5�y+����ى\�7���p����g�+P7�!�o��^P������K:�qp��n�����E���1u���tJe\]T��E�u�����S%�A��q�@�Ʊr�3s�|�쬠�G��Ԣ�;���yV�Oe��k�B��
�F�}|������}a;��
�`��w���`L��y�r{�}��#)�pП���#?����<�u�Nd���#~TѠ���=���x�aÅZ�kl��Z��wR���9(���x0h'U��8�{h���N�+@UA����
ȥ)~2
��FN�x[���J�1�Z�Ԃ:�U;4�d�������O����H��;6+Q������)�ےT欟*��Pa9\���ѣ�	8�������U�c;x<*8�}�$��Wc��S��$�{�i-�9f��M�Ԏ�-��ptW�ڑ�w��f������pN\������2��;~��l&Vm���s{������@���@;�}��8j�`���zz���'j_^�âS�U���Q�"�1��K�a~,�W_�S�UC���꯳t����t�F2����2e�b'FC��|x|(�gw:���������b������#�N(B�lF]�2�`n9�Zl)Y�Q<z���H̼�B}�k+��k=s}.�AK���(WG���X3��22A���p?�B�X��Z:�oA�*��؟��9y��O-sǻ�.��<��$��~������<���,��7�6#��������������N֥7+���M� �̲�!��gT)�o�x�L�|c�������!P�os����dO�Z�>{<. �*� 3�dvV�x�)Q�<�2��l,c���J&�������ݻ o�"����5�q℀�!$G�᝞˫҃ӑ��aS�� ���c�o8ߟW��r0�$�Ɣ cm��5���s�p��Ms��7<J�`����F~fҷa9I<�ǆ���-�37:R�B�ċ:��"G4``�ǰ�L��ߢ5�4XEc��\bR�SO�`���w�������쥗�gB�����\:�KU�%9���u�a״#��hB�,����6bo�>^1߀�f��cx9��P�u�jbM�i��G] aV�1�ր,�R�,��K��֏��&؞���qH�t8��y5Z/x�dI�@��k�K1���sK�v�9E�U5��F9).������ӊg�n���?L��O����?�l{���>6Ծ��!�N8u��(�L ��rz�Mpz�r�pn1�;�`��= s+�jŗiۛ�=!�M��iY��j�+��O�E�l2[�����,��˰î��-"�M�$��1A��*< �K� n_M��q*x��%ZR�1��q�����Wmp���S���Zn+��e�Q��<�'��bBE�goV��"���up2�Sa�Q��,�j�D�q�����J��R$��޾�@��J�����~C��(�����L�Ů辴��0�o�Aj�ʙsA��J~��V��hѻ&Р�FT�Eco1�,�{��T��L�yc�P�1-c���__��,@�����y���џa�������C���'�t��a�QbV�~/��k�W��Ҋ�%k��e�Q�m�<�V✕T$������阠�6v����}���6le,�=z���V��ٟIo��|�&�Ђ��^2�#�᮫�B�b�F?�rmi�m7��X���R���iL�A��ٯJ���ݤV1�Q���Fx��V���'���^)�����E4cR��ʹ�6}{-_J�S�2
bzW8J��	��������bPlSE4o�|�{lS�~�d������]��Ep�J�)k�hrU�^*�3�ɬ�D1�D�i�)��}UR�t%�Se1��ʎy�X �c�X鮍c[�x��
j�2�ic- ��wLh&{��%�g��v�3,��=����#/��bo�RQ��|����L�q�laI^�b����iF�q�W�~K��
�T��JD�CX�u�*��R�4z�����Ǩ6�H�����h.��������n1Ծ��[&� ���E��#���u
�(7��nz�:3\	�0�Q����j��:���	p���;I��k�k��I�t�+�[��_X�����	���y�[�$�d�\egDPg�~�d�
��hC�ɼ�*ȵ;��Jf;���Ty�ON����zi���^X�$r�H��VdV���Ӵ�GRvD!፼H��'�yD�D����-�V��� a%����V�����8JG6��}��R���mo����D���N@���Y�%wM��.c05����W.� �&��f�o����K�MO�%�:J�!�ѧ��Am$�a�R�=���Vp��r���?l��x6�C�I2�6��Rs#.�ޅ�b��2�J�U;n�n��c����vb��P
Rә�I��n�救e���9c��L��T��="O!�o[��>Y�²xC!�lا^��w��̱��Q�<Uo�n�Tܰ�h��ڻ�2I/�>I:U�Y;(�����P�G�s�F��J�) ����Oׅk�3c���A�@c���i=l}� �����ON���ɩ�++3#dy�Ch{H�ط���jo��7��������wr��֝��3%�;di@&���3����빍K�2�Yj���_/#4���4<�����25�?�u:e��+B�b��xa�S�(
F�~���J�&j���<�Pe d��ȍ4����R�u�T��If�9j�e�B�Q�T���)[�����R�ݔ�����;��֤��(��w�kD�
��l�Kyii�x�mEh1�Au�̀ �Ʉ��sHh&�S��Dd�O�[ԄU����D�40���V���}nnF�Y���_(��i���vH�m�z��&+P/����2y����iZ���	O�;�6��z����w��
+/�ܿ��U�--�7%��}b���)ω8��������u��]E}-�Β�/� �>܈��I0E������6�2K��䍍�J�N���2u��(��?�,j<x3t�-�mZ�7b��T�u�*g����S�47bM��25l��t�{!P #�!	z�j�X�ͼ�pf�5�ٕ���o%;�>������� ��Q� �:w�q���$��R���]�^@j�%+�4�Qu��0(���ҥ��dt��E�K������&Y��5��Q��	�z�x|C|sxfS)��������ʯM�PP�o�["�+�0�.~݄�u��@2
�|���GT���)����!����4�M��d�ǧ��v}a)��x۔w�-/��X���ǟl�A�>�-��¡@��N�>����R�(���D\^�?�>��S�V���	(������f�a�K�5U�;3�DIo�֧wU���L�Ｓ���y�"K��⯌��G=ʜ�hᗆ�
�]�"1?Ƀ^�1a{X�[~ڏ(��q��Iq��gn�B��2��W�Jȭ�)j��O���[�d<��R�=ɀ�wS���-�
Q[�]=U@�����JJ���(���eE)� +\]>~t�CI�%�zT���%ӭ|n���m����
6=�ecU.Ψ�A�,y�lu�U���0�)"��xK�S��Y�*�䓒�6�*�`P�*��5Ϳ�K�m8��πw-(�C��Ǵ���]wqP���o�6�w�(���
���ۯGȯ앙~40*E62�˵}!eP�9k\�q�}�w���q���9v��kC3-��+���&�����[�@��#Z�^���LT7$�����T����_:zG*�?F�S�Nx�:c�#�,��|ᾏ�P�`������qC,��jۅ��W[W�K�U{��z�vD�葵�����S���TR/�6/�cɹ�}��f
C��b���>�3�⍜���:{��� 2��@��E`x�T����N�?2�`�P�E�ꌗTZi�㧧�^���WgV�Y�YW�7�Yӆ 9Ki���
�U����Zw���˱@�(i� A����9R��iUIG��#؋���7]!�9 �Z�� �~=��qt^�ׯ'J/n�o\,�)~q��Yep��[:vK. ɑ2�=|o,�EhQ�:�����{5����K��A��z�Vb[��VK?ܯ%�	L���k��
^-�X	ǒ��H�M�`���_�7�{sU���V���a�5��,�#������L���y�SN��<�f.G��9��a�.cw�ɗ�1䷨����4O��CO��h��P�3�IhXL�>�FSQ��Zw�v�ٕ*̢RW�Zly��Ċ���d�gk��BN	����w9~���Qr�>�VX�{\��!~�_#^�
��3�CCY����ö;�Pk�:|�B��y�*��:��-�g9fxs���_��c��/�BZ���F�&fo��8Jʠ�x�jꍐ��$U	�U�mp���v:���|�t��b컘Sr��{H�c����{������'z8�Q�lZ�uJ(`�ŕ��Ґ���fFl� �Avw�K;�u�Kܻ�hh� ��/ _�%J,���0���ΈyIQ��l-��!�
7��4�M�:��hM\�ڤ	���F
��,��b����&����O�C��м��y��$���F�b{Vh����E���*�#\�}��դ����*;������?B�X�+F�ڧ�w��wA��)�Ӟ��x� �'y���G�(Or�ח�Xmu���T��HŔ �+iS�H�b��D4�W�T�`FD�P˪�"����U#Z3ϩ(��?ۘ?��4.$?�N�v��~hn�%� -8��ԩ�=oӈ�G��14�	U���"ATK#)<Y�M��$f��)�(h�h��0;��q���4IPC/�w?g���aW���4�l��>�����_c�uau��jl�A�^nu6L����P˄����!E3�������Ѽ��������Οa�0��r�p�|=S�ꔲL��'R�"s�[.QG��R�	ͅ�$��%`�ʦ����h,�޿D2m��ǤF�֩�aY��؃���S4�cʤ�2-9BƯ>�S�Am�t�*V�fy�Ly�Cs�@C�)��n�`3*#�8�}4ު�_Q?n�eci�EA��?����m��ύz�K�^�i��_���9<��;Y��|�x	56�5�U�L;5b��f��c���}�X-�{��mN36���]u�稢�(��`LH ��z�]\���@yDdHx���6�!ȥ�2ɶ$����B�A�nߚ,���Smtn:D��e��K���B�[�"H(V�{�[��e�7Iz�Fi~Q$1ZA9���d�Bs�/2��d��S���u�`" .j3�4ا�J�A�Nl�{�f��Э�����d��]�+���o*�R���t8�z&!	��q�E�韇m0���54L�
�z�`��� ���}UGh�NIo�P�����b�=�$���	<֏��X0��|tˊ��?�|}� ��y��P 3㕬ٸ��b��񺤦Tp����q�/
f���(k�m��G���
^f>:��cO; X�<WxI�e�9��ox�*�]�dZ�S�f�I�[�"{6WWp�\F*�|�!i|,�F�"��L�w���Ф�dV��m ���c�6"��5P��R��b!גR�G�*XE,m M�>���>��}K��ǋe�����Ā�v��?�����-]�^�6��Y�[���	S�]��d������_��湤ϘX1��=�b3�a�?�d�� G�kN}1)��;:dyͩ[������1�Z��l�WB�=��O`�P���hV�6�i���*��=��옌,3�]���j+��=�3h� 4�&��}�nưXL��#ު&��Ha��B�5�х����ap�⓱:Oё�&g���N�2�d#M�Q]y����n��-!�D�nz���zC�ѓ"��G�c�A쨥dkӸy�ǒ��5���7����&R! �������?#&������'�J��`Z��μ	�fLXK�5���X�b7�� <���u>���������I_νsi)b}S�%X�l��@ШRrb>;�<���}�}�)}t��D��`-'z| 4j������Y�"J���s�iZgc���T�s�iuՖ��q�h@�6t��������O�;��;�)��iKn�{�e9�5�����X �F��\��\�h����͜��獨�w_����b8�g��OJ7��g?&�[9wN����!���"wK���|9�W.$��B�QB~�#�xT�%a[�m5w<EՌ�젊���/!Sa۠�_@ö�������55_Ho���dE��Ԫ���SI�����Q(3Uk��������J�XU�N��J1tT��w�H!]C�kݍ%�Q�O��`Ѯa���f��mG���BC�!ң>����~��e�v���rZ��Y9��/>��H3m��X/k!���͕~Mœ�Hj`�
8�W�ٽ�Z�sz�/5�G,�a���F�ͥ#ytm߁)��n�,����~��w#ca6(o�~8����^o0}���:T��zi���N@z�a���2@���"����EaoB���I�0V*� �năK
?ݾ��1n��.�W	s_X!�G3*IHjv"#���i�D�S��q8f�BqS��2�x�����'���4�u�R*�z���s,2��7>�"�sb1aǎ�G�wx2�h�F��%U8
\"�1�5Jv�cd���ȭ�<=QX�����`�7y$�.��2Q�a��Kxb0��\y��g���ae��V7f�q:�s��y�/\��>#����y�C��d�ƾ�="��"�I���	Ob�� $�3�G��j�W1�;z�Μ�E�]�C�E@�d�p�!O�%k#NC������2,�����5A���r�k��0�6��ʮ�����"��9���3?q��g����b0xE$�(`Sӽ4C'R��E�J��v��
���_7����i�C�[�掾"��M��e���	�Д� ��4N�<ŀ�3	b�m��5��0��Z����_R6��DѦ�5.B��7�(�(AVb�P]5-9�l�7g)n����˭0Ď^�����C6�V��W*���H��_�b|f�#�Ð���&Q<Jk}���Wᎆ��-������pv��
���I-�|��/�C�Ն�����zK�ڟ1`�H
��9���cԥj0^�~!�*�M�ͻ]��t{A8>�c$��o���gz�-�V�f���ل�]1����\\���.�aQ�gA"9ɽ��@��Fdgm�j=��]�ޤ�=1R~ (J�7΁c��R�B1���l�Q��T�ÔuT?Sz
�֮8���
e��E�.�
��s��;���x8A^�~�5���v�0�c��h�It\���jUU�G
�YfR��C�0�5{[�������!�1�6�m�e�7���zi�=��
�(���f��Ja�^z��	g%&�N+@�e�|����W�t�b�j�jB�7.9�B�#h��d�����I%�f���oudG��L؉�`�����US����;{Bk-3Y�6� FK�N7�m��[h�-���W�3*��_K��@��!UQ��!\i��"��T�*g~Q���kTr6�����1
�R|BX�HLK��L��ʾ���8���x/�8:=z�my��ko.Q?OE�<���c�Cu�s ���ԛ��+[!Sqt�]�J���2���։uK�	���_Pngz��EMX4'�߰G
	�-o��"���;qF�,,����R:?��Z���!{&�{��*�h kZ:���7�l�!������NH��Mg�ߍ�+v�7F�����GF+�ɤ�6�Z��لI���v�-F���N�`�'�!,0�@Pjsv�ؿ����'�v�P}����1�˂�p}*�m�.�	I�ā��د��=u�ęp�LK{���\�l�ŏ���
�I�� �c�X|w-!5��׀0flD��&}���~�}A�DWΒ
Z�G�(_�T;�(y�W�,�쑝?�.��-���d������<1�/"e ����`��`�>|��?��1L�oF���L���|Gc���YK�nڛ��]�(��~���Id�jUN���s4h�5�tX�xc�D�t4��Y^��Y~�Jݣb6C�'9��}V��])�8 `�{f:�Hy!UiR�ʶa�E(LN�.��(�j�k���s�|�B����`�tF�����/%7�g�a^iyD�ط�L�_�S���p��gH�.O�o�J����$�c��Dc�Fj��E�o4]2$��/<-���M��I� nTĳ��OP��;��4�2�mG�����|�$�K��h8=mL�I%��av��#�{�dI�Ie��E^�Qse���O���?s�����g6�
�%�ȫ8��H�f'��2��5�yBcː�����s��0{@�va<��`��e!3�r�;�" �$}4]��~���^�?��JJ��� �h��_�� ��4�o�MI�Gf���:,�_#de�zܨǗ: 9q	z��hs �7���^2��]:rN&��&���4�P�a���)~Ԋmm0����Ǫz���}���嫐x����i���|�P�T�x���{����1#�5%b��P�-d�� �ޖ�
&*���'��g���nj�%Xm�؛���zR��uڱ������.��q~�@�#i:�������$�X�#���ߔ����Ì|��͒��7p3M�ɽ
�6�Q�vs���8In�1�Z+u�>Z(�W��y����o���H�^�(?4&�pv��b���,N����CI���a��A�J@��Q�C��1Dt];�@�G�o+���(n��\,�Pf��u�jT��&4a��G�n�����_?!-���a��X�=���8��;6���:`�ͼ7.+�刡�B�s�dJ�'���wP��)�"�e��/�A�09��Ez/�
Ր�zF6��淌N�7�H�=S��g�R��|���P�S�5�p����)���ɇ��P�1�P��d=2꛷���i�8�k���g3u���V[�iU"��"w@i ����7�	���4t���͹���M�h���u��*�?4>P��g�D�M�{�7q�w��?��luGy�B}%~2��1z?��9�'b&��o�Q�G��C=���j��N�m�s1rы=w�_����䂑�J;EU8�wj|���y�N�[s��veݓ~�GBL�����VA�ވ���lM�v3�3z��V֌g �_g��s(+�Bz�`�����4�1�y�5��>AT���I9����)��WT�?�(�U ��g��b�`��ǫ'�IlҊn`cLT�%���䦈��C�b��N��<��h1+TJC�J3���hK$q�7� ���s�m�mE�Ee*���f.�Gw���:T	'�V#�2�`oyB^d �0�2�<V���AۋE���	���+#"m�d��ѼĻH)D:���㍪��~��iQ3�Й�X^���<��|~u�C���y�Wi���5��:G���X/�����ҫ�R;E�F"�L�^K�uL��R��1��<>0o�E�7_4	��d����nW6`�Pf���Z`_��4�+��~&���[_�c�{� *ҹ��k���e�D�;��&���C���#��t�3�����.�ώ�cp�=a��X����@��p�T����0z�1L�d�J�{R�`��#wȘ��I��!@���Z�hх�?�|g�3s���:�����'��𝕻��H�,2߰ƺ�P�������%4錽���J���(����..�ǆ7�^���~ xTJU�6ñ��� ��s�	Q�<��!����2�C7i�h9��O|�=	� q�"�"�d#~�E&Oo��F'kV���N��Jwo�C1B�J}®Q��w4���"�~���A݊�w����"���b��b��!"�0�\Zj�*�����V��ElE&�+�y��&K~E\��>��M��w��S&F(C��������&�+��c3|q��G��r�^_�&oA�(�A��`����JF�\�hr�� �0�t��0Hm��t:��S̑vm�#YNt^��;�~��
���Ɵ:jf��>��q[#ԄP���}
�*�q`4�����S(�Ǐ���G�.�t�O�t�˙�����"i[*�8�m��5�B̵*P�Vܛ�"aX���#�~�A0'v��ҽ�WRw��}$ yO3�w�+gV��+A�qp9��Ny���ɔ	��cn<��3�hVE\���*�O��/�|��g���NTT�MI$C���䎪�r(؜'��& �4�L��GiO�vc�=;-3mH6hU0J8�c��Q�le�OVi#wބ�Aw�k�s��f����%߾'�������cjS�81��/ k�����W�[���<9�v�e�6