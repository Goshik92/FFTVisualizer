��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�V��:��X�o������Z�t��)�$�� ^����hZm��xJ��}fK��pD_����;G�)��N��h��`��Y� ��v���/�5=��*�.�(�`V�\�Q<S�O<��}iդ�o8P��V^�e'�g }*MQw5e�]�a�x���gw�W!^�a�zqq�1�H�<�E�чA�"�:��,��l��
�{^��i7��a�Q�W���5�n8>�}�MB2)L�on_Փ}�,^0�O����G"6^W�z�Y~S-�k��S}�	�>�}�`����2�[ ��:�9��M��>
*�T�܀
�~&
�W~��3h�nr]����9$j��l:x*�y�s�3'�ch�,�W�(p��L�u9���
l9�?(��1�֒��;�n9ITZ��2=���0{�$yy��S�-lԅ�0��؉gG]�T�t�cW���`���YL΁_�
M�2��TY\w}69�=U1��<{�W����l�`��+-��D�yڳ��.}��ڦ�?�?m��j�7@)�2���5���U]=/�H���XlN�e���SO���8��UD^�$B�c<�k�MK�	��d����;\�nv9;���t#;�83�Ds'��7�ƴ����a	ѱR&�C��ch�Qe�&+��`N���{P<��Ђ"�Ϯ�Ĩ�ȓ��!Co+���~�A&9��{���@Y.z��0Z�M�D�N�-a�..��2Q{��(?ӹ��_���$�?}:��z~��nt*��l�
�L�����	��^6<������?h��ޫp>���Oㅽ삑�ЃВ2P}��щ�{|�Pt�	����83����=Ҵ䒮�Ņ��d�D�ZWs����t�}?P��i�1�A��A*�c�d�S��HÎ`d�Nr\ET.��0Y��J�g�t՚�w��g��,�����b[���R?)��7�T]�Etc�~�fb���H'X�n@Z��Pm{.y��v�hw@��	x^�vZ�*��U��0z���ڳ 8Ӣ�Ǹ�gz~H��"$q����)�㮷(�PLe�%���{�n-�b�ȾW��d*���'�H��[p��"�Kth�6@D��S޴ͫI�?�-8���ŝ����� f�94����V�]���'�G K�^�m举F&Gx�%��,w���&TaW�Ezx-�{C�I�I�Ф� 1!�-�ka��:1H�UHpAR�IΚ%�8�(�8;v�����]���ТtlG�\d�Hf����jj��V��R�!q*��m�̂����̬�O��&�6M�xe'ޔ���W���}[��`T���l%�v�$�p�4�ɰx�Lg~{�Q�K1��Z��~�x���D������w j�bG����iЬ\����]���@�./¼࿥�D�K;2����^ٶ���8��bzT~jwu��}��&�m��l:�:��Y�k���"�Q�_ ��Ԃ����oP4<	���x���'wA u<
�䒊��M���b�u�ө=��r�mFy����v�y�:�/`	u�=�G��ƥ�K�L��
�@}M(�P7=㢨���@�wb�[%pv�h�$���႞��SE;��ͽn0�NP�2}H.�o� h��@�49$��������\Z�d�A�Ț�����&K�Ƙ�-{g���B��J3�8RT�R�
��1$.�b���sW�o��TGb���_�\����|;F�:��&���ۯ
�-�SB��ۮ�^}��*��,�����2����PAuv�C��`���0ˋ��C<+������]D?!�BO,ts��7`�{R$b��Uf�f���Ws�*�m���<bw�j�c���`
H�3�����<�{�����]P�'(���t9J����϶��$��.����$=.9}��qq<�r�-�O� ��l�!4� ����.N��|��
Lޑ��7[�Ib�{���90|�7#�}Aݯ�բ��F:����>�iЏ���t��"����Gm�L�ܝPud�֠^f_Z��w�{N�;�ӱ�����5���'.�����~P��ߕ{$�֐,d��)H���Y�Z��s�걱�/>]�W�P��
��m������xhr��wK[l�&���T���tR�8����<m	Z�2�B��0�:�&#���J��V�r���|��kj���lof/���{�\. bN���y��| ��bo����l7��mhs/���/I���������s�U�
�ee�G���;��N�k�t#ܶXz�+&�����a�;��WZ�߄�d�A=»=��̄��NSc�w�u-���_\o�X��H�ð�.�?��7�)D*{������+����s	�T1胧����S�,?N��l�!��Y�4��\�i��~�s����1Dxߋ.Qb�ц�7����28��thʏ"��[��&�	n��3kX8e��U�>e��z��y�C;`w��!CQ�&����1��%IseMx}��K��7���i��8|�����)��x���Z.�A�mgUj����]N+���uY�iEL�~_��tLJI�9�t�:��.,�ˮ�N�d.�7i�o�((��sT*FI�b����0*t a�0"{an-V�\��J��e�1ͫ��}��/Rk�	c�,-��5��|=��,a���� (o9�?A��x��͝R�н����9�u��6󝡻6�4�	ť�]��zx���9F��J�/� 8;r�N�����4$�(Y8����^C��c����*qRq�P�>�t�Jݖ���C-��y.g�}�])��%�ܱ�i� ���g��)h�Tl�{b6~7Ҏ��{�.��RM������IP���d�RɆ�v)�H�D�`u� N�nMe�kI�ż��)�Z66y���P���È�%b�e��rS�~�=E��٢�B�İ�l��b��n�(\qA��_�VK�
U�SP����)(�6�N��A�]����,T	U��� �v��YL����+@7E��ZA��kᲽ
��@'�,�D���$�16��M��=�+I躿��b�� ���kW�\�V� ]�~�@V��T������f�R�6WhLM��G���.K7�R:��-�(�=O��S<�L���k�Zl?S��F0�S>^:�^YIŖ�5\����[F�H K��J�4-\G�ī1�<���s!f�Q(b�+�e�T��1=u�dZc������Rt�#9
�7~m�K���!���Ɔ*���],/��Z���z���v>֤v�&h���++�f�L`jf�L�(�S����e�#c"�������T�-��Fe_���)^�_�>�N.3�ZKs�b�~I��������_�'�����V���Bΐ���O�qD�,a=Y������l9�� �N��#l�\8z��ϳQ�B���Rk�-�p��D�W��-��l�q���C��qшw쿊�O��c��s���f �,�ġ��⵱�M��6���*U�F�ʘ4x0��mZ���D���U[w����
V_TtI��)m�ۦ����P�ۣ4W~:~[�!���X�dUx�$��R��/���S<�*����������*��\q)��,[�}6xEb�?y�b�甤0�0�h�����3�f��'��N��tU����|��Ћ����%��y<�GA�����������m��>��S0���l�K~��`9���{St�.��D��_��0 �C�eL��ա��a^�ן�2��ڿ� �R� ��� �֘��ֺ!*��n;�X^�h`�K��QX�'� V�g��Ϊ�9�;���*��_�1u�i���Ҵ	�\��~*������&]����	:$3J/��4�4-Ɗ��g;�|��3L5��4
��F��r8��@��\0>'��:h�D� ��j��D��f�G�Î���y�̸�E����&-�ŀKͬyCAtV�R�e�e\��2|�E��x-�*�y�I�y��w@}(}�2�*�6�~�JO�jX	o��u�F\�8	YSdc�FM�g�`��%Z��`�N�{W�J/�2�_l5�����&R�����-"��
��|��*
b�8��X<±�������8^�a#7[�c@�*\�ǝ��U��jטUh�8}l��.�P��w���$d�|V��рT'�ar�%��m�d�e`/��B�B�j�K5�b�t���28[P��Oī^˶�Y7�� +:�ekVA��8�����`�%��[�`��$R��k҇_��ʊ}��M PE���re�I���0u���nY����ߐ�,�-�:��%��� H�G�-�<l&1T�U�a�GX�զ���ds���9����s!h��<��=s�!�<�T]���u��X$�`e�^7
��h�'�L�����S��By�%�S�>��qFPc�(��ID��e.'D��=�w*+�u��oZ�g�x0�� 3�ּx��E.&:]T�pj�cKx}o���@'�8aΞa�݃�;Ѿ�3��ݶF���J�[���w��:sI�("[U����[�
o�S7�O��f	�YD�9�o�2"*�F�aw��&��?x�6{o�>ќ����%��AIf2�3�-�j�1��ޣ��N!���s0�S%�$��)�.E]jlZЬ�I�P����LUL���q�剣0Ib��СX�0��Cd�Y�+�_�:ϛ��j�!�2�6�/���:��g�-�J|L�K��d�\������a�9�m[8�ywL�h9�!e�_;� ����-�>n�3�K�h�H첸�����S8�l=M��7����τ�!_רcV�u��G��"�d����n��a~��������ƚء�H�����jS���p�όr��#�NtO@����'���%�����c�������r�H���@�\�o�OP�
��%�P��io�b���d�h p=��-��WjC���ʋZ^�Tf�~W��tr�B��_j�E�s����z�;��!�̭��!11ޱ:��;��D�K�̀d:ST՜ͬ�GnP[RW�C�&z%�cE�]c)�F��{I�Q/�=%>˾!m�sa����rǉz��b����/$�+�"����`��C�ݜ`iR�(W��#(�V�C���L�H�#Ӧ��7��[���F�W�����ف~�~�����K�$M-'�z\�-\��Y} onW����Mk���� 
�=�8{!���9"���"
n��q��#FЁ��'U���� �h���7\>p�~&�<��R����U��%#jؐ<Ѿ�i����`NӔĚv)NO��GNװ�Fr)ץ�b��r�����B=�'R�e���MJ���u%
]D
�'`�C�i���%V̈́8
���`�B�����&By���I�$�a�����:t<as�6��� �k�/L5g:���ػ��<b�! M�]IVk���$ҿ9�tyrf���WHqP��N�f�SE4�e�a)'=Pr	�([H�.�"��>�/rE�y�Q�_�A�aZ5<���ґiI�r�7X�۽/���U<�id�^�ig�So��[���37u��Gp�l��,�b�=7'�+D����z�7�廪��&��^�@@DA�u=�h�c>�)&�	As)��)xUҀ ��CH�o��b*�y�58�q�����qi�y<��SSj�f)w/��X����5E�m�����#���e�K�c��*�^��ƪRX�l���\/X���"�Q˹?���
-�=ͭao��>��|�P����VV-�Я ��nƩ-�bp�4' ��ȇI���z�����u�q��~���Hyk�v3�yc�H1j,9����"�l�c���m�?��8��й*���+����&�v&e|�V�X�
�~$cH֊W�c�����?�+X�I^����/0�]q��8��p�E��2y�,�PΫw�h���Dl~�E{Km�ХP	�O;K��r���� ֙��6{�\��-N7��qk��:g����H��e��nL���*���4w�� ���ROu�1m�"�֋ݵl����!�~�?�z]Æ�Y
R���P�Na�{b���3w��%�b�P�&R�z�Z�{�j�Zl�A�(�e�;#��.��ա911̑v��g��	��b�������0oJ����k�~,��W`BʚU�$���?�и�XV��	/�Q�\���7Z�t�H��"��H [�o/�'�j�J씸�B���%7d㙊y�k��d{�m[��D���[aq,z��c��2��+��ɖ(��v�*�J%�7 ���J�T!J�:@�-h 2�f�=��Q�jO
m'���6������W��6>�c"y���B�s��`.��	�}���jh���'�m���p3Ȑ�"QZ��ћ��]T&6�j4��������i�?v\����w����wIE�	��%��	��\�Z�{e�[P�>ɡX?�pC�x�V�u�6	�K+ bid��)�ڤ&�Nbr�CD5o ƍxז"487�z�y8�-#u���d��vn�].㸆z��Gb]��JJ%����B;),/����1v��hZS���^`�bo=(kq��V٦&d��%(�Rw�����s�#���|�Q1dߑy���1��7��z;W]�v�,��ǚ�G���_�rn���Ԏ �����w7���-���=0��	�zP;ΉmA$o�����1*�k��5xAz�'6՝���SC$>�BQ�V:���_�pi��$U�{�#0Df��o*�����?Vӭm|���8P��*�>��%��($-���̂3J7݇h�&l>j�w�j!��*�~Zg��]�P��
�n#`7���mZ$O��Aep��]��!��C�{��ф�s���)X�r_��{���G<�����{���%�����_��~�{_�x�"�=��(���6?�o$�O'C��8Z%�JU������(٬��:%]�ő�Ug�d��
�����dE�׉<��ݽ��5�Z��_C�ޟ-��J���Ue��� ��So�{J~��}c�!~����� �`2� #���N�����[#,OW%T/�+�0��o��W���*c��F�d��_�{�������-���M�io��ה���'�?u�{)~+���%��G���/�,[8[��a��=Y6�U�7�~�CC��:G锣��3c��Ԫ�Z�j��d��������{y��3�U����5�� �����et�e6�8�@23Lyfe'c��c!�'t�5M���X�E�`�MޙaI#��d�^���������!�,p�Yu4��ˏ�$��94u��┉~�Nhpϫ�o+�*Bhw�j)U����KY&0=0aty�>��3�)�9�\���8�S4���<��?t���+��e�Et��I�I��uO��F��en�9ƹ�a:��/U�2�v�4Mw�\��`��SY�Ka��<�ە�]sU����y�1�Q����d�7Cz����gz��m�	��� �F>@8�^�>����4")&c�R}���"�������/�[C�VZ#���Ɖ�0��g�'���i�h�FC� /[���⨏�Ѯ����A=pe|�xr ��xk��ľc:5��ܢ�ie�R����]iw��OaD�B��2�0p�o�(%8���O�����ɋ��׀JY����}�J�n ���U]3�s�T��05��Dz��L."��#����!�D�,J��k��hO���~����#{al, �6	/|1����><�X�5L��7�^�W>�������2���9�4�U��Ѭ��sfh] D�*�� ���������:��B�M�Xp�c��������d>P`"�/j�j�,
�^R�{)~tM�A�)ȫ&�G_VqY����^�,��r{Qr]@
��.3:�)�c��ȭ�����ڦ���BB�,���d֌�}���W�&;�K�g�n��8����Tˆ�ޥ����� 8��k�����"�~h��E�YR8/������YO=�ڛ