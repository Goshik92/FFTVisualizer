��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M��*����g#φ'����T��6%.^f��8{�^v�wK�T��fAN(.�oC�Yt���Ao�>���� �h�*��9礩[s�Tj˧��Y���oG� �'!�D!�#S��E3@b����}��(��ѣԿ���:+��rYV��;��6��!�iG�{#�Rݕ_����JkK�ݽ4\�(��.*�[{��+����3J��� ���J�S��pթ�`�]JX��X(EЊ"����sZ�Бx���
�Bo\Q�t�����vw�ջW����ccσ�*^���%l���N�rd�!����Z�q0G�nRu�4Q� ���������㜕�f{$u�6v���9,(�)�8n��N��	���]� ŉ �"�'x�Ε4�
��=cE��%*�Xϧ".�Z�x�Ro���[":��id;K������j��QU�^m6lr62��qʛ�a����� �Oy���,�BW1�P�6F��<�ot�?�������PH|?�
����ӳ�|by������#����OE�L�w���p�
H��鱂��M��cZ\�K�L?PQ��	��脤ѫ�ARw\~
S��ҋ�24��(� �.(g�:囱= �d��0#mw@�!�Z��4B.�6�X�ИH?ー5+�SI�]x���dS���^��n���Pq Sn�
��0�y*��8�O�	�߉"E��s��H������*�����s�Й<���:�&�DD��j�Y{��◫�ڧ��b��PǩғŔ���\��cc���Y7�T`�T
aaq�g�_)��m`�,� ��/�D?��h�'��PN�s3�ܼ	�i��4�y:�	�Cٳ�д�?��'9(�]�������jZ�L��5�{3k�	�x��շ/�#'�u�]�&��)��:%��p$v�	g�jUIm^��ߕ]ޥag�`�O��Ia�.�h��/��el+͆)XO�e���<J�ͨ4� ���R�笨s>�7�����@�u"�;(ߍ3�/��뺙��k��amc�Jc�9M���h���*.;8���P��Z_q��q�L_%����"�r��9�Rk�]4%�(N��=W��e�;�R�*���81jC�b�s��U��+�gJ�#�$�8a���4V� �1�9��
�	bv�`�"lJ�)�}T5t�Ѩ�Iwe��.�2hD��r������K�s�Y"�r�שB�m���V�k>�UM�6�ԡ���!�2h%"C�RJN=��|Q�&TA�};�ma�U�)
�&�с����m��4J︦:��J���
@z�5���H�s�,�l��d��b�s�lMM�"}��C�k m-T�[��OA{�)�V���1DAg��.X��[xL�Q)�������A:�Ϸ6S��9?Q���BqM��V>ݴ����_^�^U�I�kn_d&��J�� �.����i�ǹ�;�_��?!G����1z
8�L�W ����f��V���>cn1yV �$�%ո>�Ǐ����:Z[]�VX�z�Y�)W�,�#n����~*#�u=F��. ��K2�`��A`�?ۭ�q����� �lP�=V���?�?M�ɭ����`6q����Ma���k��ZԿ��ِN�v`6c�I�_�~7<�p��qf�Ie�Jig.G1�]��<�͌��/�'��ե(���?��b�(�v�|ر���������Qܼ�C�[.% }f(UB�-��7jq��'���M��$*@ѬV�z¬�eΗ3;Dߧ���D঄����sqN3,,Ʌ��FĜ� ��eɪ'����sz{�
O�n���9�-ρ#&��vX:��TZ�UMj��#%LA+�w�T�T3Q�.�+ϣ�q��(�T�%`J�]A,�@�̞�VI��n�E���=�M���oz�v�{b�,�3݇:��[q�,��0/�x���|��stۢ�R4�p��)�X��+�n�iBݲi�h���f���C�=JÅ�틁�Q߼\�h;���$k��s�'�L��~��s3p�n$�Aa�Jը�}�� �|ۃ.4���]���F��p���#���O��;�I|X�����:�c|�)a��h��=���x!�5��b�4�?�8��0d��YW��S�WR�1y���b7qr2�W��H�����~q����z�	�{wu�1ZR�	��퓟@�{uNȈ0�K�?I}�.ÒPtG&���3$et��;>(�*��Q(:���؏8.r�?:�i�}]�<
�J��� �k�P�Ȇ�����W�ߙBՙ7��E��&:�E�F_ʚ���v�)w>���Fn�W�M�=���/��J/���"�ܶ|�&G������9�&<��
�@�����V<��m��>څ mݙ\�T�b�֒s}�����Wk�KԋH8�n~M�w��4��,Tޫ�ek%�t���\�s��N��B�g�����%H��2
�#ii�����Tx���oY�d���3�P�+6�P�w�VMU��Eő��l���:�2H�<QF���tx�<�JY�ƥӱΌ�]4�{P���W���hffL���S���(n[q[~��v���Tv�Q��u�Zvk�������#J�8��>R�
b�Ƿ�fdY(z��\�]x��;��~_Hdn`Fk6Sx11�ߘy|'g�TS'3�2�����_-���V��>�D���#b���[Fz��d��Eg+a��L���H`ُ��kZv_M0�!��Q����4ͬ���Ҭo<.B��Ϊ�"��#M�0��9L�� �Nْ��]M ��U@�M�D�B�;Τ��gGw�H���"�M\��m �ͅ�4��Qc���f��ĭ*��zj��y���(m��1.?�ә�=�;�c�E�z3���nK1�y�+�����0N}x2�e-�����T\|�)�CK|�ޤk%�9Ax 4	/�c���O�5���/:nf}y-H5�B��MKy�հ�@zxk��6�
���W����0�Q	ڑ�����B?�F�Y����+�9j��8�������Q��	�O��r��ƋnZK$]� �5��,��<���.B-?�Gj�����_ !H��{խئ�i�U2�?<gp#Z-Cբ��F��l��j���v�v�g%�i��$��R�O���)=�yI��ç>�(� ���A���U�>�vߑ�@Z�S���N�5Wv�lN��Ⱁ�հ��>�[�߸�z@^f����\S$1t\�P��W�r�r�rNhW`@�E:L��%N���]���H/�n@���%W�8�f�1�?Oa)�����F����hGÙ\ 	���}~<o�fA�y���&~�^~6�������1���.��@=�pu"�Y^��ju�X�X��z�P*k Y��ꄵ23�1f���j%�!p�(κG�Vl����,<N�'R�v�^�Fb��E��C��#�]5�F ���ٌ����%��&�hAg����*���ݶ�0xۜdP Qt��P���$f�4��kY@\��)-)|����1�Cb5� �z�HY�:�ajB���o���܄ƻ��i��2��O�{u�*lx��H ���ADTA=Ϊj`����i��F/���~�6�	�D_��<���1yC�	�o;�]Ͽ�߇��. �@�\��c�݌iD��>;I.HK����"J�Y������^�}&XR�3ڢXm��j�1G����Dmpaj뛛-xD��$��)~&�k5���]�� H�%#�4I��%���yÜ���/���3�#���.f5�i�X@��=4����\��M1�2�ՈF~���O��:zb� q���J�Yډˤ�3r��@r��f�l9��+1ʮ߉T="����k�Y�7�ص�L����1���`6o^�u�N���� ��	*�S��&g���;�?�$��(�.���3çp7m��r�0,dxC8�����1 �(�}��C�&���kQ�/V%Г ���?^}4�8�̈́3�n�A2�|,�@� 8�˘cDe��]��'*��L�ܮ�Xz��{���a\�v;-�?�
��4HΎR/���cp���Dq��hf���ɵ��)�4�<��'�G�����	$�B*��6fң�� cw%Y�;�=mh��!��D�i�Rc�e��=����% ��� b܅
�]����%<�7YLQ�q3���lP�[�6!��g%)�9�Vq!�o�3u�i�U�K����(_���l!�Ώ�j�0y�m�U�t�k�1��,7a����G�OdYDM�@})d�,E��ű���Ԅ�AF~�Ɯ�&.��􀞬 KI��|������8o�Pi����B{��٪@�թ��݌1�}���� m��+^4M��&����j���>��D��!�J/a�&1 Ü�^q5�xsF}���.��7bcz�BC�cѪ.�P!�ɓ�7saSPN�is\�~ixA.��l��(��ƕ��W1��@s]<x�j��2[��.X'b�f=�9�%�%RZ����cz�d���y��5)�X�Ǉ}"Lu]�t�z0Y�7؆g���~�WR���g�1Ҳҕ��@���~��k�^3�=��Qs;��&ύq&z���r��t�!��(��@Q]���FN&�\l���ϛ�	�_#kݐA�_yR�B�-\y�ŒDo0����	����3����k��g��ȶ-`8��%�Bt�EV��F�Ƭ�gB�qDXo�%9���< cN*#M�\�(Y�#I���R+^�7<�C�K6��m����(���O���B(��E��U��1�F`��Sn�gmɤ��M��pRߣ{������Q��j�|��%09�>��L�C�:�I��pN�|�l��}(;�ڎ\��������n��������#�8 y&��߱�cD��ͦ�r� [�p��/�dq�¦�Qգ� f�a�%�v.�����,��0����>R֏��Sy���N�d��H��Gr�x���e@݌�����A9:��ze���H���M��K���)���U��
}�o~�	c�C�/��<D\�n��3��ltr�����ѓ%�Zc��.'s^��I^�0���pq�3��Y�uU?Ec�<#�	�"z�48N����[dg���=��l�)ڭ����R��g�d��F��T�n��W)�f��ƄɆ��[�F�Z��=B<��&�G�£���r
�}~}��{l"����f?C�zK?��q�.t- ��QY,2��g6}Ov&ޅ��_� �-�����Dt/�¸{1�/�ErǧI�%�Fz6/!$�3˕Ĳmz��������l�u�Z�YQx�{ګr`��ٌ,��@�(��j�����~j�ǽ�ĸϸ��Qo�D}m���z�n�S0���,��|���O�
��q=X��U��4"u�e͜L�I� d�~�Y�W�'�5����=A��eolJ'��:QJ�U����B'���~XR2�ͣ�w�#�6�jL6i�O�N��$���P��Z�������Wv���"$oX�ιs�O�Tuaz)$��K�]���v��U���J-���'p��z�W�Z�����gS��㇘�
�P�T��?�	��������Jj�3������Xs,���8/e6`��쭥�6��U�����՟[k�6�~h���rٔ�K9c�p �.����,_-y{�|Oc�\-" =57�-ll��] �E&����s��
plG�i,!����|�9C��}!y�9O�����gO桬H%��>NQ�Ŋ{��He���Ǎf�$��s�	+�+��Wi���o4����6y��E�Gtm���П���m��?����^��q�6�g;�D�d��i
�RN����wG9c���Щ��@�UN�ˢ��1 #ٍ�P�k�g׍�b�xp��n%]�ZY���B4���0�íRO%�>�W���oxi�E�ۗ�_SGu^�l����s(���7ʥ,�[�#f9X89$~�*�6�
���+6L%��sԕ����1~d|;^��o1<s7n ��I��"l,\}.�X^hG����Ց�� |R�7�ͩ��36�ஓB�����9-ē+��gL�)�2m@H9�*�zq�����UK1
�+�-\�����#���䖕�;��88�?x�m}Kg������t͹���S�Y6���?���ۿLl.�>��˳��nN��Zp =�� ��@��5
33֧59��e��7wz��|��ٽ=-	��Q�\� T����m���7}Iũ�@��x�K�����_)�����cR4".�2!#!�i; �s���oj��b68qT�ϟ,��9E���PC:���$-�|p����?�a=|Ez%�ٻI�>��G�u/��[��J�X�+�-�{�4���｣@���V��3�������9��"�������s�(��h߬�O������;}���E�?�BLMz�xؔ�)��7�|��)M��>a�Լ�`�fl[=c���\Zz�=��R����Y.�׻���=
"K���� �\c�O�/���܀au�ԼS{��`�*������Z����|������5\��$��Y�@��������󼿕����o��Q-�t����PXT�>��jBjV��Nd�
R��*p+U!�v��m`��c���h���{c��:��tt�{��į�z=؁�zP�j���%�䏅��mΘ��1��r����7�Uv��Qծ�fT(
Gn��త[�nR��e�D˧$G��4ڝ�Vq?t�a��$p�_u��s�S�]/��m��x$�f7�5R{���a��QE�!Inr;��K�jF$ ����<u�KtdD8�>巍���i����<S�Z���-CM���C$e"��(�ί}����.нO�8��N_�E� ���՚��|5�ˈ�b�ș��~�YP�g]��<�S�� 6Q��@7�����O��1(����{��o5�LR�MI�6��g�2����J΋�v�9"����S�߹�$�F3�����i�'>6>/�ϷG$v�����!<��<UD���-�l��^y O,.�4V9<�1p��P�h�hs�SO���w��481?_�\l��,��l�������D�v�]�Z��?���kX��J<'�{b�EC#�V���vd��e�s7��[����~����B+�'Zf�.`7�`�BJ����.V��j�B��JT�:��D�\Y��(_/�q�`g��@��]��*�������ߣ@{�����������Ξ��ڠ�iUڬ�ص�2��|~s�� $�nߵ�Z�Y*
�/�RJ?�Wr\��d�)���e��af���0��lV��rq��wq�A_zH�q:u���y��'�UӒZ�v�XYb&��^��;g�Y��;��vVe&@r�[�% �Sꧾ���65�mTg�TsP/~g~7r�u��v����A,>/�(��T�vd׈fn(�V3������Z��CC��Gw�/����I:�����s��K��0��oɃ�zu�o�4��T^B��\�tn��~V�Ҽ�B���s?���Clr�M9zɍ�vΠ�?�2+�HG��m8�����i7&�c��̗�"C�`6�J9	��X�@��s�C�n��c�`�97��8�0�WW�������tXbJE��ih�+�ya	w.G,}8O���g�� }S��U�b$<�V���؃0D��7�]��#��`��޷[:V�}�x�K�S��S�(�XR1?�������W�^�_VSHK`z�
Y�����I���P��Lt�E
:ؖ�A��f���a�y׹y��գ>�����&��1�y;�P����?d���H�� w�~�h�%������x7���^btl�o+�X����˲6���§� Z���}��=���@��������	�@�;4�h�1fH@�W�23��K}�)���B��_����ݘ������\�v��:�:��1�C]\8Z�5�]��t(�I���t���h�<��kD���� {&�t����	�2�9q��`@� �r��y�g^��Z*s�᫥9xL��'��8��i��E�_e�6q�p�5D\Ywߘ�DA�̘]����4�a�[���ܛ�BE�����.��'7Q�$�L�)�˒���A��ʘੂ���ͼH�"�����lhI�b��tد ���u���.��Tu ��=��e��3�g��Cˤ�ĺ�ᔇ��3���A���Nx!��x/0?�:=h��Ǔx7/��L����u�0�5�.W����5�L"5�R�[�|K0k��&�O�
U,c�4����iM����]]��m�۠[������714Dsfb�����eb��[�A�*\,q%{%Xq�����o�E-X/��q�1*Q_Y�#��^|�tq0��X��u���Px�A��y���/�|M���8��*g���ܓ�Z��;|����J�0e5O��{~]�b��b�Yx2gxq?Y�� `m��o��²[�q�\4I��,AՋ�u�G�1,3I���H�!��6B )���L��[d�Z��,b����Ȥ��Չλث��^��h�Ld�W(���~�.�X|;�Q;t:O���z�<`�w����:�M;��M��ͼZ��/��g�Cl�B���mC�*������و	DeR�w�(���s"�zb<R�4z1��I�7'�������'%�h؋��}үcj�/r�uf����ɲ�G�de�F��)
$��X��a�BTY�,��_�O�;��DiԤ���"��L��_=2�tr�\��������9{>>#}^��gΥNo�ù��B����Ɯ���EC|0���f�\�}�2�����SŁ1[	+mS�z�`-NP����@=�FC��eR�[d���E|[<W|~�M~�p�������c�2��wب�r�8`R읃�?�� ���{����B\.���E(xwl�Oע$:�ty/��!�B�������J6�w__{���ܟ�(�4�r�� �!�k�&x���-+�M���H)�\����Y�O��B�mw��{��� ;�!)lq���YП� �ȇq?��#�ٗ���jU����t��s}�O��P�������3OSed�6~?�9G�2F��	���a�����ZAyilT�<wb����d�k033)���w�/j��V��#��<����"ψ��$I�l��ˠq�-z��w�'��i2�������V]qȫ��7��v_	J�]��
��o�ʎ���z�s� Dh�Z�"�i9�ԍ���>�ge �s��6�E(_��Ha��+���N�l��bX���9a�>�am�d�c���]\^�B$1�8�k��֨��_����B��gSi�U��A=Om�Z=�A��%s�@��6Fe����:�F��>��D"��Ho�W�/��#[C*�/򷱔�#.���B���|��3%�S y�o��y9�|[�5;;p�v� 5#T��m�Y~�I��򃘴z,5�t�Pn�d���`�&�!0ɮ)��@гp��]��t���}��X�8ńu�MI`��8������"�,����b�)��0K}$�hM�w�2R~��9z���O���5�w[:cv�M�A�HꚀŌ���y�!�Z���_��p��w��rる�vv/4V��G+�|��F�W��)3Bt�豄�Q֦'�� �������" fѨ��y�-U�f���1�*�Č�b��  #`�Af�!�e������5���/G�=zVE�x�K�� �U[��FP��D�A�c�4�C$���J�B����6��o_鏼��챲�J�:��ۙ���u�)X����F���Oi\��Rސ�)�gLj��#�ܓH��U��S*J=��Ղ¹Qy���D���*����R��Dp�P�,!,Vb&ݍx/�:k�XG{c:�Z7o;H8_�T�ah@ƙ�?�~�[�� �� eK������� ���Ѕ^�9-��"dp:_��b_&
=���N���*��^��\����i��$����.yܧO� �k�!�ϸp����Rjh?A�1n�0��Y������%J��S�/��%�a�k����tȬ8D��Wh����h��ugǜ�T�õ�J_[~j�7���	�"ԏ9�:{C7���D����Ȧ���8?.��M`E/���e��I�����I�����U��Q��amb�ԕH;&wG%�P�
�,�
���h<-���p�4���k���T�F�K�H��b^f<�m9���Vk��M%�o��^����� �9�l����j����)$�*u4@5u�+�'�M�΅#[�?y���ח��]}v+]H �U�L�=��L����3�2���M
��NhUOb��J�˽�aۃ��9%�ː�����_OѠ��T)in�yj�.�}j�h��ι21]�Qh�a���;ʦ��(��-������..���5����bwV&Ď2��RZ*C���Й-$������7���a0H����'sk��F��-�p�&�ε�q9���x��p������I�_��2�\�����0�U��ho��h�*h��Zb��*��9�����������oz͡3�c(���*ze�&�q֧�Zv��7�l��ĳQO�7w�VO��=i��]�X�4�J��2�WԳ#n��j�K��!V5C|١�u���܃i�F�����vO<d�m��%�@��D��=k��t0}(�
N��,}�R�
R�r'B=Feڷ�����XG%����_��������|ONAT�7`�g���G4m��� ��oeM��G���^/b&�"̛��{�wf��;���*&ǋ�Ma;PU^a��篥M��b�%/��p�jE�e-�<�&�`�@�#N��O@�x{���D��/�d8�nToM�Z�1-��Sf��8��У�Pi�ɬM�7Si�I5�:�d}g@�V%x�/����ߵE�Kd8F3i���L"��z�;�&'\VI9"9���Е�����n�����+��I$��p �p�8[y d'��:�}��*��<+���
_r>$(|{��/�'N3�%�R�	�����lǩ�U��h~�x��o��-{�w�K���K�!)o�;Y\�d��Y��ٚ?5�����1�\��\��"2�G������L��v����ׅ�!��X.O�9 Sw�.��č̘-��幝 ?`�J���C���(�0b6�d���L��̼��6��y0ho�)]t�өF)�(���p�MS��G��\c7K>7�c��9�*0hoEe��*Q0�u�yj�9�ա��1):���L��E��v��Bk���eK���l� ���ȿ��ϱm"�Ѧ<o�(lW�)[��\y%���য়1'#iB`3��jO��z|@��6e&���z<��w���`�
Zt�5E?*pq�5W��ge��c�6\��p$�h��ɇ�e���}���UaFp~�l����R#\��G/ʒu��;1뉤=F,5y2�w.�|�}v�!FE8+�0��Cg	Y�����3�{��؞��On��y�<��v�OU�
�q�d�dn��tr�
a=��-z� U�v�7��㽽E�Bkh����X��R�l3f:�j�颵p>�0���pC5T���WX��l!8������K�/!�0�8�h�}��%�Y�7�U;Y�h *Fj�r!��քI�5���o7;��o���"�|��Fa��@pYyGv�#���Y`�֤슡LR�B��� ���u�^�D6����q���I�g)�}]p���+�c2'���QL�n�Gצ�8���[�H	�ԇ[
���ޘ�����<z݆'����#~�DO�W\��:���0��w�$TV��Ē��C�?4��Lk��%B�1�dx]C�)��T�0��WGs|扷��F]�]� @9����g�ړ���o�P����f�D��m�-q�re�.@�Ѡk ��x}��i�z����+)���u���/\�V�����j�[��!b8�6r��{Mm-��$�����z�<�L���i%�O�61B���7v;�2֍
w�� ��aL%׃I������[RW2�a����6�O��ш��h0������At-�vn<M�aP�v�� k��M������He&u/�E6{���>�߃�S���%���T�0$���T��>&����W��Q�+\�"WS@>�;a~�[���y�FV��o�z rJʼ�_�?��ኁq�%p�/|V�k�M�����e���F��ߜ
�	�#),)%Ù��Jr���77���e�/�O[X���0�5b^����C�NI	� �\������K5p99����z2Wa�^���i����Q�O�I&�����OX�PgQڵjɏ�GYg�G���\R�g��f�/A
a'��o�ﰤ�0���-���{�Ɵ�c�׺���U-�L;c3�{���I����B�7tn��w�121�6A��l�<?�U%�(wi�Bv��P�
Ӗ34��Y�*�/U4�\�o^)r�v*��4�@b�i�'A+�����ʅgRHvЙ�(Ѐv���s�T���`!��cd��d�	����[���������\���b�bCa��Xؕ�5/Ո=]%�9���� t��֥��y�p�ڣ���=5�;0�?t��@�&}�]�`��w���p�P�p�SGm��ZQ/�.6��vO�K0�P���I:��f���7���w�\��=9Q���ܟ�b�n6^�SX H�;����n��.>B4]E�(���8���(Qs3qB�v$�1�{�8��͔?X�W]�8������c��S�������2>�˹m@_���G)��W%����@K{h�z�":��ϻ�z�xm5x���[�;�a��b�|�>b5D�,�x�i��_x�$T.�	�H>���|r��/BaxP�`�_҆�_�A���~K�-�N��wJ�;��mFU�T_��%�=�̎(M�Pb�p!�8�뽝7�� �h����Ґ���T6��;~�c�},]E���q��3K�c��|W�����el��Y��2��ᐕ�)Y}�4���5}����t�*����>J�g@�DS���
��Ϲ��׮,B�6!Υ��I,���9��F�W�����+jL�b�C��E�>�8��D��k}�ul�7x�EcǰZ���ûo�g���*\Ҭ�"��l+H+�3��0�t0�����Ԗꊭ���WM:�+1���69Q��\�$֛���V(�?Ns�n�Q�{;Ia�`h*l~bM?�s㡄,���g�ΰ1P�\�'x�HB��Ʋ=����Ò�:��o���36�k�y
�-Z�.����S˅gя�\q�kTD��	���q]������_Q�PO�?G��wכ�	�戃+7�4�q���W����)�C �^1�
؞�[4��q���D�R�ƻvᾢǥ�|����j ;G��
/��B��'ۜ�.�c�@ ��8Ay%�K��ms'�L_���rQ��WS��p�C50�g=Ɲ,�b����mZ����v
=���	����~й�T�2(�K���{Q���>=j}t��@1 Y�t�i�\�МYr-�G'Xl��4�A)ҝ+�	�`�»<���g��t� �����ɍ➋�v����P������5Р'f��b�#�p�dgΕ�Y�|m����M˾vC�弚#�	6z�7u�����P�� DF���+�7���x��1���Z\�c��h�D�`���� !aM�֮��:*ڎ�ehDT.�l�������Br��)�M�-�\}ۅ�rm��5����_�u+a�jvZ��rP�� �.!؉����Za�
�YX.�7q_M?��(e�}����N��<�6 *û��H.�L�s��
#L7�G}Q�!�+)1�OX�F%���k��:��6	 �~hj��oL�f�����7�i�R0S�^j�;��r7��۲S��}=5i�	�2)��~����̹�GtB�Z�EH��6_�t��UN:6 ��5�_����[*�c���>�*,[�ל;AV ��"{B����o�f=]a���"��,+��NP0.z�R�f�#���`�"���e"G�{~���)\�}9հA%�Ɩ���J�N�����m+�VA]a�����Ûk�����'�]1� |�.-�[��p��?g�Έ~+ �6n��.�:�[��Jd<����垐�S���e�{�J�lqT)��,�@�@b��IS�,�P�� ����z7*%0^>2��Y���@�m]��ܛC��`�XV���%ƽ#=[�S1��"k*e����p�Nd�w HuV2�,�$t�D��߀�~#?3�W�p��4/$��6�G�"�}{��GK�C�Dn�����ߔU@�N�4cH<]���&j?�~��}{o�?̀�5����^�q&��������t�hh����t]�� BQ~�xuF���(s1��"Sūr��(��w�,Q��Y����$��W܁CJ�A�X)���ќI��Z��8�˶���/�#���Y�%o��$-�#\a�9@d8����w���p�je�+〭ʩ���f���8�(�f2���gV�����2,��e*1Z^��m�s)��Ҫ.uu5�f�f$��N�μ���0�G̦�<#��o�JgVϰsѢm~8Bt�y���)�ص��A��n'+�dY�

�/F��TW"oc���O��g���p�۬�<�z��� �r�38�Ȫg��6~/��O@DI
�2��#�D�����k3FK��m�b�"Q��N*V�%^�� ��5	�Y�L��,�F%����E<mvH�KO�~�9�B��ph�i��d�>v��)���MM �?���^���*��P��:�M�R ����Q�ge"�=�G���Y9�z�Q�Щ�V��0���y���E5=�8:������В�g����ޑc;Ha��x��4^q�� ���	�T�P���_�e?Y�J�ҟ+&A��M
l�:�Bj��V҄�"��)�ݱ�;�]��^=�01%����/�zu��O�f_��6 �����B[t��U|k]��rh�D榲Jw�#{p��6}Zp
N�������Qg��^q�GM�C�� �e��w �#��u����=oD3a��il?��=|���yc��I+>B��̠Z�\u����<��L�41�� !������Y�[=\�!`N�쯲4��"u�K?��)�u����d��ҋθ�%*�x�o�<W�Azm�`�d����c�'JsE��1��#r-l����7U��iIvJ�$,�.�A��.�jB\�T%hUy�H��Ui�����>�����Z�)|^h�6ll�Ԁq���*�.��rj�_���a��-�A�%�!��HZҫ'T���B�x��@9*9Y�3�(���j���-�*&}r�)�V m��P����W��d�75��}��֬o����>���X>�9%la��\�V6C1��B0�|=�P�+�0���V����]؛���4fG�h�b��c��y���׻��4�&��n� ��/�h���`W��:�@%L�87QZ��s+��N�2C�j�{K��^�}��y�"�B �"y��˪��@��X��UV�]?.���)c�(�Rs[�8z��QN/�s����Iu�QP�dS�-J�c+���5' �d��ũZ,�L���q�L�V\kv�|E��tO�If�Iȵs�9JR;7ِ����N�Z��ݏ��� �H�Y�r��S� �Ī 	�y1h�j����dg�m����� ����j�[�Y&ę�!���~�]{U_��k� �ז\�!$��ȵa\�5�� f*}�!&�
����m+F{���3E��:FeF�P"�0XK�'z~
���@Jda�,�����5:�#��,���u�3-��,=;
�BGb����Yթ
�f��H�NÎ�7�=����<�	¾K ��2H,m?�P"�I-���@���3���	��	�.G��G�>�|_�^�1���)�x|����P�=�D�o.��^��(�dp�`�	8�����2�]-,jE�f��u������e6ќsu�X�њ|өs�rdg'0���U*�+1��c�o%�]�N=;�:�Nd;��{\�?�H� � ,$PZ��R){҅\xO��!�M����UƓ����S�u�
IKoW��J�{�Oa�ɗk|5����x �F�+m�<�3���ڼ
Ⱦ��� �iK��.���	��`E� :1�r�{"R�E�O���d�E&��u��5�����Q�"�����q<�'mfb�s��p�vtr[������e���r[�^��� Ϋ��Q(a�$x�ys�s�y���TXh���ެb��P�>����af]v 9�y*��Z�ҷ"Wq��+W4�B�b:�.znh��=�I�M�uʹ�'����n�^�Ìf����\���>pʥ�U� ����!�t��!Q#��S���3�� Q�&���LDI~Jc��B��/
2���w���w[�=B@�yj�ѽ������|��C�G�|r�V�r�ĳX�������dFh�5���YI{9&5�I��N����hv��d����U��	�����
�ܛ�K�
^L��E���M�"i/��cz}�;Y�������H4�����[H�rW�um���l�������;i�[n-�C+JᤓŹ�dH��f.��[�����-�X)�\�H+���������s�N&�X!������꣣��M[�/u/�j_�h �����L9u�zSH�F�]�n%fsm�	���8�_#�p��o1��d���ng�����iRЮ�F���C�3� 6@�h�^��w���ǉdK��"G��A�G���z�	�Uk��,v9�K��}1�&����#3�7�aeQ<(2�{z`.&6��y���2�=2.G^b>S�,�C{f���Ϟ"Z
��!B��<q��z�{! �i�a��qsc��t֑߬ ��5p�U��x*�����3�z����P%`�e��Rx�l0mR'�q���&��7�}*���W�Ѩ�9�^I �&�>���>�����д��wϳL+Tr���s����v��������.?iq��=��.�{�MIl[��\�Ax�1�[%���t��'W�/��|q͑�/5T��y�83�׿���]A"�q����/�K�5G𙉈�:��@b����*�T�Y�Aq����]`(��� �^&ޠmX5U4�q�a��W�{��v�����5(�sn�L���'�}ѵ �3d�,�w8o�� ���*��Γj��B�]Y�w��4���wt�y:�$FN��;�#�6{;�D�n��eѣ����K`�	���29������@��Ya|yH�^{�8ݩkU|�j��5�����=p��^�O��<^1֫��࢔A"8|�yMf��G@�����i�u�9�ǖ�'����[!6���:>I/�]k�L�o|��i�6�%�V���;��+��Je��ݫ]�E�*Ч��Ѳ_����,��E6j��:�\�_�[���V.³*��-����Vof�9�Ƥ�� ���.��]�]d;��m߶Nz�M(�R|:;�:-5�,����cq:
x���D�tx��Ћ��W˕a��a.�����/��-~���qt�:��i>�d 1���e^�>+�Kʝ�˯Ԏ/���LB(�T�v&ѵ�H4�ݸ �B�H�,�E�2x!��9Z��u��(�B�e�'w؋��?��M��O�^�kN�~T=Tɤ r����J������+�	w�NL6�P�#��f=������[cu��%���U�$&F�X5V��3k�w>�U�b&�ł�@�,�%2�%f�ዾ���֓�!ad�ߌ�x*`�U��S�R��_���U�T7^���	����ſ�)�TZ�$j�Y�d�XKMлF�ܤ��+�xg��;QIa�}U\�����P%��P�o#�w(�ôw�S�i'����u����k�\>��'͒��ϯ�`����00JMX����hV���}�uŻa�m�c�.�;�6�.��r�Jp��`��G	5;�����-v�'n�$nal���GP��{\8m���yq��Q�r�򫞐^�����E��_I�ט {�b
U�:x�$m�C��R�Uܲ�9���I�Br���t��@Ï(m���/���!������-����y\.B�d�_I��(�������8��
�Z�$�T�*�?w�G*����Q�:S��	9�R�r�A����&E�2��Ѣ���[jM]�Q������^+_ʨ^�Z�sJ��A�?��`�FF*w�q]���� НJaC ��|GcL�o3r�W�f(B#w�����Ao0v��ڃL���A��%��� L�e��<�o����J��|����X�dK"?���b�D[p����_�^Cf�7V7]OK&���h˟�������8*�����t)�{�O����~~%���0K��	���
�6���7��oi8�0O��xoa%x�t��iGm:ޡT���I�geݔb$������[@�BՁ��1s�|��9@��y\�����n+�(C@ŷ+��"�"��\��XK�w�`��*d����Z�7��ban�=�ֹ��ʿ^Gn񁐎��-U1x�#�~��+�0�y)іDja���v�j'���r����z��1hG5;[4yG��>O�ZB?���(K-	x�	ܓ<��Z6f`;�	�3&]DL�d�e8�O���W�1`5�s� ��JN��y!�.p<)�6O���Ez�!h9��2���G������Ѵ6���9 5�ɮ+~����Ϭ���������<уln��Vpp�2���p�,cI3�h"�]'�4���IOv	�w�c85�n��=<W�3�Me��z{tG&=A_�.����� ���'$��H_��i���ȝ!���td��N�1\�����:�=���ޟ!���V��W$%Mt?6�-���ܿ�v�xJ�ڳo����਑Ey#**j��]��f�"�=��x,�7����eqjH�"XY�{�C/�ȿ͈ ���}x�f"4�'�G���1Fχ�6dR�6��NZ�Yi��c�Q����
�Y��$�r�|k\7>���I�L��*�����O�B��|sGՍ�N'i���]��
��u�`��i�H�3�I�܀��9F�Y7��'H�]&M���*�&�4�b��(=���������h��]����Y�[�,�F9�2#rӮ�n���jԺ� .fV�@�Eu��]�(�xx���
ϔ���u�2X%:��$��ҟN��D�S!�}���.�u�%��u�,�]ƶ�uئl�:�ԏ�>ۊf�I��wy2�F#Ti�ux�2)�`rA3^�n�HW�\x���&2��K����ޖ�%q釃���qPS��tYQ���M|J�����uSm���ht����FRG�Nl��<�/���=�9j���}؞�a���^86��c�;�Gv�k<t��H*dv!�ת�(ݪq����#�hn����6���x.�Ǆu�������Ã1�y��|���=����g���LM
:�t�`� ��k^���b���O�������b8'q�b�����m2�j��+ ������Ӣ+�7�@'��|�d�9 gm��w��9�&��pT�?&]�7�-�N�cf��A�51�yw��2P$��Dú]����J�R�p{�Y���-�W�q�@�	�m�,Trd	(^K�fz��Pp�k�C���j��kV,s�9!h�*NڣCq���M�q�<�}����p����T��6��"E*������6���G8��4D~u�[qsE&Z�Oq�T+F�H���̬)��pl��.������=���T�����e/g;�B*֒��i\*~�8T�[�"�Z[{�r �&/L<p!�W�q�L|�@XƧo�u1�Ox��&��g��5�Ew���T^CW��e�S�H�����hT(n���>����9R=�c\9�)�58��&�cJ�ON�S��H�|$Jqd��f���[�B��V����k&���Бy,G��� ��SI��=�GE�&���|1e��e��'�7�}4I��oV�m����V`�����L���wlE�����+��XA6���L �80ԓ?Mݙ�V&.���l0<�G���8�r����xv��-�3��\�c�O�D^�!�&�[_�Q��P4�%j�'��%��`�v��g%@Bq��@Ji�	$a�:@s�4{RS��d�~�����ÖD�b7�2u�0%im�i��V�󋈤�xy�ڤ�_�%�3��v�4u@�ez� ��r0�>�d�A!(o\��I:y��m�9gj�a5P���J�C>�6��q�Z0Lƈ ���-|޿�@5���.��j�goΪ��ț�m�?y�x�AZȶ :Z�,�G�}P�8���j�U�*�sX�B�p��%G7��G�:e���Q�i:R��I�-A����|�C��T2b_�	�%H:��~Z��"��; h�*��>���sj�jyq��a�	�f҆�;&~� %o-ZcL!�,n(�W�=��V:��|�a(�R_t&����@@w����/ �%J=���|a\J�%�6P�Ym����tF��$�L$u�g���:�Q%�1S"����� ���X�a���8���X�V琢�q��7��I�r8�ÁC��> S"2��N�F����dĨ���OI�ƕ+w^�Q���6@��C�p$�EY�e���y�K[>�6��C���
��g;ך�\K(C��G�D2ev�]��������Ըd���
2ɹH�-��y�vd�O���Df*.�:�^�Ss٤j����z&I�Q�U���bB��:J�H%H�4�?'�,�QN�Ш�iy�e��|.���Ԍ�S��D������BFf3�f��	�*���i��'�!{�$��p{{FϮ+�Z6b�=��%,������>T��0E����lKOJXG���mqD�Q��k�����Z���U[���^���C}�睫���V��4@��P�d��}��Y����k�h�/���Y;�<�ָ������LO��8������|f���3�McFw�31��F4�4Ã��կ�8�m6�{�	E%F&wh��T��n��S��x�'�T����^�+�yPmz&��p"_���t����A��a6�q�,�x�cnҧ�%��}fl~)��W �5�U����.['���?l�����Sr�ɿ�Q*�c�g���v��~���[�K�q��s�5��pIU��x��瀹ϏsX�1�E9��c�{�'�M}��#���Z-���4�s\�H��`�:lI_����I���7+T�� @�H_>�����u����MK�#���I8�.���ʮ�Y03Y,v*$�ϭ�=
K*M��֒�����B�R������-��۝u�Q�2 �%$l5�<e�xR���V���]_e��6Fh��c�ZT��N�ń2ڛ�1Aq���=3���������Sȭ���!d��o2Q��ԱX?��pl�^�+�>zb�`SA�x���v9Yؤ�������tF��K�%C9��C��-#o�&H�j�+���Ρ��d��ґ��Y]�dW�L|1��yr/�hpq(����w7Ǩņ�޻��oq����T����|�����ŏ��Z�e]T�F3����G���Y�zr.�DI��+�5{��U�@�eӧ���Gӌ�9G�pm�׏�`3g�\����F��v���[M�7��ũw�u_�E<Ȍ������6�*�O~$)�Rh.��z��0+�d��l���y���`�	Ҏ}����)���� ���4B��ve�߈��hA�'���l��x<,���q�}���u.X^3��~�%V���:gE�N|���GBc�ȥ4Y���L��u
�2�X�d�] ��1�ޤ\\u;k�ҍ8jY�z>E#���V�H�o
�cdִ0��Y�ꏊa����Br@�ޔc�br1ꨊYJq�cI�/���ȡ�~��0M;����$B�����`(���ĕ� C�i�7O������#��Ɛ!�$�־����g2�@�c���"3���i�;��$Uͬ=#����e	%��>t��Qx.GM�;h��G�RC��a��������o^X<�9�3�I�n�1�9���[
���8"�]=���Z���%���v��I7�3P�|���3�ob1«�E����-���Z�΀��L�N��u�ZB��`����z]hK� ���Nxז��s�q�Ώ� �u@~��N	؁��� to�������)hg7In�Z�}\^�����m�ݠm�]m���$�=s����S6��3�����t'�H���3��\R%�	����jћ� $tr� �Y���o�*$^+��-A�6G�~���VO��B��"#ܘ
��[�U4�p�"ķ�f%^Zd��&+<��z�k� ���P��Y���e���#�Z8c�܊�[�<`���f21��*أ�k��HfE����9��f�KFi��R���L T`BG;��I�y�eO��yG{+k�Z]ę�~�V�9x>��"�Q�[o *+���A��6:�s�B,Rd����bį�ܒ�~�e���\��7��3�V�$���é]y��H���F��Px�CU���Ɂ~߄�������,��Нa-�r� ü�ykܿʭ��v���?�M�s����2O�A}d�� � ���#7���hb�㥙'�n�h�}��*�������{��� ��%��1=�>����jR���ek\Yf�g�{M`O�TiLx�m�}mW)�bk�8jtH�Em4R�-7;�8?8��]�iPx����|1������^��SBP�]�h}�l��	ve��	j��)��Rk��FS�n�|+s�=ٙ��gC҂��ݭ��eƲ ��~>::�Q��g##��O���8o�S��ě�s,�ʎ
��7/��K���7}	
|�+f���r,�.u����gu{,-�Hܛ� ���*�	:�1�9Rix'T�p/݆d����7�v�,�A������D-�#�4�e�Ag��:9�S��+0�?:�߀W)@�I	�2��$g��!D*�Li�*��<
����d~=.m����S���}!��Ypp�+ �� o
5
���:��$��Z����,��/����^�8/���T�U���=is�_{Tt��T!3��?��=�Q1wH�tw�����O8��a(Q���llC�����I�-��	NH�N{�����8��u�@e֜}�2)���ng����&T;LMrZ"g-I�;�j$fV_��J+75��>b;�1(a�#�_�$�K!�)��ݠ
,-Z�mGth�i��/nv��)��64��e��XP����+�0W�?���xUYd˯�QA�ș�T�/���t��8�[V66�\ͬ�� ��8�� �6�
YN�>:>x�߲8Ɛ��|�.��ֺ�=̗Gp�~ƾq8�����~&�Hw���[�� ��f�Pp��1���
����_�qH{�*�A�n+
�:0����o�m.=^SӍޣ�gcOB{�kw��'��;�k�2���#��?9
 �ۥ��t�vID�`��B�w�F��Vy�����4]�z�Mؒ���B����qbZЈs�xGK�Yr/�߁d�H�_}S�C�P9d��3��*��Öh����{<��R��!0�w�(U"�N?���$	$Sh9�\3F�"�!l���d��b���k>@_�x}�/���A�ɘJ[��1=]��2�ak�d�9J���p)�ADg�����1���]|����d�l�IڝSj�l�����2_��ͣ�=%`/�wB2�k�[tܮ����Y�vv�n���1C���e�o���Bv�?�;��� I6d�MjN�;�d9�I7���[Olθ\q/�N������(��{�*�O�
E���A��h��iL�kE�����74`OC�6Q���w j���-�&CL/�\��a<�|A+;�C�E��6C��_�]�&�L�ek��@�L�vs��k��zY�9_��d�%8�O�6��� ��Es%�.�q��6�s��*뇃vی�ĉ7�I�ÃpNM��G�r�K�ÏlE����S�AM�>���O���N ��
��tg��Ʒ2 @n����1w���l��/B���n��������V��sN'6'�Cd�Y��
ր�{�M%�i�8|]�<A�bX�fu�-��"ȍO�����m� ����2U����mE��E;[˼�A�C�bm�Ƀ�i���ۺT�%H��G���f��}�_����*W�[�b��4���3_R��Wj��+ڔ�*�G�yH4l5�W u�����er0H֖?S���]\�]�Vڱ�����'�DĒ�	����?H?�a-�K:J\k�Up.�K iXE0c�����pŦ?��+J��V+	2t�B-Qx�����P��'�0�s̟\�Ǐ�3R`	%�g��fkP,�9֡�Bx�I��Hq�~V��q[��t��G�X`����${K�D��ـ&�Ì�����R�sx/�|�;/Ś�|���/�fj�P�����d0��5��X��}�d�Ovt>�Gc3�� �|p�Ƨ&��QP�� ��,���O���kh%��q��S�q+	~��	C�0�c\�a� 3�{�n ��"�������e@�� }�rMDj����9�U3Ѕk
�(�i��rR�x���dbbs\���f���#X�ĕ�+�&{R=��2,|D����Y�/?r7��]����)�q��`�mA��Q���WR�V��z��b�{I�������,����<�~Ac��h��sy��Û���<�R��}Cܚ2�{S��q�����S|)qB˞�V��N�'8roڍ!15]�D:�U���܌����R�(�����v#is�*����/����L!,z@�`�F������� �N5 � (OH�!�~�.�߃���xq�u%��D�7�e��#"�S�kP�:���nm
��)V>��0��;qq�[T�e�%���Q{#���B�.�P��P�U����|%�[KM�*�(�4��1��#�r�3�����SF���r��%�6`� �y�U�7Ly�O���gr�;1_/P��W��cr��${��1����8���A�	��ε�!@Z[ѥ�ʦ�
�o�Ig�P��m ���ȅ<���a$jh�QY��ڪ�����L���_��u���8��p�\$Mm"o�:�E�tYRa�ڈxq�y[��ЧV	�J=�Y��� o�eSf��V_Jcs~�9��*4 *غS4V%5̀O�_v8"%�x�L��/��Al�"i�x�ĸݕDK΁���8�<�Ls68L/*^EՉ^���}EǱ̘E��}{(LS3ā�O*�Bڜ\#�/���#^e���(��y����ۇ����C����r�������"R��.%�&�g�^(ǏX�lN&b>���R�0�wS���e��=2���ã`���M1^�ԤF�d�p��D\Ϝ��d��d�F�� �ho�gG���ZH�&�~.��!|�E2}��$�A�l��uC6&L��{��f%Ո�sh�Ps&<��X��96`����9q��Ej�J#�3�Pڰ�H7$7'�"��߹�=��.�
P{�>:}ym%a�"�(�,�#����0�a�La��WH���@����J�t���|R�����x����pmU�o(U��[�Aٵ���'d���f�����x&�q|���_ۄ����J<(��kf I�ҭ>.�`����k=,�00o/.V����^�7��zm0�Έŕj�r�@�^�n�������ʹ� ��`{���>Mi�O;>c�#�.�J���f�:^�����d̻�rI���j�A��𖟼�
=���vRp�=a*���Z�l'B�ݵ��3����齋)�T���NO����L����K6�줞�Jȋ�����k��ͺvs�}L��^L��瘔��p"���Ľ��a}dS<�C)���O�,�98���F��٪ޟ�;e@��K@��A�Ey��Žf�� �<r�8�`�{�!���ۼD(1Mn�_P�� �����wG�'�#�k֋��#�P0Xi�����5��mu�S� �|7*6j0�Y�����G�X�1I\!�L�S������p+�
cg�1�]�V��R�b�>�R���4Vx����J��,��S9	�*�7%s>о��Gu�sD�Xܔ�7h��zP�qb�\���*&�vti�N�JJ�p�UOc���Cp�K.޷�|J�P>.�Qx�#+���;��n{��D�wV�s) �'���±^DDȀF1��x��cd�Y� ��Cnu^�M�frN$Jr��h�\2��x��:vɞ��MD�D�z
@'���'a8k��ԓ<��)Ⲁ�+Ǧ�\a��Q��cYf�zK"�z���G�� $��{�&��2����P��+9�:�q��,��1pl��w��D�yDo���_�rO�w����bA`�@���U��n_���l�ޯ��=���.�Ư���?H�v ���^{�͘�`,q�Qi`�m�t�%��E�k�i�2P�r���J�͇̈X=t��Ș 8ʸOlX����<���?E��q^G="�4�Z��M��U\���זt,�2b�Y���\$h�y����(�a�q�l��n�t�j��`�~]R�e�k����[�%c�`�yӼ^/��x&��ꣀ��P
�F頊2�o g"�mj{�-����x���������y8����rRH~5m7�=�79��Jq������DVc2gS�/�"�����u�<�v+���>d�uI�)�!����X|�>���{�d��1˿�F�;�����K�c��ծ�K���Ӏ�y�Y��zQ�(����ci[�>�Ν�z�c���<.�F�)"�n�$��WYv���o��Bj+�����N��G�������[H����<|��f�PC*�(�پ3$y�����(��/���*�:\�Rs:g޶�fP=���	�鬅������Lj�Q[�H듧�&�	Ø����v�z�Z����2�`JU��W�2��?F�9e��
�E9K�p��{�HZ5����"=��I��s��gpb�+>�-���3a�z��ړ�ey�X�y�ύ�7Y{@��8v)�Y� ��n�'�J���]c��'*��ҍ����CN=)P���k�T*������P]�#�����J:�E��O��s��^��7�:�u�˲�I��Y/@sj��|�F��^[���4�����ÕtR�; ��ຑ#�FW��� �'+!��{��V�: ��Z���JJʦ,��Sp�����^�Y�R���$��s`�9�\�z���g"��|���*��\�`��|I/�20��p��9Ď��>�E=�:����D�~ο�Pp�X7�P�0���;6���zqpݱ����������5_��݈��
��1�_�=W��I���dp��Z�Kq�-�fRp������M-��q%C�#$������j�ja��d?�	�vY�<��=�m�dz}��T�D����6D�T���Ul��Qi@F�!�q#Z`]�{��e��6	4�����8�3� ���4�k��ԋ�`�?�M�h����� G����v��p=��bL�sl�#��J������HW�Q"��r���_u�4S�f�7c{��ufyĒ�������ga���G��J"��%z�7ꕉp�;-�h;C��5�a�\��W�e@��I���w�MB�g��8�*D���Q9hm��m�X��7E>�]��"}��q��w��5�}R�s�7`!DGgeHM���΁pOTH�����Q�H���]��u�	�u��Ou�hp�v��s�������9G�B@���ogaU?�&��<�O���r�G��캊�����>ƪ��+�\�D�4�m.�ȿ��qx|�.��hZKyQ������8���xƴ��PI�lL�A��zM��,�]L/9@�*�e�/�%5��C��t��(L�}�Jy�zi��hr�h��3D+�6�y�IK[�Ԛ��i'D�W���}f<ضҁlՂ�$�:��	ۣY����7�T�R��O���*���c ��lO`:$��솷��\��f�_��ӈ�#)�ae6M�Rp���u�áie"�zvSaG�Q�P
�;��P�P��N�cO����m����7���>�A�D�n��3�>)>4$��!�/�#����8X��#���L�V*7��3}��h�?���]'�h������ha{Qh�",�$FL�-���`�M��M�������M�7r���������V�>�@��uT��w�y�R6�%�4�0XT��Ih��X�pi�5l:ɗ�,f���r�]�{%_N�e�b�j��D�D*3Zm�rB� ���ʷ�񔠂��-#L���nV��z��	ESq�K�
��}���.Â��ܯA�� �&E��Ύ�C�\f�^38�6�@�q�܉]n�<B���Ԧ^D�G9%�;[7~�96 ^=���M�վ��\z�D��~�-�X��`|���S�*�M_������M����-��" � �_�Y�|��)��[��H�N"�:��k�-�a4k����ɪ��e���%~|g�]�Ds��0��=�+z@��D3u��Ԯ҆L>x��� ǆ6�J�Y�ґ����I��s��b��KdG����`����c,��O!��z'R����m�?��G�(��Y*���z� �����r�_�t��A����E7+�� ��Tv�b]ˍ�����7ާ�1ua�}����v�ɔɇ0������4i��D0}W3Χ�pCo�s����u)�e��"�N�����@�csҒ'��>p^G<+	u�2�[IW�l����h|��� �r��X"�������J�~I1trF$BP'6�Zf�r�vS�a�aJ�e�={���g����^vhl� �U��c�|�H�J�" ��L=�q��g,>�� 4�b[ol��.��d'�;S��sH��Q�d`8^�^�t/���O���n#��� �T�[NX�7���s+j�ý��}�������ܡ��!�/��)+�=
��!u��l�8j6Ah��e�G��d�8%�٭��]�}d.�Y�8O~���d#�N�}`wQ��TE�����.o\U|^̌v"���@�V��I�i�C�ڞ¿������q�)jc&U���L��=���@0����T��5��;�>�%"�2�¨&(��T�l�`��JQDm�S+tA]!{,	ypȒu՚��2ґ�cb��M�^�����s[0b���k?�;�n9����/���n`9���BU�L��e�"��ڲ�.̠���C�$��B������`�u�9mPU ��� ���$̀������9�h����f�>R=_�$�kSM%�L	`����	�g<�j��~+~�_G�����q�'�m����q:¿k��������@� ��ͺ^��g�!��*��������+�iLy�h8��l��0���ڼ����s�!K5���	?�[ƺ�'��7a>FN�8��{��c���RSλ�y�fuD`lh�N��5��f���X
Ec]��~��s 1����s}��[/��D饻�D7Xʳa���Uaڦ��=j�NB��|���c|?֚���gP����E���}��ԏ����.O�8�4��%G���~'�Ӆ$J�ڜ[����
��|��+��F��#B���Q~P���F7��S��s���ܬ�PCW`�419`$I�~�&�G�-`�X\����(��Ϫ�b��Z�� ���5
d!\a��,��pM��dr����h���tQ��b�]�3v�iHHIo���eL+�d>���X���;Ie]� ���4���J���������
݌o�ޏF�����T�f��+��)׿��&�tAЏ�y@lr�*Hr~A�6���7aƱ�޵��`Y�?$�fʹDq�rz�D�T?��i<�&;�����X&��n���
L���L�k�/�+�p<f̪N�mpk@]�3fL��"x%7Z�8�8FG2��cR�s��h�Nӌ��[wY�؃����l�~�� Nk���e%���w���"��r0�
����"�!*�M�:�n��
��Tȷ��,�,�B�xhfK�S��t%Bh���'�[.0�|':Y�OkaQ�d���t�"�0R��A���,�6���U��P�
�`�I�B�ʷSL�d
*7�n�K������8e�XQ]�P�ҐggX,\����
ZM@�Y�%���2�h�i���;��,��ۖ3a��w���S��+mWҧT��ʧv��+����s���j�^p��]���ԅƶ&Q�8lxh�x�{j)}V�������������]��+�\4)��y:I�Wn}�ӯ��i�s,i��.�*�`ߎ�!��O��Y~�P��?ۄd� ��Y��'~�����p�9��:<?���BF�Y7��H<=��,�Lf{���zr��-���B�cq��;�*F��׫�G嚈1o-�Ka�-�wϴ��fZ��+>�9����< b���A��.�q�C��q#�yH �C�ZW�<������*-����q�H�Z�!� ��tl�{d�)�9�Z���c���2H�<��r���u,2� �����7�!�K*�&�ܽ��B��氓����g�<��ο���P>�� D�'8B7<�<|�2�.%r�O6�Yz	����t����= ��g���	���Y���T�.�l鈖4��!��!�c��r�5����"B����Wo�v���ה��΂}'���ڱB3 ��7����oV��5<g�"�+N���^  |}�����R�J@�¶��^� Q�'D�뉫��l���k���iۼ[-*fC[04�8����`m�з�4o�����M�Lכ #;B+��ٜ/�T���>�^Y�q`eQԞ�����������hE SS�3A��UV�Q�	x[K�o�q{��iN�X�@�"
��~4��ZT"F�v�2�ۨ�P3M!��n�����j�/�4�B�#GM�5>����L�C&?pX0��u�����^ܬ�������u�'"b�`2�1��9�tO�(�)������~<�ݑF%��}'�զg�6� �}��
#[�^��q�ZB��z��1
ا�K�w��?j��6y�P^q��i��15TR"���cs^�I��Gw��#�q�p�Te��d������?�h�����	&���!�,bvy���|��^���A��}*��ym�}A�rvv���?�q��ҧx��tE�����U���w^�ܞ�~m�͑N-g�]�[���U��a��_��ǚW������{h��2Z�߸�7��/k*�����v���$�����jť�3S����(\\,w*��}6���@7і]>{~/#���F� �m�a8�̦H�BZJUw����Y����<��A
�k�<bO(���/%=_�+�k���#�7��k��I/��+ߢu�X��ލZٕ]��2��E�Ʌ�}#^	r^w-�\T�fHv;�?�_�p
�\���0�(0<zb|m,~.7�8�(��>7�>8=�hh����@��w�dB:�mz�����C)��f�\ꍍNЌ֫/�h����i����x�=+�͇xP��ڜ��"KT�8D�<�N��S�q�N�WR[��W�W��],��k�Զ�n��� %N;ǋ�F����
�P6�����Q�&�d��f�X���O�,�!���h���^!�K0lEw K�a@�X(FXa	�o�O
��e��۳�9o������PyG��u��q��A�������UPK�	�Tc�Zy1�X�j*(y+��+հ$��d*-n��f�<������EU�*�6N!f!�,z����nA��3#8=��i�f�i���J��n��奟�H36&
�>�s�T٥���45���n��v���	Q��ۉJ���.��[�ю�"�-9`+D1ӳ�VW�z����p�\�𴪱�MF9��L��#*���Gm߮d���}x���z�wC���QxŪ��2Ǖ�w���[�����e@u]�ޖG����&�o-�����ya�o�F7SH�L�\���j�#  �6�l���˃C*ԈL6�1ô�R�>z� ѱ	��NaƆ���ԃ�j¤6����KY�a��9�|�l�r#n�J�7�! 'VW#���X Q�V����A%�<wH��;f��/5�'��	�<���O��V��(��h�{�B��v9e���a)F�R�2�F��>.�F���:�~_p*n��,p�L���'��ݓ#�Ɣ�'�[�i^���ND��UE��8����9��g�,�>�,�_��xb�i�%G�פy|��ڂ�bN-dMfx��m;��6}����!a�׉w
���G�h��ddD��!G��@����P��y��<�B#�"VQ�WO ��a]t�(!�e6ƝU�F��]�c͊869>84�~d��	QY�&M�	�F���s�7L$\���O����꯲S�uJ��"^���͉���O.*�|���t��R9�V`��|�%<sde��FkC�'-a�d?�4-�6hx���GƄ��'?tg�k�p���[NA��!ZX#��
�T�B]���&b���,$�	O���z��0��r���4+?G攙�*��l<s?Ԛ�S���E#[��j-�/Aa�-o��j�pƻ�S�+������6Hꂭ�woS��D�h8�������ƭ鸈-T�w��Pk�<�a����N�Dҹ���q�� 1����A�G�kށ(W���}R{��>�b2���F�c����9Z�@���t��h�q@i@�&��ݖ.D#��!�W:�9�y�Ϊ#{6P�P��:�2��p�[ �.��̔�Cߤ]�*���:>���dY��X5��]�E2S�[�2�^˖3�$�8t�����I�跣�t:&��md!��@�FԸ0�I ���2ϣt�y�U0(��q� Q^"m4{[]{FB	Kq�H�B��̷�З������[R��ӯ�$�ñ՟�i�QG�|�n��y��W���.F��R�#��Ynﯖ0py�#vihab��u+�{�SCyA����˂�^�f�{��.f^�w�^ߓ�<-������0g�ꤜ#�K�&����Q:�Q�5*{l(�1�=��F�}t{b�g�R��g�ƚ�Q�K�v� �# Tl�k?�j�
�z6��.;�L���2:�4}s}9�e�(Z�Yo���]w��T><*fDW��@>�`q�F���1�t*@ꖴ}�����;&���zPk�?��;c���"�jl���^q�qa���a��#�������"k�QFO�	��	r���$�����{�+���8wT̒v�3S�o���F�������#a�G�_	�u��Y�;���ǜ��D�3%��QpY]���ͳ='O��[�Q�����-y��9����4	�㬓��-2�$_~iZ�[�����)�E( څO(�z�SA�Ab�۹��>��z q��y���x5j:=�=��Qm�c�_T�6�(�fmJ(.�R���u����l����Y�:bB� ��4Zӟ�i�d΢t���d��r�Y���,���M���"��7{&2��B��g�%{�ߓ���Z���pF%��#o�'��zק1��F�0M���7���1#�Ǝ��'ط��u�Jv�0�b)�;�ia���Al���+T���	�@�y�g�ϖS���ǅ�NM,k�2�.}���<��Q��g����о(��`X�y�K+��_�[ye0
�5��1�R�C���˽p��ֆm�+Y9��JO}���h]��OX��3�:�l+�l�I[zܮ�BP�X�9��2���ö��ZQ��U�V��eO%z������8���q;�����,o��۞�'�J���N&� �ũdT	�.�����&'��XSc"hD��ʦ"�0��@����p�zE��3�l�״��CxEO7$}��ڞ�x�"R�^���E�t��M �M�n��n�RD�2�5	1��<��aď���*G��v�W��s�c!}��S͢��zl�=��'[��Iz����H
{� Fj"B��g]u�:1	K^K��?r)D����͛�x����1 E1�O�V�]��P��+�GAp�O�����us����;�4��y��k�g��.(��D�FvHl6��;��ߗl}���ԝ�8zK��b;��k~��O�e�9����ή1Q�Q�X����GHgKmL|�>�2i��a�Q�t�)O�3=�=(����i�B�
7�����t���D��'r�����ТÑ�)r�-���}�+�.ˎ*��B��B""H*Xt�g(D<ֳ����~U]6��®���v����kO��l�ǂ��Ȇ ���;��= ���Q�2��-��­?�����v.f2P�I����d)!��_O1U{�[�6X�A��s�À�>�a��i&{E�|�~IH���N��H��B�s��]�t�!�f�����D-O�O6�k{��(�W�Siw�4�Y�Hr��lO�7՝�}���*Dd��A�0(e���湪5����/;�8�<����Zf�������y��^���MD��b��Rnrȕ���4�(�[7r������$Xҕ`\�˝T���og*�9�0Y-��OT��'m?tI��X�7|t��C/]�AALʗ� i�xҍ�=�|��@�|���o�B�ſ�U9���zH����#�6�k\q�zѳg'��a�wA?蠆|�r/�����sf,�|չ�۴��6_���kzq�H�
�|�8P�R��̻/��y���4.>������7�Y#F����y���D9v��~C!K£WcMWa��2����A�_�j��]��������n9"�V����q��p`������L�+>'O˹�<@�6����\�Ժ�r����(v�Fc��Ǡ?_.�=>�Y��|k}�D1s�М��\����A�S�����ӝ�_j̏ȁAe9)�y����#���ܕ���(3�ZF�, - ���?�w�cI"��A�����=:/����u�%V�{SU��E���{ɓsl/ѳ3��u����w���}�M��zb/�K��e����$A��V5,�7�Q�<��?��%MA>��ǣ��{*a��F�H��-��N�O�wqM�W���[�V��������g���A�[�Yu�M�1:h0Ͳ������qQ�4ΠVD���@�o�bYIf��е�N��c�Jk�t���'��o>�>�>��*<i6�/�sp�*#���f/\+&���q��+�.k"�/�w1ҫ�-�l\�j����@�CC �KS<h�S�+p�T��w�:-8�]+�D��$���:���fj�%𼼟�����y@����0�?�����be
�;Yl�����@��I(Hs%.�78ha���i�^��� `���e�u�l�c*|���N������h/���¡�����a���	,#/j/>��Y_FU�[ДK�@���f��y���U.;�rbFK2�]��P�Xb��/�=
�#�#l�^!`0Mƺ
��9����Н=j� #��dbj���'Nqi<�Tu;q�N�Q(���ܘ�Us `�l&�
��p~y�����Iנe\�T�bL�h��)�y��j),�׋�*��Y�qq+AGf�����`E:%X��q7��C��De��IG
�Kr�>����.s14��o�[Jx��k���;�,D�Jz���9�>�� -�V��c����~c��"�N��z��AJ��М�ز�
@V�$���N�rE�E1c	�Q=���u�_(���G�)$<M������&+Q��=7���d��2p5�)��D=!G��N:Tk�H�H���B����u��(�'��{�V����Lx��AN�n�$/%`t#�QTi��n\}^�[6d����&�����8�s���|H�e�P��-gߚ�/�ԗ�0���{M��z��:��u�Cg&�>-�Vns��Zb��\�bxwf��p�	-.Hs�5u�����/&�;��F����Lx���y�c��E*G� �E�&2s$�1�2�3˃�NTqA�$pJ�r1�������`'���B�h��D�afH��\ܱ��LoK��Q/'��j���μ�0?��NF�TmoD3ר)(�4_�:v:A�	��|�-��x���c"����q@|�Sp�?��-a��)5.	��-�����ui���5�yf���@à�*�}v.0��_��|ɱ�}�@�g��Q������O�z6���m��Sl(�5�fȚ�nu��k,�V�yx&P�?������J�{��`jʾvVL�ee&�����������Y^�.�X������5P?@���_T0�V`��2%��ɡd[�{�y�t���L�1��2�{+��|��Q���х;��G0u�
/������I�\6#��FJ:�-�+�o����<�f�����gjS���r��B��W{K,�����\���r(�U�?�#m�(�KOJ6š��A�t� NRڹuQM٩�]z��GR��s�+�0���/�NSF5S/;�II��֩�;! ���	"��4g���?"����
�ƈk��C�f�^�R'�U����VK��(4����E<�(���A��h�`��i�>���7��6�M���3,X���ya���DBZ�Fn�u��?����y�"���SН$���4����~�%6����=X��
&��ǂ.$m�9Eu~*�a'��-���u8T��MB�t�(���X��ːk"�|!oyt@�=�P}��Rn`�%+=�o8�^\~������!��s;*#��v���Q;L�8E�YT��e ����5`���*�wÍ�3xM�Kt�o�ۖ��ֱ��#cn�{�M;��,��W�&�∃�$��|V/���*�)�3ڜ����s �t��$o�I��?o8+$`t�%�ہ�҂��AN�d�S��5旵�Ŷ�So���X1H)׻�:�.E�f�_gտ��>��j]�����2�F��;��;'zEw�A��3���� �4ё+�y���ϲ��K,Ԡ_dV4�+����t�R�k���&�ŔX�^�9Ӥ��Y�Z�ۦ�ѕꤕ��0$u�?��|�q��\��Α虶#Soo����-�!�õ>o��u^� eߠ�|��e!��ǃ�������&_�8���G���*�w/�л4 ��,裰J�T�V�N��<��v��m6Ƅ`%��Y�3�rȦ�C�@x+���v��!��$:���F{2���K�>(@�C>E��|�9�ga�i��QD7DNt�WB@\KUk��]�E�m/)�\�g��<���]")a��$VV��dB�VyEk$��W��k���S	V��e�4��5�ݷ'���� �53򧱰�k�=����_jh>x����u�ZЛx2��k��\/$'8u��=�}>�D9r,�&C�$�A�6@=�-��Cb�ݻA�+K!���g'�Q����T`["���u?��^D�n'�vR�X��U�r!�q)''z�n'�\��{#u�.�n���=u��1������w4���33� �zF3�6
,~�&��AU	�����TF�I���������������5 �����P����$o>}�r��.?�����5y�ħ��L�W��'{��V뾓tg�K�0Ԯ��m}���3�U��p�o	�Q-���o؏Ԇ>��9(��m;�^ERZ"�F�׹8l�9�\E��νNHGӟ(�/Y6��߹Q��90/(��4-$]�k�-��<�ἬJ`��@�$��	�ȑ9P�Ϊ瘾��*��1R$�l�$S	x��?�%!���/�I����A��u������C�x�#s2A�~��pZ���,o�3��Nt�?���7���7�j�s),0zM�
�y3'��yh2��[��� �c��?UlRZ@�a���j3�k-X�=�&����}��S+���:d��˽�%�/՝�I�Ek�=G�8���f��*shw�he �oڤ��0�K7��Hw&�5��)���Af����Ó;�i�n��!ſ�շK���y��K�*�V�f�,�9y�Qj-8��gب��E�ĉRj��U��p]h��YosX9ԛ��Ƹ����W
�O}#H�6��� E\� ط6c�x����zv����b�V9{6'<OF��1ը�d�b��?2�W����?֫+���5� $��e���\�E�<f�ξ��8	� [E�8X$�j믟��x�3�~��ύkEt1m��7,o�:"�<�W4['��-1�s�ý%d| L�H�ڀ6ˈp�"���a"AT|���$�M�����`hs��3�7�p>�rH��?�1)�VS��
��0ehVũ1_ ��ѷ�����y��M��3��Tk,�v.GS����$��R�^���!~1h ��������J�0q�1����@:.-U�']7`�.��)U�|N2��|w���@�V���8�ͪ�Qâ��@��v]�!M~+��C�Mhٖ�p�� ���J�E�_٢�XX���	���`��aδN��)]*�� ~a�=�Z1V
~޹��hM���+�z��L9�uX2M̕�H!�'��-�z^XL�e(�;3���Q�
F6�gC�>�y~�Ǐ�q�R�b6�B�W'��4G�Vg��s���{����,tpa?�?���'ഔ[���e��L��<E1C�kSPA�\�I�� �br�%�Ec[)��~Z1�~�]�<�Ay�N�q�&������ .dMdq�|�I�UvM��X�����#�E7
&ݴ%b��F��~@U������obv�9vˣ�=
=�XlL�����]��`���
�J����@W����e�A�P�\v��
�E�B�F&E��&���e��(b�8�Z6���S��-�2�?�؟�G+I�m��@!��N�w27䰿�e3:v쮫nsRI��~��_Z]��q3�@���O���vD廔���8�&`?q4��� �-�頊A\�e�[���E�+��xϷm�����dE�v{G�s�@��]�J(��I� ��GFmM��i�l<����.7:��:tt�Ѝ�b��P�['ǲz,�>F-D�t��$�_p��?N
��X�xC9��A�, "!bJ2�t��.+
�_(�?�1��δ���;������kv�i�U1_�z�EMT���ҼZ�\!t�a�"���u��� ��\n�ut��U�} ��p-��>W��y��g�	H�M1��
�D�9��V+P�&Ҵ�!o�5B�'l�����_�
�#g���Ѫ)�j�Z+Ͽ4׷Sb�'�g��� ���^oV������8�a�A�&��n�f;��"$x�<�%�U�asf�8�'��f���krr�5��\xȖ¼�}9l��U��F��\�3��OA�~\�����CGWM-y:��q�}�ܒ�tgr%t2a^�M=�RY��H�jV�T8���	��������z���[�#�RB�Ս�\����N=�Qf#���HA�$	�H�������k��6�턅���Pq8	g��Z�l)�u�
�/�II^�BN��IB��<�W��JG�͂���{t���ʅ؆}�f��^%�4���B�,�e���<M˰�����Ws�o����Q�j�Þ��]�SF���DJ޶���w6ٰ��wS��_�9b�v�|����^mᭈi	����� ��[[���6o���O凨���QҪO�Զ�3+��)��4[�>���,͊�wc�~�M�-�L�,���^�vz�ǅa��&"�\Z���8%�
�����ۤ��d��(.8N^�6!=�j��$�y7��n��殿��I�PE��ru�'�N!�j�eq$�+<O�S|��ӝ��0���}`��ٛ�@[E.�f`���u���Ff��G��N��}���2�X�/]+���{$6ҩ`�N�H��C�/�T��Ь`����k`QZ6lp��t�m�����'͠N���f4����*%�&Cת~U���4��5�z�/�����m1T!2(Ҹw�[�NfI3C����hK�qa0��@0���lkA��=�)��'�����o��ng���3fP�I
��~܂��c�`Ms�'e������
����&@m�c5e��%^w��JTߕU�we���;�R������̆�'�Sض��Y+�n:���76��&�||N��K��z��E�G��e���򸬖E$!b~�gm6���"������#m`�����j
{��&���1:�{����bdY����8��H!�u'qZSq���"�E��(ޱg��7,|�c]����0{����Ӻ�FK����9��e�3�Jw`d��9ӕ)�Aw�f"�Z�H&>L�e�3��V�K|B6��I��ci���nRMN�*S]u�ゟg��:�y�AxcP(���)��Yq�q
�	]�
!#�^`[	ෲ�����
�M��ofDZ���ׁI��{
F��k���΃g��c��sp�r���@�W�IA����l�T��<q�� r�4�jx1L�*qqKDH���n"OS,�#���B�B��"��/�dv~E&%b��8R;�Z�J�2�^���{�Z�@|�<���4!���[Y�!9�V^��S�h&������q�������p����$\���$�[����I��Ѥ������lŘǢ��p�&Ed�L��a�� M�=,="�����]Ӭ�,�o��4s��'u�8jwP�v�i1K>,��@�8���t��:�sJ��<&=Q�T����ʛ*g�P��ӯ�Y��.L�1[�Y�*{��Q����1g��$"��	JRr�R}xB��r���Vz�M�.%����\�=wG66dPw��օwFG���y}����ʲ�����H���(m�[�o�^�t�U��T���
w�S�]'��C<�`���hj)\�m���|w�Dh�cț��k�m�4�+�"�KY�2F4�M/P��KXd@m��B�m�~��=�u��B�P�2s�ٸ��&zy�=s
AK4A���T۲KT��{>g4)o��x̜���^��(fDm ���9�jW�
��q&)�4r�N����!�-^m�� �X|��I��]j�l�6D�_�~�2�