��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>>�Htd�	5w��O�̽�]�ɽ!d�`���٠�L�3��>�TI��Ft��"�e�3j���!|�x�����S��D�|�<���2�5���cBQ73���ƭ!=�҂M��|$�5u�Ly-������a��^���r$���M3d^����H�*���-HQ�w̓�se�*^�����C:��#_���������
��݀q� Y.vQ���3R�a�VNW���j�&�V�c�O7D��ؙ�Q�T͔�֎�:�Ɛ>c\�^o�z%Wڼc=�a�+�N��W� t�5@n�4�<fTy_f%����@�V�t�=�(H�G�$���>�އ3��x3�[_�YU��/�_l��Q:�C�g�� E��{:v��rn��)W2US8P����_{�S�k a��+��H,{��+�U7܇dO\(+�sN�Vt*�DS�JJ��?��%��$.���g��!i���9b��N]~D
O��)����ۃ��Rͣ���)���=�v��Y��)@(9����#]��֔q˶LG%�3��1�D=� s�G@D[|�E1�,�h�޸�G�H��4z̙>��c9���ZiK�8�3��8aoʜtC
Dl�a'��O��zޥs6� �Z��˺{@�����
�h>����%�oA�l}�Ba����x����r�{O3��wj�%ߥ:*w�s,5-��kn0���sr�L~ڴ�i�i���+L��s:y>o�J�v$����rlu������NҲBP
��>��!#����x-�zC��<��Y�F<\yh��=,�8C���zz��!�����U4��/}I�!ݐCL8�v�&7���HB�<��P�4D2�qҘ����}�/��Z��;��y���ŝ>��7#�dvs3� �z��2��/@��D����|��ך�79Y��EA]��WZ2���.����ob�<�����U>�O%'q*k��)MF�;���n�}|ec
��p��ϙ&�μB?�5�R)E�[��剈E溾�%%R�ĉg�f�sjTa�\����ʨ㋎S��-�)���B��Pl�y��C�!G�#�f�-�x��R��;L��J�����p�M��e}�ku0@K&�c�E���Q��Vxp�YP�.���,���]��[��Ö��p�-L��b
�6�}�k6���L��o��1���������Չ#���f;�E���q��{�����?��i-�:�9y*��o
~EXDB{m�[���\���ΠY,߹LMJDm�/[�*��
�f_i5S�+R��oA�,�jH~G,3��t�Nڊ����"�CL�f,�8l�"�j�)l)L�|m}c�}E�c�v����B��-K�=jP����榡�6m�:Q>ڢ��h�Bf���� �V�Y� ���AaV���L������w�/�|K��+#�%������{q6��c7$("�.�U�����{=�o%Lor����6�x,b|���z�·b`߬[�������+9;C�d�8��`��ޤ_oj��)Ι��,^�ˬh�"*dGOf��-^��`�+�3�M�DI#=כ�W~A���SȊ0���F�'"��Z��">�M�E^�'�e���Y��6��h�t;�yk�x�����Ċ�W!ˋ�9C������q��x;uPDP�O��b]^g����
7�O���Q�(#�&݌#���rG
�c� jF2�"���j����U�>_�]�G�`6-�ې+�r�ܠ깰��|�^���{�4�5��j�o���F�N!M����`�8[ڸU*L]=ۑS�:�+�eJU�͇�[YAXAͽ�{?��	*���dP�I�y�O}-�0.#�;s�	�d�=�� q����R&"������d-{d�dJ�Z���\>�$���J������� ��S�qшfb	.�߼t�JG���^�MKnD�Q�,������� ��\y��;���m��ghro��^����%E�^31{=o�Χ�u'M���?u,c�s���WF����>($�3���`��Y�YL�2R�����B�r��=^ekiwH��(���tp�z{A�_Fd��3T�])�-> $����ϋPr�]�'����f`�4�*E%��ĺ�0��9���XD�j�:�ĩ�r��l��]���I�!H�I��	S�b��M;����Z��3�s0E�L�
�HK�lA?	�jf@��RU\k�tJ�2QT�����n�u��k=�l��Y4Ņ��v |�P�F�Qjv1@IꟂ�^%�ju�7*|_��7���]�.��E7�Y#�FiƊ̔]���h�"�P�O�5S�q
LE�HFA�\`���b?q�A�x�G��G(��	!HH�N���J�k���>���K)�Dxo��Z6�t!�"B/��7��Ѫ�!3��R���y<(cx7�r�B���_P �m�8���3�&?� �6�[�#Y��Vwv�����c��7�b>�~ e��,"�;�c��t���[��qߍ���>|����u��bS[����qg-B*�)����W��Q �g���y��c}*�����G�5�m|�e8A�3Z�+.{����$�+99(_	�hu�=e��#�>�צ��`Y����tO��Fe��	e&�)��8o �8�ߟ�T��_!�!�5�B�Bٱ�q�$&3P�қf/�7��*:�K�4%�e¹��ۭ?F����";mT��0W'$�W2K�+���R1������J ���U))��/����>�3���Ʉp� юP�M聪�-��u_��tr��k�3	�F�x��r����B5�҈w��w	?;��!��PU��)H��W0�P�0n��*�@��DX�N�� ���Pv�xS"�u9v�c�Y6��4C_3�"�!��C��;&�fI|F+Dż.LѮϻ��������*��-sR��8P�$�9��"Ϻ_���l��]K�)f�9NɃI���(P�~�����k�P���i@ޜ�,v^D�Od�%z����+bW�u1�#ʈ�G�H�Ի��3n �Gz�I��@D���ݜ��	�����]�ڱ��[��'��n���5I�G씃K0�]%Mk~���3;�����U
'���瑉G�~�:R�5�eٙn�^	���R���'�ͬ����(t�0��8F;.��>�Ѝ?P�\Um�cl�+��A8��BE�)��u�]��ض�����+�Q,�忚���@�2�#����r�I$Y��_�[?w���{ʽ���m̛|n�<���q%湊@��;�U���@�R��)���A���S��ր@�=5�7�!{�WA��Z^p�C(�<�D�qL(�\�u��=l.�����