��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn반lŔޢa0�ݙ���'V�߻��i��mx
T�"zM95&Dq����gMl�����s�V��P[����.,��ͪR�"wߢ?�=�z�ۖ��kk���Zr��1�g�{�7F��������?p�qR�\y��Bq�a@�҂��4n���z������}�X���Q�1+�n|�̏��-(�,�����Tn�(A~I���UK(ܕ� ���g�.n}�j�"���S���x�A�s.7fo{�V��y��S#:I|ym���r���~]BMD� y埒�尮C��Mz���	.���@��Y��}�2m�>�݌�i6G�t=�����()-U����b�j��!�KjMʒ�&��4`5R'���̼������ ���s$����Bp����^b�~sF�L�w�o��Ԍ�?�M -�dW	���r�Khld`w{Y����{Y0�Uؐ����ac�󵯒:�]x�?y,�a	8�D#Xׄ�e���7��o>,�b֟��8A0��r�w����Ѧ�z�o�;�BqE�;c[ի;�ULst�Ҿ����N	�PJliw�VW������fC�k�ڴp�7y�Н���6!C�
����������J|�¨x+A�"���<.Y"��3_��uJy�}��c���\�SQ?`?��MMV�MV�vn�?�ld��%��,�!b;ը�l��"��=�
V�/E�\b�9�g�v��?�ӕ�{Mء�=�b��W��@o�(�:�at�Q�r�?y4��tF����4�n��>����x\��{�$B!�5��Q�gi�����ѩ��3�)ً��	��UDd!�S��� 9�/�)�᜾�sU��A�AT��&-���F<��F���-j�u��S��8�$��������z>�ʇ.��a�l�8��@B��`X��M���q�?��7077(E��"�K@�_���D�X	�\\way����G��6�@�j�?��+QϹ1��WpV#RW�zn3���a������� 1��MԎ����+����f�d���a�-\~@���nGp�7���J3a8�F�2z�z��Ʈ�;�P���:Za`('R�P�6�|Y�x$���(��BF���i�������^��즞��<x�˝/ՙY[2>�� �@�e^W�8��M�*�����Վ"�RA�Gd t����@u`�b-HզYe�R���h�bL����F\8��‛������_RY�B�y�c�JFH���`�.H��p2�p@ɇ�ʦ���9���3`UX�6n:<%��{�w���~v��!ϒ�T4ؤaJޘ��!�c'dЏ<�]���_uB�DZ�h���f[������U��n|7��q���'�#��cV�:�^���?�6�s���3����������W&�?�A�����K�o�6l�˦k�٧���yAڞh�
 �X�A����G��F{�!:+�����~�tB%ҡ0�H܆�y�g���%�h�T����d��7���ʱ@�������;�����;w�v��4M�k��ɠH�a��<��3,�@1���8,�$A� t{�q%��m��xӕfb�g���fӵr>�XjA/6��+0�O`�6a���Go8�r~��t�`�:�x��fw^	�).�{��&�=��Ů	s�q��}O;��]<}�3]9�ʩz��5� M��w���x�R^y��ɺ�o�[�B��b*���#���<�:��{�D�'v�be%�قO>�^(�ҏ�G�[+dUT�`)M���WV���*�]�+wl����<�)!#�t�?a�ĸ$P�x_JX�~�f���m!٨J<��Q��r��������O��
-3�f%� ��`:���oEK�$ �X���4��������H��w>�s�$�O�#{qB�Gދ��3���E��0�SW���(dC��6a�,�t,d���k�z˿��OZ��%}.��8n�5�\��DI	�M-E��Ú�W����s*��*���Fj1��N�T��˃��P�cEs�[Z}R�pÙ8�-��}��W��~_g5ŧ$uc8�e��B��W�V�R�
��G�^{�	�_��(�'�F�H��g�_";��v���;���m�'h�6c�9!ܩ�����Uח�%`=d.��1�9:It8#�K�c�ˬ~��!��$rr�Ԋ�eڌ����K wQ�w�Ё�o\w�7<}�������vJ� N�`�R0y��kc�"��DE-�+�cB�o �cc�Iv�.N
�L=��K�᪡�^���у�Q���1��q�k���N���"(��Am�Q��l��p1z��w�j���(�<T�":�8�M��]�A?�����>�Epꕾ���7��ޞ�]n���j�x�N�Z�=�\4�ޒ1�E��a�[�����.J=�������.)-��N���O��~�����Y�����ݏ1��kp�M'�ҩ���6>��+T4�=ܔOg��/5�#�H�F�1p��n�$��I\d��v]�z;�ざ4qO��k�b9�a2b�M~�k8�s���t�h|�½��j�L�4��I����P����F��24�G��?�CS+�GDx��uf�Lރ�Qf^�YS5u���5�	�Me:鬛�=�ޝR�@�)$����7�rQ4k��J��M��s9|��?ݼQV;�r��LC�Gz��#����:�gv�@l�n�������]�����;��%bn�pBڠ��jS�N�b����XIYN1������F���	��/ �|�Z&b�P|��<�HP*�����cO�(��!&tYj.D ��	��s�����n!5�Nz�nS�9�VEt��p�z�n�/�ޢ&9����[���Y������]��fZ���%����r�[u��5ݾ%2wo'�6[�K��L������Pn鎤���?��\	_%F��ݞRɛ,���e�o(�9�fR��Is8>Xm2���e����s2�j�g¤ 4��жN>�$�jRev��w�����N��a���؊��e�,�(�X�˂cU�E2 �c�p�O�˭��,���W��r���۽�S�o�Ϡ紩r���R�W ��j'��a��?i�G�#�����~09�^ݥU����������-��쇽��R9�a�;������*��zQ�5�4��u�;�!�OT�F��!�$W�0�����9��N�&��Q�MT)�?��7��²�)/�%�lP�h��&�.`�=q����jF��~��VJ��qѴ�P��o��|\P�x�3�x�i����r4�&/f}��� ����?���7�p�����7�)ᩏ����@�D�W�B�E%n���䖚~�Җ��{�?Y��6J�XS�������aueR�v�ɡXs>ā,�|�o�%�/e�S�ո4��{��}I['R�1���o�i%p-ۿ)}��ZF���-������l��ZzH�Ӻ�2�h���8I������ΖJ"u���9r��� �^Vy��nt�[�|G�K�k{�$�����5l۔�:��8��F�G�`�rB�0s�%6�>�� �\h#�鍚�V������ϋ}��<��Ę�s%qdH���m|227"�4�����
�d�j�
���H�C�$����� n�N�_�F>�~���ZZ��w!�A��Aw0R��U@�N�Ϛt %DM�;_�h5�Ž�dg�p��i��3V����܍\33w����r����yw{��ً�(�|���Y:�^��}3���}KF�@�`~��1�5�Q~+;f�X��'2z�n�orH�ǙD�y`šh]�p$��w���V��R�o�lɎ#�f~蘒}Wk��KsҎ�����#@M�'�Zؼ���![�ڮ�м��������Z�7RkQ֌�6-߀�Sܜ�ҁ.����SY��׎�]`��C� ��A��R'�M؁�۬��9_��g��>�J&��z��q	6�����]EC9��|.&��8�����~�>�#�U��1�Ӈ�*��e�����G�]����B��D@2F`�K��'� 0�����8ο�|iuʛ�����*3��ˇ-�'	��lyX�c	�턾-ڛ�bN�����V"��NO�d+1[.�ұ���A������5���Æ���2�����wC��M��L'8�������V�9"�b�L�)\+�vğ��=]=릚Ӊo�c��|����P�m����r�K���O΅�`�t:) NA�47 0���%��7���Ɓ�/�-o��p4�_�G�r��bX���>V��,+�NP�v6���#��w$��v��<X��w�� ��X��ܓD��Ja�Bɘ�I\}Í?<ݤQ>�����⍝%��CDo]�~ �ZI�[��/M�ɓK`��Ya�6o=��M�;�DvP����ȥ1�#�MA>���x�?'p&�)2g���Ic�6�s,���.�ո�ǽ���5S _r{n����7;��V}�}o��`@����f�����1/�z�CV�g��0�j�q��F�3n�9`���ZDN56osn.@�y�ݥ{)���i���OV�y�K��ީ��4�#p���H ٻ�rw�!�S�X���"c��Є�WZ�j��.�}1a�m�P��
�Dm#}\�e@1�b�9��~T�pM�0�u�4kz�R����g�/��7G��ZX�z�F<��qcv��)�+j�bs�k�H;�I�����RE�c�B�B�D�ʝ�L���.��s@��aK&z#QXa=�v̈́3e�) a�Z4�6j� �kY�+�ד�6�'��`��'��ǋ�K���I�R�B�v�U��P���2�|b^��>J�M��UN4S���Kj�����q��8�ݻx;f,��笤9�F�SIjQ��?�Wp��b�*�h+��|H,�*2Y
��~K8�m��eF��!�I�[ � �xs^Fb�M��Dvv`�6��l�9߫��7B��F���\�ﵜ�WlnD��z�!��V�rn�n�'�U�I�]�3���'{�6�Xc!��jI1'�2�~ȟ���6�7l�$8{�~JP�ܽ����_�6�.KK7;M��$`��Y���L�h���)y։ݟ*���	��/�q�������C����S�]A����%�D"	%^8����Ly�3=��v�n{_(�bA�����y&V�K�_�s�R���U�퓨Fxrk�X4���-�\��O4��́��^J��u"yA��ʂ��#q%^G�
�A*n:��{����,}P�j�v��VI��=L��.�V������ ��<>C
�Z�&j]x�}�Z�2$��u���Mϭ6�T3���V/���0��8������(#S�0]0-2V`�3�w��S�saܺ��,Bƚ��ˮ7v��[<�cyFx#�跨є`�����
�c��3�U�Ó8H��">�v/�QU�VZK���i\�K�vR�Í�e�Q��p{�Py�:`�>�f�^��K�RK.�O�OǄW,��쮖#Zu,ᡟd��&�~�c۞�g����F��N9Uɠ�� ��ҧs�p�&�������;��~t��fG�0�N:1��R��L��l�G6��!��P�}kH�"�8|c7�t�x]^#]���7�&���5�λ]p�$2YkPMقz��3۾4�RhZU>P�fQM.MJ#��B����9��{��M�J,'w�_��(�S����r�t�=�m�w$;B�j�{�J1/H��Y�<}�c��g�Ȯ�{���]��n���dv��MC����U��� ���T���?��Q%���#0�Y���)²�'����9�h��ú�Y���<�a���q�����I}�bu�o�����7	��3�lF� 2҈#�J ��A���s:�Mq)� ���_������J��f��N�Y���lHz֍1�)
c1�@����m6�`��|,]�+H''UE5S|�?D�Q7�9l�ꡏ=F��T*o��K.����������@o,u�%5g|!��d^��Y�An<b5�)ߓ�.�^S���w�m:bĨvv�g���0_Ew��N���p��5nY���M{�A�]�F�������'ĆH�AQJ�q]@8@*l|���W2^TU��9(oQt�T��Ҳ�t��L����-V!;[e���i��^[�)�AR��~��kW%ЕX|S�ԫ\���_섍��s��j�]�8Y��t�� � +Q����nk�X�8�s}���RM�ja��ڂn������˿�}�F%�fR�+R�)�9��j���:_%��D� b(�[�ɬ!��vJ*fh�G	��R��By��C���v�(~p�f3/�.�� '�{�n��4�}�Q��(��ױ��a�P_ioH�k[ �b*7�a�L Ko@�����&N���谡&(�n�/�`�M�9��t���P�i`6��w�\^r���Nѕ���Ό���!�ݻي��4����A_��y�x�������{�h���L�6�#�.w:Q3����dt�{f�֤�[H�q�{T�dH��w?c�e@O���SG��O �Lf�Y��c��$���2����/2H�9
�<k���rE����^_�����^Z��r�փ�0��k@�4�s�����E�ˬ�h\��BV�w�K�g�63�����O���y�ַ��'C7����}d�+����v#�����,���N��8l��Bx�(����e��l^�(>Fi?Ӡݽcc.�~��B|�x����`${�#�Q�~�%�K����J =`�%�35L	C�Nyˠ~���A�d�aRR�)�8ҳ�FW�єHg���xU��S����^����P��{M�A�¢&�f���no_�.!z��DK�3��,)��̵���^~n�;��� ߘlZ��#�ӥ!�h�Ya{ר���IgSS�0�2���t$��@�Jz����� ����1,G�C��g�E��ĴNׯ�í�eJ	��>�Iж$��T$�*��5ԃi���\�߯��-���M]|Nع"D����Ox�'�R3V^��A��fLD׍ǊP�?�ٯ�J�1�����`tw��Б���ߘCvx��B������(�p�?`���K�����:e�WP�˔����~�;h�c���!��N���)���0����+��6�Wƥ�( ���yU4������p��8�������r���!��;s�7Wf��2�����W΢<!Ӹg���R6�ul��VW��HvD�^ �0�WW�S׺O�2R"=Yu�Y���R�ļ<S��d��a���۸S_ �9�������5`)�o��n�4@�1Am�ƕt�K�js���V�c�Ϲ](!��v�gzo�i~3�1efFz��Q�`D�/�Kd��2_�<8�a��N�/a��Z�0�V��uk��z�9����J	�M���T�+K�c,	԰�D1ڀ��+���'�@��2le�)�1�0m��5��~�qf���Է5��%���� �f�H?��f��-*�v;�F�*�`iSI}1`�!��t�]b��_w��v�Y���x\v�p��,n���>�@�g�Ӎsoy��<x�6#q�CVː6Ժ�,�r���r�:���P=#4����L�~l���_d��Cp�Y��ϋo3S��N���mk�������͈�ژ��Ը,)a7z��(�9��r�nv��'�V�@�0����v=ޑ��b�~��ޝ�8%��D��u�p�������Q�]�����ݮ����Qq��-�1�_�Z��,�_�pߞ�k����� ���B��V86^��Vo`��LRW�dS�w���pu��S}N6��]B�*��2P�j��Z1�5���1��E�t����ݴ��c�}&���{�����ś��?��k�E�o�>QW:9A����$���riF��Ѽס2E=�"���/еL���0����]=~��&O:��+�����&�B�S- A��.4���Y�}�\ݢȁ�R�|�{�/9�ܾ�'غ�+���5�w�H��j�xU4�}�m�̬�HK��̶����2�,��󾲜�T�fv�K�V�4���z���	Rԩ~��1B�ٯ�2*$�ߜ�{%!�ץ@�����`I�t���-@_�4��;��B��R|�F��o۹hn����zv4�9Y����:dqCL/�I�?�{�ۿx0�G�,�uxs*�Z��Wq�����(<���DHa�n�����)/�F�N��-$R��4f�k�ˡS���s�I���;2�)�J���9�4bWQ�Mo8��jy�>��A�j,���;e�=�>{��|���?*�[�<��H�f.7d� �
$�ɿy�S��+�R��}FAQ ۝��y�ꉶ �x�w�]y�׹r%�ml~N��&[��TcT�gL�p[���UI��'��4w��{��9�g3��Q}�n��.�I$ck�P.T�WlD�~B\��!ѐ��.���L��޴�	���)�V�&r�i�=J�8Ga1��3g�<It�:��i���*x�g<�O���C����g%���oCZ� v�Pd���G��D;F��<0ļI���W�c�22�(�)B6P�+"D����#������e�P���F�_&8l��Y��D9�w"���g��?`&~�R�q��ec�O?�%�h\��6���|ly9x0_֐Kz{�
܈'
G�[�%���Fv�|Ц�����dχ���p����r8�tYګ~�x��P��D(��aV�a
{
90�w�¤#G٧�/1�9�"�T24�"�sMV�ع��)߉���,S��b��b��ε#u��Q�W���ф��~���L�:�m�K������{����ՠ2m3����@��S��B�M{��(�=���e��	-�0�E҈��:[I����m����>`|*3(���_~N`�_"�M�/�<p�5����3�}8n"VC�\�~��,q=�	��$�fI��[�8%��s�'JC�:���Sh'��sV��$`t�D��k����u'�=�
�	`�p�8eB�LR�uD�070;�c���j��0`���m08l-�%!g9� ����GG��fi�.�cf�ϴ��oY�
�ܥ�yOX�����Oi����?P7P��'����n�A#���*,�o���򖦍t�|Oԏ>tK�)6l�-�^u�h�����/"��Z[硟�S�2�ȎGa��ӗO�"Ί%�#`�s��B�nH�A���ⓨ���~z)9��[*�&8��X���o������~��V9S̛���/ֈ.�\ج`dz�c�j!s���q�<7�?X�+nD�qU�^��J�"�i�inZ���� 4�T	2i�yQ���D-�#�@��ou�5%�D%������۝��u�ѓ�P ��՚��F�w$"�;Ѓ�h���T����s�v�☵�E�g0�A!Mc��>��|�}�CtK���˙�X8R+6Z�4��M��tcM��Rk�E~��g#�4	7�z�(���p�� ��,���6=W/���|v����[�I��I�5|]7�Z����:Y�0Jk�#M/���J�Ւg��S���V�5�����¥2Kb�����Yz��_���y��V��ޅ�j���o�����*�w�A�'�7P8���JȒ8ݘ"_@H��Xc@n2���`�
=6G�O5T�-��=�57z�C�7Nxs��]Ǳ��9܎����x5��>>��::��/�'?*U�@G��=��Xb^����#:��l�?
�4��?� �C'�a�D��bڢǣ#�͡mo�B`e0��c���2ғ��y��4��٫��",����h�k��� ����'�D'�dW��L-on��$}\��2@x8��8pHP�;(�;u��߽u�X`=n�N��Y�9罣g��Uv�����mB|�X@�����ݦlb�n�Ɏ6�������r<���1�p�y���1��(��"#�{�>�X&���f�L�<K-��:�������|�7o���P��G�?D�N8�"Rs%b)h���m���)�����/3cT|a��M��^_Mi��� n��
݁��}_��2,��Uf�	�P��[|�P�ũ��t�����/H����ta�GO[�mҗO��T�,�+}��ON��#|��@�.�`���*Hu�8��*t�1�6j�'��4��hYt�p۶��quo8-As�.��[�2��*���t�u���n,��0�9��8���ּe^��"�u��$�%�O ��!�׌9�������n[T���\'�y�����l�����;���k��]?��զ�ʁl���0�q��qꩶ�آ=B���#a+	u��فx͸�(�h��1˿6�����!a6������vÒDt�/le_8�wHy��5���Ѐ������W�L�p���xR����:��R:W!��(U��2"�:4hM�xƓ�O
Grٟ^dBf����	��ŏ܋m��t��]:��ׅ&:�pgČ)E��� �!��W#�_g[��x z�f���;�g,kr{�`��Ә,�S��y��<���q�T��R1�����yJ'}\=���e�d�>�
y`U�] qr��)v��zh��Ǻ�orX_s�s rᜌp^H���	�"0sNd3�4X���)1'hx�n8����+Q�Kz�J�:}F�]ۤ��zQ|}���>r~��f�f�c5��P�qΦ�j�(�N��o�+��>^'��:z"��ۖ���Z�� Z�Ur��T+�Æ�R�ɭ�%&�AoK�M��e��U������6А�?�� 7I����cE��T�Nr~�B^Bp���߱�#���	��ѭ��T��trM�K'�>�Op%=�D $I&���{T���`�u}q���~��S�[_���n��{�6�Z��(ĉp�|�AʫD����͛�#��U*P��?�8��"҃�W�u-�63f����c�Boǃ�ľ�����:%����NM5�D�Z��>!m���.�l͙]/F����&z3@d�R�����T���&`��;�׉L�93v�[��z�w���}�\:H��L���G
K�;O"QZ�$�kY4a�o���f2�dF\��j<n��Ô%3�S^�J^(m4ٮH}�f�m��xc;W\wȐyG<d@gnFQHC+�����↬�t�����-6����Dyz���4�?)�ݱ��M���o���Sw��*A� �>p.!'W����-r3ǐ���w7I�E���ʦ���7(0K���'B�N�Tѱ��jB?='zf�:�lOW�c�]�`��Ʒ��:!�?'��$t%�ȶ�FF58�jtz]ŵ�)(����e+ꉊ��;H�2}"�01�U�[�6��<O�M������Oo��ǍA���HUs�y�`TQ�	f
 k��?.'#s%6u�	���ё?InI�]]��dB�E��E��Ul��[�Ǿ�@H�dOك�]�p��uo���a�|�}׈����pΛ����_T��<F�L'#�u�&r���m�����П�HB���e \(�*x*y�X[�@su�9�;zK������&7�g��S�{.2����F~�#��A��N^T2�w��J+�[�t,SS\���S��
w*۬ ��Z�Z7�BiEK�;���ƑTƿ�	�[T�EOY]���@-�y΀+����g���ʒ�B
�&��L��/�+��-_��'��R��=��-���Z-5�̺'�9 O;���?|�pU�Wh���tDS"�����ꍝ�J��T�@W���'��:V� +B�r4Cܻ;j�L9�.o��4�^g9����|yE����_L��Q�h�����a�Wa�{z�曞�8|-+�FPS��,�5�N�84d۞��t���H/�m�'0NN��,r�ȬHL�{ӳk{sK��X�(ѣ
M!�3��qpi�!>{�T����T�׿�2��3fgU|}�; 0����nm-h���p�(b���. 5Yg2�gV���(	���y��swNnJ��ַ=:���D4��t�F1�p�9���[EJB!g7��X��EG���x��q4ө�%S��������_��և�������#��8z��7�9��6�����$��H��� ��]�����v�#}U�j�;i����)�^ڳ$�	��.��^y�b;8��*x)�J��r8n�x���J��q���ɭ��ţ4B	�+ӥ���v�㫎�������Y��]�A�����a?Ĩ�������YC����|��U��D�!ߤ4_U6�1���T����c��d�T�~�M��3���d�0(�TT��h���K��=F�-�|>�h�an�A8�  ]a� ��x�r�ʲ�-is�9�e��o��KM�X��G�{P���Y്�ߙ�Y3�q�(DU&j���)�,lf�.�<ڪR1\���2�Z5y����Kr:	�2@k������V}��pO�����2�9U�X+P��@�6�����{�#�=⏦|nRg�or��<��)"ˌ�O���������v�tkGb��+yѮ��{��Nvs5=�vvg�qv<��A���+wIu~H�o8@���x\2a[��d���������R�׹���ވ\��񻍜���"��S*����%5�>
���u�*�)d#�_�M4TP�0�v��R{����5D�m9�mt��ɥ�Я��j_u�v��!���t��fw�7$?�	ɖJ�7�T^�	�vS�~��\���;V��M�k��.��O�wC���ñ �'`��u~S'��5f�%W�i�c�_Ev?�.0I@5�l)�����o�u�MX/T�����V�t��u�8ׅ�2����5 ���ۋ>�Qc�SV;��7�Pɀ�_b�cɿN�%�r���2�f�%��n0�ﰬ��L����*����4�t�����T�"��U�<�F
��L�a�ĠUё]�ZR�g1ﺱ��7�����1�w��噋T,F,sǂm&+���i��E�\��$�%	Sw�_ ө���,V�I���Gփ��=8ny�����l͈}�<�Q��O
���Sȳq�R\�^�0N�o��̈�ͤ�~f�g�q1�_�A���>0ӹ��QLv�-X�#����L����&�Uh�jߍm�L�����zr!7|�H��}pֽ�zb��2=�/�\x��ַ�d�Q�3�V]P���>Z��%��Sٛ�p0G�����Q2��o�w��IZȗ�響������)�qh����)���x��.�Xr��������2�TZ�;e(cq�.�n'��>�&�G�'
����҇,<���t`MP���/RY�V�z)]_~�
ͫ�?�p����D+� �,�qO���ͮQ�K뇗�d�E$�?�3�B��W�+�m�r���i��>|��+�	����l��>Y�|��N�(�K*5��)r�=���.[�dT`����ŷN�6����S��\��7 �������Ǔ{��J��S��Ū"��|��^k������������;i�m6�Y��{*����ra���l|���Y��8-�2���N�%v� ���GTq��X9��Ŵ��vG������҅��s���X�ā��	&�L�#~|�9����1q��t��0��2�0�T�;��e&��O���bf	��)��PV(O���a��Ө��T+�SI�Q�*�0���Oa/�s]%�N�7��*�Û0�X��Vee�l
��&�A���b���O��� ���}�;�Vm�|�<l,�m�J������?�X�9c�hes�e���Dk߹*rh3H�t��W��T��I��$���׹�SH:,���׏ߍ��Y���I�7�G���r��+u�����]<	�3�������y������HL�8T�OQ��U���<��4�v2K��9碗�G�� ��G�Ӳj�zG�F� ��B~�`������mQ�(�����E�Y��&��}�Ab�����\��wbL׼�G_�I����+C6āˢ��H��禉�j�=�ڲ��&VO�w�φ<��r��W�������B�n��Z� ^�#F�<�i�m��!�'0&�}��\���6��__��۲���%����w�u ?�y�A�TW�דּF�]P�~e�R<��a���r)��] N=�`7��R��3d�SB�3v�Z�s��+���"���d3���i�:9\������O��l�e;�|N�#>'��&@V��Z�]�1�����W1\������v0�L/O�Ά6o��
b�W4ǢBPOye��n��������-9�-z�XOH_n�9=�I0=8o��Mz8/}���,��C�'9'��RK��U1n9v��8��~m;� 	'��X`�o���1́�����x%`��9ɔ��H��ɉG���9>	���O���, ^eY^d�
�R�5���w�:�A�m�2�P5�;N�ЬF���J�͖�}��+2��GM���I�����۸����h�t���
��p��w��j(��yhҴG�1�g�wI�X����U����M�=�4�i�N8w;��� ����y����,�Q'���"�e�<H~�����!@c�^�^~?R���/?Q���+�H-{��<w��{��#-d!�����܍uR ��@��cIكI�e&�O��C��pd$���^1��Z���׾���7�ȇ�7�2�{�5Uo)�?�`�Km�UE.�k�� ���b���9u1?��Ϡ*�C�^�0�
*6"�eL���hv6�?u�6��.��.AW�[���}�G��^��l�����Kk{],�u���Z�z~6�'h�{
ﳩ�s+o��Z��p����盧�ή�ݖ��_0�t�G�"�3�J���i�{V?�B1G��ش��MZ�)��/,�����9��QUz��/x��G�R���0
�.o���t��f�̒���4��
�ҠC]5��m��	:�G�m��E>w�Y;�A(��m�+7�$�+���Nz��¸<h�P�l)��je��ׁ�r�(�G%"A�zW<�B^�z��>��Hnb��z��sc�n�����ڗ��ڍP	�\WlX�oY&.��Q�����bO&����r��샗�*�v�4�AX��+�?��w�t?���'����v
D#d���g�yF�=;Ⱥ��@�S�p+�O��. 8I�1U��𤗼��Y[���#��|	�y-����〞���u����b��F�_X�I��AȠ�8YpTf�B�E�~��Dv���:�8y�Q��ع�G��3J��F��&9�m��s�χP���l��
���V��"�N�?}�N�i�)���TF!}���%cV�D�酒�tWbDS�2��h�P�ab�h=$��n�4A��S��4�0;jy�F�0������&4C4@�X�i���%���J��Ǩ�-7�
� Gq�҃�-X��zŃ��z���\��7��\d��YRJ��3VbGV�_'��5�k�g�">���I�i�w�,����\��I��xʲ��#�;:�H/�;�o�޶u��k~��7�����V&[\N�c�d����LŜ���BO�3��m�V����m�,�[��(-��e�87���j*��F̀ ��W���N-���[S;ۋ.�A���]�f~6(?G��Ń�^+[�T
N���;���`���Q��f��^1��YI����Y��$4�6�E��`�Kѣ z�c�Wq��tiKS������(�F�Ov&�ɐ����'*zV�Er�Z����� `F��\M���ty�,z�{-2x��}����i{9�T�ߑ(cĆz]�A�׍�P��!�i�;�?!�1�#f�2G�Kr���u���a�[x�mN��h�������`$Ic�E]_O�����5�sJ��\�����Jə6�x��j���},,�[q9ϳ7�������Xk�O0��	�O=����	1��KDzC*CA!1D��O!�'1��������r����rd��l��ՉX�yO��I�iD�\���7�#�n���ዌ�ƕ��6�0�O��1�E��~�5e�L�%�f��ޛô�U��O�VQ5��J�����͹��U�K�Xi�oЬvZ���@��љ�����T���U����k	M��o��!TXH�-����9#Kv��d���]�}5.���y�a/��-�%�,���U��%�#���>�7 ��y�Ɉ�N�O7Dxu�D̍,�\��L�{dZ�6�ʝ�%>�L�Yg@Yy�.r��H�{a��}��������d]���L���+�M�/�/6H�1���;�`��d� 45�G\!K�/���m�NOr��3G%1!���T%��%�sPEMr&}a9s�y�QEK�7�߾����^��{�[�u��/]C^{�wI��
2{�N[��G�;�����jR��������y�"��hA��o����"�^�G���S�&�8���>L��9�-�M���#�	��Cj�AHͰ�f �zs�+,�"���J��R��3.�z���]d�	��=´�{��WP�}C���=v�����<ZH׆&�73ͦFQ+�: H��a�[���D�{Bۛs޽<�7O��$Y��`��M1��Q����n���,�y��W0�H`?�K�8�Xn�h��?��et%��k,Q��+�WǌSީ�Ơ<�?!��U%���k�\�����<#��0�zk�#���ƌ������^O�h#�UA��^'���d���U{)�2j{���1����0�`��f��"�hɝ2��aNb{�_;�QLQH߲8���8(�)l�s�J�7zi�p3r�	���8���5��-��{�����|��G���y2���Z�ů��f��+�6�n@lr�k]?g�P��I�V �P�������-�J��]��uR�P?�����w��d����Ю�2���&�A�!��)�;�}����nߴ��}�΋�X���H��?��������`�<�|�w�U�A��Y3T��f�jf��mJKD�aaW)��)Z� Voވ`��s�¿gQE��F�U���`z�"W|������B���	Z��6n
���'�'�kGWIcث$ݏt�k�W'��K�1�uN .�f�_���+v;{��5J]O�ظA,�XW�5���b�(q�7��5�`���㧤��P C�Nh�4-��X�'crl(X t����.&��5�Ͳ�)f\��,���גc�S��E�o�.��w��o�a�ؠ��g"j�jp��o�*ѩ1Rh���XAXK��0� Q6�UO�©I�e���i/wɸ���ꨓ/�_���8��P��R���A�D)�Q=]�l�U
�h�7�s�16�& ���{S =M@�/x
�����>xN���ѫ�S�u��˷v�T�>�@���l��|���;�z@��/�~WK�b=���J��ޔ��h�c��l��'v:�3�I�=�	 �8��ӱ6Nm�\>DV��P����D�5�CǬ����Z����;��K�T���v�۷�?�����U�[�C�d�`6���ǤZ��e=��f�PJ���`��,�D��V����y
�ym+�᱉
;P��*�6/W�S����)�{F�Q�R��<�J$\�Enn^�9��{O!�ͱ.�[��uȐ(*�����Q��m0�~�C�oxXL%�NCu
�$d*���e�������I�=��{Aq��y֧�d�Uɋ�Xy�]�O1���N(��4��V�m��`�z�o�e��=74`:F��\�X\{��Ƕ�r
��U_�B�z�	��I����ܥ�T��9��x��oP��c�
�����)��4�ӿ�Lb�׫n�.����R�������sq�H9�r�x���Z��x��K,���<Ժ�[�b3� �sc_б�Ө��(Ɣ�ɺxBat}-�	-,�E��5\��̍�J�s���<H��h�(�E߷�X�ԭN�F:���u1�̿�6���^Gկ�eG�2�2�I��MX���x��fv�e��i�9ͼł�%�4sjD��|\�R~�4C�?c*~3���a�OX+`P��j�4-D�������{xce� 7�2i��=�\"���j�����0J���☸c(�� H��\��A�y��Y��{t�N9ő�<���l�1p:��\����m\����ܲ$?��*9�R������DK2��
���F�����gi�7b�@~��sc�ޟ��Ȯ��y��2 c�H$Ji�����r�}��t~�5>����7e�%�9֭�3�U�&�-�VA#A���ę��v�<��ʉ��R7g&���$�$�ԋ-FӁ��a���?�q樸�Ο�3��ڮ��b"�!�]�E^��@�JF�khu,u��~97x�f�ʕj�~{/�p��<ȇ-�L�8%��Ǫ�g x�a�MĐ:	x��
�+`w	�9�
!�9����9��T_b'�a��%1��VYأ�_��c1�@*��R�V���>EF_�9C�e�(#�2x�?{���J@\�M�`MNv�w�(R��T4�l�����)�Pςx�T��h�R~�?6x�t�vNPթE�ř�\7�S�65��]=[�.AX�"9E"ʎ�.�l��6�2^�P�q��Z/�{��ɚ���<�o��Z����ѧ�r�0'tQ��Eo�T��[rb�����Q�gǌ���D��|�1"���O�d�����	�|t�s$���8X����N�G��n5J���I&ݨC�I��1:�	^�=��gIe��7Ja0�ԯ�'�.c�&K� ����P��}'^Q��!���җ�L��#ˁ�O���5��c�<�W%t��y��>~Kg;)��j�l�+��u�*ؔ��~ȻiS�k0u~a���o#J/�W?J��.7�H�&U{0<le�������*�]��m�.9D~��xp�r#�3Op:�U��O�յ2@���~���3���i�R����<��#5]k����6ouD�!�%-^_�`�:��R��b�貉K&?�'�,p*	�-A���K{M������w���U���WoBm~޵���pjN����\k�xH;��5��  �z]�5`K���Wn*z!�� ���Ⱦ�Q͸:� ��d�p{\n�E=��>2����6Ui8�|��"|y~�ݻoO]c�w���J�
��!������6�b��vL|& ��N��x��y���� >:�䛋�;A	�,�ي��:��;=�=�*���}9Ғŏ�M\H����*�L�D9���cV�uܲEQ��j��e��%Su��\�(�'�3�C"F�p��72��c�O ��h썕��=C��Q{P-5��'�$��K�;
5�%Y3|�K�e�����V���D�ڲ}��~ܟ��A�;?����(���.W�lDs���J�&���Б��c%_'�i]JM}�;�A�l��1�54��>3�v�ePn��G���(��TKddt�Xl�"x�G{�
*yҝ@�(�'�$�$w�p�j��>!v�k��߾��Ȍ/9�J|����R�DB�{��%k���WC���{#x����]IK���y�GCݽ�A8o�3,ˏ��N�#Q!VD�ͳ� p����7����Мc�4zk���ލ5�Fp��B��k�F����+�L�Z1�VG�����p�j��o+-��hВRfɺ
0�����x+�m�đ�f���v���-�����V)%��l.�l+����q�~C�B���+�av����iT���!�;äb۲<N��
��l�� O���)�a^R�m��	�:�׆���j0`�NhB�*���&:�;�;�O�]Z7?�SV�}�qf� xՀlζ�N���iW9�m�|hNf�eK���D�}t\0��y��囩SJ�UJ
��������U�jg����:'�J�����9�ʺ������a� �k�,��"�'l ��I�u�s*A��,��U��^��G�㏌2l�z�E��=�M/�Ğ��m0"|x�H.z� 8��mnv���G~�TV��m���0���&D�Ċ%��Q,:R�����}�f����Fw�w�G���7&���
ԈE�3.��_�@C�ߌ����ǕTS�E	@Zk��y%�yu���,V�r^!xي�!4��?	w����|]T��ZEm���~g�����%v8�ء��r�ޙ$��0va�>	�A�R���ҟL�ѐgb�̢lp��_��oMM�멡�`N7?t�9�Z����W3���4ŞM_a�N�s5�ޣ5 �$��S��D�`���fqdm�����E�1�3�J�>	�i�օxw�C���;2�v��ܴ��/�lO ��8��z�J�*�� �r�{�Q��T�p�	ǯ�O����?�W&8my���Z ~�.E{�Pu>mA�"f�fb�Wh��p Q<ǋ�5fP���q����Z�����m�*������^�B�����u��,|��$��\i�_�No�Gf�K�Ԡ��Qs��xN�O^h�=<�������Bn�fl�I��c�15�m���綺#�e�*�q�H��x��x<A�>�oc$AR��;�[r	+t(����ǒ*�����K�J���{�i>.����8��Q��JC�-��k�x���6A�~�t*�V��-C�cr����#?���~D��*�B[,����u�������(m�b�}�Yռ#���EvJ{�g���3g�,�ptDۊ<��E^c��N�g"�ԴXBH������h����u�ITaS4��$VA��x���;�b�o�n��~������(�+3�a#��N�r(�U	GD�M��G/�r�$-��	�a��v�=�Y1a�\L���˦X9��Փ��ƴEaܱ�H���fQ����Lf�^yVz����u�Y��b8�Q9B�A%�r`?Q�XL�C��,��^���T"rv��9~�D:�����8�Dt׹jY�u���#>k���a����&�`?��������: �'��r<q-B�@K�gY��Q4d��SM]_?A�,{���:�y�`��Sa�����/��ƚ����cYJ�_�h��,�9���H=�c���XQ����)v�~�P&Ğ�Re4��]������7�Io0�n�:�p�=���,3@�u��_�S�M�1Qa�r��%&uь5O�����N7��O�f��MŚ�ˍ�����{RB�n7Q�@;RL>��]�X]q��� �C�92[�H��lQ[�����ǘ:� j�-'%������<AP��F�����(q��¢�YF���:��t��ɳ��&=k�c��` BG_L�b/e���&���t�!YC@f����FY�h��F�op��I9���pi? �T8���ش9�����7܀*{N����RTk�s�m[h[̫/�$�i�����(��3�nc��>6i��^�.��\_Y.~�d���H����@T�i:3jo�Cs�a� SIҐ�r4���g����)�h�,w��:Xd�)�:��\���5��Z�>�CGH�զH���0D@T3w�~�Ќ��=��R)���Dq�N��X2ج�[ZW��-�Y�{�chF��;ȩ��p̱���
p�Z�Y-bN�H����/��cKn�ۊyom���gp���PlC
��z4lIw���󍍮�3[v�m�D�i)U���S�VzӰ	f��sL��t���i���̎��@R�b�2�М�z�W8r2���� ���U_Ի�Q�d�H��wB|�< � �$��6/ȹ�љ<�+3<�~��H���B���77F��P�/ƏZ�#�N��J�-[���XɃ��s*������P��}�+q3\L��,1c�ER�J��b[<�o��3�s��x�AVʹK��H�-F;��7��_���[�љ�n$�6���_)�Pb�Y�tS�/P��_|#`��:���V4�:8p;�<�'b��pOö�t�߾	й ��6�O_��}H`�;��1y��E�5[�E�o_����E�D�ٹ掵)�JO|�rX"w��>:��uZ�����z��^q̐�ާ1�)4,|j�^�Z�N�h]�z2�ߚ��G����s�(l*�<��1��P��(S/T�聡Pp���XwL���A�_?��A�NT&�NcB�";"3��(-U�����cU��צ�/�h�,_bw�ղmm��L��*:$*{L�h�I�P|��P���/�^&���j�!�V�i�3�!��\�}|x
7�o�!�Ɩ��ݤ��:��� ���gTGک{����EU�F)N���/���9�q�q�ȉ��G�Y�^ �f��n�ҹ�/�FBW`.�f�i��X6'C�����9ק;7�f��V��7��	�y�J��dӆ���ΛN.��P���A���<�
�<��Q��#|�:��F�n���7�~�t����*��S{�o�Px��i�(�#4軹�tO�<�.W<��|�ɚ�>�*�� '���t_��A鿶y��v�|3"~#����}G~R�qq������挢��QA�$�#˿�Xɣ�H-ͣp.���L?���`.$���^��|X|5{�^p�`��_��Q'W!�|�U����"Fի�G���{ߏ������8�J��ᴁl�ԃ��t@(.�zn�CR���JXJ�����Zُ+�l�zbRx�ppw�}��,b"�@�U�t:�*ߔt�~��p�"�$��������X��k�[ס�KIbG� �p��)h�&��tv�h�5�h-ܔ�^���{B�?��	�^oݯ��R���������փգ�T?w�*�Z΍1��b�2l9�4*�)�!��܄r��΂R�X�`�N�m-�q�,�HYcn�j���X�yJϬ/a��ъ��
_���gwÍ,.g���"�R��܋�l8�����=��x{�i�e=�����˞nWΔE�����2�Y`Pv4�B>U��5��P�������.�[�ė�ȈJԏ����I�\��Q�%���}�y�,����8C�pC7*�q<]M���]�	�i����Y%��P���3L���V�DJMV���rw�>� ċ�C��o�:�/
��K픝Rf���Y#�:���e�̓�B��T��&���1$���s�AXԧu��UX�Y�/���F����i���z嚌"՞K�:����Z*G�H1�D�
�=��X��m�̠�531�dџ^,z2�Ȣ��o����X�# 9�+;)��m�)9G��(v�=a��i�YC+�Ͷu���E�L�ؒU����?���'[�{�_�^ �NS*pe�e�єz�����f�kR;9�%��-*ڔZ����ǵJ�p����e��P�ӹ�u5��򇽍��Q��e"uǨx�&�c��O���z�T�Wd�ngMWS�!��钑؀h�":��JA�v�	���.� ��%Cw�%�p)x�=��5?�q�(m�x�t?�\fV�4	q����Z2V��l�B�������_��H!'���s��6�+m����l�{(W.>s�����(a�n&�5�/bB�؈mb!��֮�V�߹��y��><@}Lr/�.���t�����Ň8���ڬmln�{��4ްe`��8�9A��`��Ͱ�	�#Π-��q\I->�J�����?AM�j&s+x�?'���9C�G�{%��"�ߌ��B8�27[��V?xՔ��<k��������_n!ԓ[.��Z?�o��)pq.��g`Qum�V����d�ɵ��T�
�}Z���i�|�W��I���Q�x��iJ/o��F���a
�#]~�5�~��h�"5��u1/�l[9�R��L�q잵��w�&AUC3�&%��&$=)�XG͙�թ"tf�,Z�������U��zv�l�����-HZr����^�<��|qPm�c��8h%N� ��6��ި	�?� whV��1��T�FXЪ~�7d���#�6���W�ZP���7�Q��]%��:t)�b�
�
n#qv��᨟{����������h'�ãx�:1ښi�gn&$�0q�9�s��Y��1'ࡔU#�7m��`J �eѶ��IğqPV�.շ7�o�.���gmj���&��[��P��$(��?�l�p���~�}���L�P�6��Pb�P��N?�~��j��D`jzs��'���v�.��O}�R���6Ds ��}�>,���$m]��� �;���{_c\l��J*��zߣX��];�k�ZZ������l���>}沇=��1O7[Ɛ���n�`�W����`Ĥ@�B���U!)�lvK�{�pu�'�3�5��	b�Zeu�$�/=f�ȫw�.O���:���k�y�=z�:}�=٭���gx��^)�x�oH�	Y\�28o��V')�*3zE�H��V�R�$F.� 	���A����sek��KM�8Y��4V����
ep��^P��
25,�Ol�A;R�?����D���?������`��v�!o�o�;:Ví_�_��c�b��؛|�}�����{'�M4 [��e�/Hݣ����r�l0Fb��*d�t�-� \��[�����ɇ�7�%���Gy��1�܏ڏ���c�i
jM$���@$�u���k3��c��#T������BYpOdd���k�O��WS�� ��_U'i���?d�M������D0<�'e�
!�:��&��w�}��� �V&"?ńs(2�j���(6bN^�T�����{���t�����/�-�9�g=�r��IOf �i"aY��m+�R*]u�%�\��c�%J3�����<f�t�*�}O�b�'�-���3�S*Ý<R��yx���i[(�N�УU�������\nD��9bYÐ�ߗ�B���8�8x��F�en�5)�s'A����.���vuap�(߃�/^/1+����KU��������/�jS���+�o�7'�#�FG9�{7�e;�:�>U(<��{w�������*�!7�{�Q5��Eە�r� N7�쵲�����-Nd1s�!�D~�:|z�ǂ���#
����tf��z���&�*��ǂ?��T[�CK�u�pN���]�0Y!�^��ȹ�eѤ�T�uԝ�b��3�]�]����U��U��ڑ��b���I���r�׾X�����)oQ��hrF�g���'4�٦rPj̞���?��P$�f;��Z ��u_���T�ә�q���i��W�r�+�Q|�
����T�H�vG�ua��u"
��[�_��H�(�"��,.��f��Bw�>*ƈ9]t�M�n��,�f�S|����N�(�*�O���m=K��%�N�T���2/�y^�^���FԹ�	���d1���ާ�/S.�q��� �8�Ň:�������R��N�,s���BU^�� l��հ.��^���<�n�|U����팷�q�>i<s��K���R;*�7:���/�����=�B5�c�_��8��>�XX�M�܌��N8�~vYq�1�C�]my%��9Wҕ+�\���Ir��M�-v�q�̀p����!aN�R��&	}��� �A��� ��$e��ZIQ/�8c��^��4��%C�rL����Ɉ%�=�K�ض��6�!�Kw#���+����^>�p*UtPBe�Ҁ=�  ���y�!�ð3��,̌��l��q�-Q�ơ��CޅPI�b�a�� <�V�	+5۫���^%��X?]��������k �t��:�	�dS��g���*��lm��4�H
�E��	���$��J}�J�5k�-#�z���c|p�}=d&Jb����S1sxD��	��t���閱����6�ط��M�+hc3�Ϟ�|�+ьy5E����\QA)n��8S.s@�x�M�*mI�M�U�������+��os�O'�@���y�.p��]����g^�m�j�dT�'_+t���aQF,��]����XF��^�㣗2����]�q�������+���w�T����b��$A����Y�4���g���ς�xJ������
�6���N�-8���������o��P�/7S2\2'.�!�r����5'a1�iCJ�]M���@�o���X����'˟�_l yB+��ޣ����Y㤯Cub��_�±}�#�.�Wi��'[i�S_�5�I�����cC<@�P���&LL�ʐ�~�i���l��P��Ȅ�D�T���6�l���!�9vG`:��J7��6���^SAv��c��	$�nf�ȃ�_� �I�:n�hH��O6�CȰ?!������u6�fkK0�c�<?�$���f��t��3�P(+.���5g��d�!��&� T��,c�h����0��@T󟣄�YBӦ��f��x�bP����UNL9�����4�B�,�M�Y��Ƀ�a׳��
M�.�C�0E'���a��H��K���%�+E��A7��N��͵�bJ�>sww
ƩJ�q=��������6m�L����6��5N$�ƉzvcVQ�R�f�*+t�ZG�~�G�BEdzg{��t��¬�~ʻ3��ӄ�!�u`M����+�F�~�ɻ��~;��ʶvɜ&ȱ�ױk�ј�֖�w]C�)�����t�4Yٳ�$R�%��v��Y!UR�s��K�D�E�@x�d��oa��v�l��r��Q
<t��9�4��:+��|����`j�S��gb��w���5��4L�ty�kp��c��;�E�O����E����&��
��'�pUܕEU�����&^� ��(rY�9qy��4p�K��t.�D�䖠n����ī"D7�OݭPɌZ!-)h��~���M\e�.?�WC����]I����2w�\	�	��v=4C�Mf*�e$�ȓ�q�MV����N-E+�I��Ѝ�u���t4-�fX}�����r�׺�����B&���i�O��ש���L�_?D[:Ɉ��	:�(���
�MJU�}&�Ր��U�n��M��bLU�c�ϭ2ù9@;�=PF��=<�.���Y�6c��w�u�Y�o��]sU.t��<��W�w�Cv��n	�`@����A�|R��ךkӳ�-�?!�}�i������f����ذ���"92�\�9����
̢� XB�2[�����Nj�c���R䕕�"��+��U�<��DR8TB���Z�����B���Zf�Y���C6���ڎ�۸Ǿ��W5_���-��<73�J�NN���^�\�i X(=@-Rvy�o�$#����5w�nNF�j�B� &ؓD�m���5������ا�s�e���{�k��̧�
�����%�n�~d����I�^`����"SDE�8�d�M��f��9ddo��1Se}��XK]?�9(D�ş����5�[m *b�l��yJf�)����:��L&��Q"Py��k\������t�gQ^���Kk�mq��\R����c<��X�l��S�3���Y��1�L�_���,�Y��~�T�Ԫ�k�N�R���a� Z����.=̵xK�̨����k�C���}ܦ��K��T����8+�U�V��v�);�4̀�S�hW���W��\��R���ZW-�PZSYw��7IF�BK�3�f;�R�(���5��=Q��~ܠ�6܎�RN\�o������1����b�Ｇz4�9&��羜�@ִD<ssy�-*���n���V��Q^��������K��L�� -����fע��e��>b���&O��c��$��	��_O��!R���ox��ġ�S�a���f�#*�u�����"�O���"�p|��w9����m�#8��<�����+��ym ���rc'e�1��ӴA�W�K`��:"����B�+E�م��t�{�:�9�e�+�!���t�c������:�7;�o�����mt�n^n�:�/Axnwd���Ì.�}�r��~��h���4���֙�77Z�ſ���c��Ix�2zc�7�ζ����v`��HT������mw)d>:�����V��n=����))j��m��\�o�4��ZP��00"\㟳pS�1��L�8yO?�Mr_����a`�A8g(S�'�j=���r��� �p�~(�GнWd���'���H}�%������ z�)l� y��@(J�h�\��C��ǟ >�[��Ku�:��Z�s��[i��^�����سJ�4Y���<Rk�hL`���e=*a�L������o B�wcx�]��Y�9������N ��j�����4��3%����v}�'�������v WUF�ۅ���A���K��/�����:�p/����R;�����=�p����b�,�sVS�������7���=��^�A�k�/��������]U��@�΀G:`+l���q%�c�%�)nɬoFf=��µ��.+6|jCS��c}�|�q"^H��<�~5D��6��C��й)d#�9�F�G�A&��X\dc#����V~Ｏ�Q�)dsɄ;�(��n/Z=�[���<o뾑����q
� �]��`�Ż��0rF�.�7S���H~v��T�2wRN%҇Σ�^�I�A���rf��(	4�K����E�� �uv�����,P�Ǉ�1.r\�����R���ά !/���i(/��
O�i��!����a��g�JA��3�W�R'��^�y��JA�DnH�Z�8�3����qH{ŇV�"�-�>�8{d��ڤ�I��M���!�hݧx9�CG��]:�˧�@������Ef����HR�r7��J�O�Ҍ�G+f1*'�Q,��f���#|�6�3���>Ӗ��/�����9�E1N[&�1MR��5�����7��t@̶=C`���J)���[*�ߤ�&�U��m{��>����:�B�h�9�^$	
o���V�uP}E-���%�����c���<K+�����G4�D:�W���Hr�J�[��<�����7�-��
\-��.��I�'��"9�;bf����S��}2?�	�R�IX�D�����XiF�h�rvH��l814Do��#U�	���A>���:��NtO�٘E�U�'3WR��q�I�m��rcم�_
���T?S���2�;�M���EAz:0(A`�9��8 ��(�yQ}/�`<�Ӓ_u
��M����%��A4�s���|}�	w��a��.4�t2���᪴��67A�؎�AT⽽ʔ��+n#����-p��@Δ�G�-�i��|E�O���s���_ʲ�}�"�S��v}I:i=(y�7����7��%��+�W9(�w���o�L �a4]�����7��́�6���Â�юgZ�F�.��)5()ԅ!��I�w��3�;]k�k�m���T�r�*yQpi� ��J��f��:>ukY��Z� =m���͢�y箶h}�|۬���Ί#cGo���pY���s��K��n��S~4�"_��O9��C��Pn˼���pH)�S�|qu�dW+�v=S��])��Dgp~�9n}�G��࿐C%��S+z1��µ% �$�{|LPY�x��D��\����qd����j�ױY�|�&)��U�v��5��9���e>[iX#����ʰ��O�<���36b�`[�F��~���@5�����tO�Hޤ߬��T%7� |�	��J�a{���Vs\���m'GV&���w��2�i��
~2=)pQSL)c��Z*�3`�R4a����M�����*����c	$N�-�@�˹,�Ʒ��'��v���t["7Dq��x�Y]?:�[�*�)���t�z7�2�=��q�s�Q9�}�0�o�}>�{�؅�{i>Bx�P�RX	�DRG�Р�n���tg���K-�.\2f4�:ӣ��f]�.�ޮxl��%��k+sX��*��n���^j-m�M�D�?�#��5�Z�}! Rߋ%��13�D��Sߦ�a�'V� ��k��if�Y�pBP��?�Ż��i<>����x��Ie��L�����s���,J�,���n�?�7馄^� "z2Y!QSHM��_"�<�_�Qz��pbZb��`���guP����6.�8x^���z�"��a����3��'{N�F]5u+6��(�B��	��5���d�j�ї���fM����.?�*�) +�4F��������_"�۹�����e5
"6�i�"���(�\�V:ধH�J���Ȩ�pK!xW�GhD�8�^�{>�-fM���QY\�������uނ�����RV"z>6,Kn_���'�ݱV9[o�N��@��V����u:��~Lhڢ�?�9�W�ž�5ᘯ�d���6r��Aŷz�65\e�9�VASt!���x���C��H�@-�7si�+�C(~���f能�߮%i��U�X���ZtT�&a�R�g��kѫH�m�s=������������ U��FO/Z��~XFw��U ����I���T��LO%Ս�B�阘�dv3�Σ����Vm�%N��)��r�"H��N��ˡ9w&T5�����E#��g7�e](�CG�C�.VG���U�g�]�z��R�%!��@�.(˴���P�o�,�V�����rZ0Ow������f�K|��I*ߢ����h]��B.���n"�>���c�������JDقo�{�5�7H
�h��L� FN4lV��2��s�L�f9���:V�b@�E�g�B���4�<��HS��3K˳��Ӈ��It�r�J�Mڜ��F��䮕-"|-���C�f�ڮ_ϊj��n�3���-sX��'���S�p��F�iI�R����e��=�pq�{(G�7$v�h�{�_<�Pܜ&��|�*�:��8�06?�bTYs�E'6�vX�B�#�}�Jnk a��.���� � �F� ه���gm���<��-�f�+Q}��f���9h@;xw���L�5#�ꌦ亐Ue��P{n���~>�n�m^#hRh��#��r�I���}��4�c(����m�h���H׫�v1�
x0�λ�����|����h"�LZ�����̮����Vx��&��E�,��lz8��23{]��t��������o��	���7��]���!��;�_��u�	��/GO�����נ$��!�P�(S��T�Ǳ:�@]R�����`ݳ9�]���n+�&�Id=�GPxC��\@z��)�Ғ�h�)��y�B���Q�@6�?vX��J�Q�U~Z��ؤ��C��C��`aT����/Al�JYA��W�J����J�>���x�'�T3T�G�?Fw[�I����9�?�CPA�W��@L�͗��='ǲ�΄��7T�b����Y{Ȫ�x����ýֻ8�ݪ�<�LjZ&���j��y�>�>9Sc�)�Ӿ��ed,��1	 �0s^�Z{Ւ�T[�c����^f�1��|m�7��O��l��%��|-�{��6@I�)����������u�&#`G����x~f�|x��m�&[��Lz��o���V9����lm��� ��չDk�Vr]J ���{�y:�S�����iT�\IruLA�nS/�E-o�_��"�lf�J�	R�.^f�c������Ӛ�8��FT"�%)���A��p+�Ƙ�i�P��LN�BR��Y��q�p��Cp�҅F��5�+\P&�U�N&Q�Z�o���ߣ�!z���^0�`5Kr����[:�� ���	� ^��n�Ԛ7��/�4623��S4��@���#\��r���
�b�'�,x¾Cü~Թ�d�~$�������@�\�4ʒ�Zt��s�J�:K�zoll����#��;5�FLp0^w��#ۻSz�z�WB^T��S��G�����v�±L�X��������\L��# gZW�T�V�n���������6/j���r�~u��s{�o��e�,��`Fr�i�����`Õ�9���|7�ُ��"}�:j�ig��A� �zy1aT�&A�q��P9���t4����S�ǘ5v[iE�T�n���;����߄G��z\���t����8��Ǯ{�}���2�oX���Q�:��);9����m�瞜�����t|�Ь�8�Ig�J8M�i�`����ǅm�5sR[���>�+��v�nD�=�s�8X��f^]��6.;�sQC,D�~A�����7ɑ��W�Ru �mT��a5���Q�lpK���u�7�O������涁F7l·ױ��1Jb.��k��X�5m,��_���q�v��~�Uǫ�Y�ɢI���/p
hA9�B<y��/5���f7sD�z�g%�7��yu ��-�$U�O�d��0�}oqMy�TH�+�TX�F���Ϥ��V:8#��(ȑ�h�7���]�}�C��柱a�k]}]�9�NE���c�S�!�t5.�Tia��}u���S\�M�ݮ��\�@�1�btś�� ��]�I��� 0�}3���P�uo��8'��iư��T���9Ux����`�75�g�V�0d�!��~ő�"�E_�ф�����"�8l~�-�9k�z���Oa��r^24��y�5�Ζ�~u�4�ݬ��}��*���Zo����Y�D�.�F+�N^Ȑ��PU�'�_Gt�{M�O�i�]�=�p �ZL�ϯ�E���GU��x����d\�duW��4�s�7Ф�����}�t
F���E�s3���r��4�Sf�*�^���O:�q�Q�+�,��g�-Xi����o��3��i���K�q����
x�z��[喋p�Ћ�8�Ŝ��)���+N�A�BϬ�Cf��'׈���&C��0�SGZ�۫%��40tC83��Kњɓ��I2Q�b���WRP��]�}�!
m����<�@�2���(��GP���.|���:OV�x��92�~8��=�>ʣ	��L��W�<jZ���C����z�<aXBCsi�D�`z�/<d6��mS{��՘?���a_7jKY�����_�'
���Ic��`�"c-IҰ	F�Fl�����2������$u�%f��o�%q.ݿ�X��cMo�q��nA!���5:��d��$��O\�D�Fa���`�`%Uk�HX����T�8hdq����7�6�uӮ�:�b�446��HufK]�vrݕ�����;��`R�3��p;V�!c�t�̐lz�YN5���5�s�53��|{��*��3ה�G�=����X�f}I*��90jg��J�I���CTt,N��x��'�\��%(�6����
��b;�I�,����5�Yuj�|�:�	�������[�!��`,�W�s�7 '4�cD�q��J��;�a�Ɉ�X������O7;Y∏n�O����=\��W��Z-M�E��v'�f�ٍFE<�_������[1��8��0�v�	"�&��5>��<�_Jn��S�aĨF���I���tD#_Y�o�~5�Э@�2%FCP��pΰ����j�p������k:�޴+3ȍ�(O�abƯ�1]g�ֿ�����<V}��N���:�d.uI�x/~�m��,j��u3A�R����/�ȴ�Q
��o������G�3b��2�^�W%�������a��{�S`m��	�	��5��j�aA`���� ����R�_خ��J-��X����};���r�{f4��Vfu����i}P�H�WS��dMjK�l:��Jy�-���E�����oJR_�P�w��.�����R�����&�����ʨ�fr�vY��7B^���O�L^ϡ
�	��.ѱ�?��2������}��cў'�-�����a:�KG&��7]��n�ׁ��T�YqTȞmi.�jD��7.�!#天���F��F�Z1`ʲG��iBP�[��XS'	޾k�9���ѳ �tOO����ۧ/�_���G�cBV���e��{]8A�/�m!����OV�� �`E�7ez7w�I�;Rj�*>��@W�p�o�c����y���ȣ\��>��� "�.]w���|�9��J�a�TV�0����y. 7o��2��_���4�!�Z�q��X#m*A��<�n�����gn�~�}c˰{d҆P���'^I�L����Ηqy]RN󣡝�3�B[��YOR�F���ð�Sj3���G\� u�p�S�^/kM��}A��ɒ;WS��������cNd6a����8@E�ӊz`]��q�~�S�
�j�cR��8:z����7����%ˉk��<(����:�Jq�Z亜+��:=������_q�z��!�&�k<P@���e�3u�H�O��#4����&�J�N iU*\5�>�[� �`���Ŝ��� ���y[�)p�~Õy���1ڑ�#ua~�球�B������Dc|$�8ܡΒV�kO��z"�e�����Y�6^�(�X:�����<@=��J��f��p�Y� [���3|��ϑ����d��UP����y�e����tѱ�BQ^]FW�;���O���߬~��^��EUi��I$1�R�0�g�~�1����I6�� �W0�?R�8��7y��!����R���/�DX�/�-��$�hs��7g���Z$&a���3�4��HƩ��5��)�.�j��;�CI�(�a[���d���+��`��&���(��I5@^�����ז$�4B:���9KDTǫ��)�L��`��X��|�h"�^���P�d�lWS+>oX�{7^'�����N�x�O���� V�݌*m�R*;������VZ#*�,>��	��9��w v��q��������i��nģ�D���6K��	�I�}b���{/l��5�չa;Ҿ�PL����gM��z��PN�-|5��6�t5d���K�ن��W��B�׊��:,�% aq�7ƺ���P���3�L�7(��GN@���f������&B���c������=�UћR��y�1	�*��5�*�Yhk��-z-���x��:�`(V}�&��>���=%�+2��N���j�0>ܼ���ᵉo?�5u#���Pb�I�� ���o���7������O�-@��^�P�ѳ�);��Fm>+X攽��ċ�X� U42�f$��H���G	�3���i����X�\�P�8��Xp�e���������K>FG�	��V��s�f,j�ٚ�����U������(>�4h)wi`�Ji�}=�{nM�=���G
��]i�1RN��T~E�.^�v��s���d�&j�Y��9u��B�l�Pѣ��l�V�\[���X��O���C충�}�\XrȄl�cW5�|�b�9���AJqz��%������kgtӦP�dS#�=�f�j*�����j_�;�(Ǌ�]� ��uH�l�p��5'����4�����������%�M�y>ޑ5�n25e�aM�FM����������9�؎�5z]�����iA�{*u��
0��Г�u�-.���L��񃾖[ȹ��1������f���XZ��R��gr��I:H(1X~G�eS�-�F޳�����I�Z����g;����y
^'�,̦��g�0TF�#��_��%]JMJ�_�,��ci-K$Q�b��4��Xu���"쳴jp8�jO���(�{����+ù��λ{Cw�Ы9�W>1� �%�j79�;�u�jSYS��Qt�{/g��+����Η���� 3��"R�u���'jX,_���L}C�Y�\X�&��O�J,��|��O�f���7��$Qs�5M�v{5��eR%��	�sv�_1�4%;��в���	؂˅_��;jvT(�UwҘ���&x��WBE��o�D`&@� ��+rVu%O���Y�G�PKh�TU:�~h�x���hs�Ǽ��)!�|^�|��	ﾋ� �Tz�I� ����x&��Ե��uQ�ƧO��+6����9"ѡ�RL(qo�z��0�93��@\����O�PJ��r$��n~e�/���[ �H��>D=(|�l/���:������"uA�/[����ZG�6#n{�ӱ����!W� S�G�� �R�dv��Hp�0�*��zG$���j���}�����0�綪v�ʀ�Mb�r���p�S���y�Y���Ձ�sI֔�B�a�T%��|��x��N��Z[5y��6:۶3y�������\�4�"��hs(�B�1M9��Ժ�\�o�מ��ȹ�<:�Ɇ*
�Ỗ��o����;�l>3�_>E�ĊZ�R��\�����Cq���J
"�
�b�t��&��p�����+�$�p��en:@_�r Wy��l���"<�C���2���������w~��,�[%����H�l5hz
0Q�s�<��;iL<����R�7ƒ\��k<��ͽ#OTU�vQ +�_�KF�ݬ�¢�����[��p��uK\��;��q��7��E�`���]�,V˗��JU�#�3����
.���k)@�r��N�<zծ�m���k혔z�3
�5��IԜn��<u��d�:��ޓ�^��n0{���a�r�VMI�����,���D5��){V �
��a�)1B_W�(I��(+8N���c;�\z��. Q'���5sY�"�H�sUu�4��L ^��z���5v���1\���k��N�3΋đ��%�.u�g���;Mz������Z#�2cĶzI�,ߎ�Ķػ;Gn��N��=@i7�u�c	��yD�`#��T�-^G��p>��2y��������)�P�n�߯�cAE��~,���X
���*����%�z�Iq�G��Wx)UJkZ�97���f���1�i���C���wy��N�?�ez��AY���}��ݢ�MyބM��"��#���<ҁ
n�t��S�6j�(��U��ۃ4w��r�?�g����o�K4t��=��BLE�������2�e�0��?�߱w#x
8Ch��0�Xfa���$����TM�:�l�ϤF����Ij��,)���lH�c,-]1��@�$#��J����*�n��%t1G � ~A�{k�������ZqtG�&d��S�k�:�A�րox�������\���|K����,��3{(eq �)e,�~ڈ
9L�t(~�J1U����s5����Tk��^mN�r�¾�����8 $㵋���0| QhA�7M�����H��"��
h�}��Ƕ�����/]�>�:�l�̥�8�$j�i���E��)%��>�%,Y�7���Z�҃���&qĢ�*�)���޿�dSG��UxK��z7ou�Juر�
~�A�!nNkptZ������27g�7���;��QV�fv�w;�#S�͋6tzHB�� 3y�Y9�@^i�.	�c�;Os	 +�=�Xң��?�;p(� �PF;a%e�ȴ���j���=�yB���h�3^0gT���`]�G��3K�VX<6�ȣ��֋+­�@$��n�`þq�r�������||V[ȏ���L`M����	1Ό�9r�6Q$���SQV�KV���<_�G��Y`_��g��d����\�m�!V�*���$��ǿo���R5.�:��E�*�0�d)��f�j�W,�d������ě��b���+� �%�H�x�uwXݚyM�N�g��p$I�4Od,*#سp�1��V˫�CZ����gFx�.r%�/���>/#�%Q|�^9��04�U7�n�~Ij����}ޟG�R ]����M&������(�6t�-���޼�� ܷW�D�����).��Xs�%�������8��]�u�'��nH&:`V�Ɓ��|�3?��m�{�n$EHCGPB$�l�+�~?��三���?����vT�:@3��c+��Gd���lV����uW��r�y���[�e '����I(���E'�^�N(<�/�~^��*�"�a2t&���a4÷HI����`{�]l?4y��{���n��ؠ{�:53��0��Y�n��О[ V��n������ |9 JY���= Li���Nm�pW�w�%�m����;3.��m�\�5Y".�f?��y�И�fT\a��v��#Rx�̋�C@�Y+�D�i"�<����1V�څ;&���{�݇\>��0�!�_iq���
�!?��@��j�r�O�����7�z�0?�1�T������[�[�|����߳��l�W��
�6΂||zQZs�.������`�����~e���,�NO��`K�Hy��  /��oZ2	�lN�O��I�y6$Q
[i�	���@'h-�����V�D��w�X��A_���^.2����0`kV���ߎ��sʶ x�7�M)(	�5�G\�Ռ5���Lզ��8_�r�(��p?��2>���'�]�eo=~o���f�L��(�	�N@���`�b��_1K����6���dH����y��0�U꼣!-�Ϗ	�S��р����W�>�Q��������gC<R~j�{[XM��Pj[�	9{՜\ǚ��tu���(��Q���W:���#F[�+�s��J������VBNs>Ã+_��`�|�G �E�%�G�@c����.C�Q�`NL�R/��6 f�?W����2
T}�Q����~�!!�?����7��T�y��'�8�Jt��11�j����*8EoN��+���j��N�bf?"���Ѧ)�֍�d I̾"L:��$9�Ytf�#3 \o�[�U' �|��2R�E�KsL:➍���w��țm���X/;��8.3_?��3-	�#���B.;�v��C���	�,"KY����Hy��XVѡ�E�K�&:@|�$��/�}���3�v��fR�y��(�ӷ��U�D��u����p�����U)J�9��x�ֶ��dAu_1'��aR2�s�6_4�{��T�p���S��5Kd���k�M�=h�����e0[���a�F�>�~��,���9t���V�/�"��)�t���C�3��g4H$��Z�٪�"�3��za���گ`R��|�A^f߱��U_�k3`5d�$�WJ��M�~����\�dE�#���k��}&���k��/B�*��ߟ�6w��зȦ�������N~G�iN�T��Wg������b��uk6�v+,��E�+��f1(���W(�$������ �62�� ���[+2��<}xo;����e	���CH�(�t/|nKCe>N��i��X�^Wh�|���+\6��b�5�V&َW��`s�P�S��>	m�
�O�� 2P|Ak�P=���U��aH�������ٗ�'A��F3Q�C//���
>G�=�����#<�tF�"�ý�5_ka�D�WQW]��"��HgOR�SĐ�&���Φ�v��I��^������`��??�hd��l��ۡl*� �zd�/Aq�G�`X��x�����@u�O�6���PϮ���l�"q�~b�0��~�5�v/�FWE�+L�UӧEa��ʁ����,v� ��=U�({�IqH��p�PkD&}$�w�(��f�)W�]5�վ��HL���!V�.}O�<q�b>c�i�)!�$����M+����/>��B~��2�& Ӟ�I�"M2?�edt��sZ�	�?��r�@��QJ�7����Rz8���ȁ�;D8}����c��?��b�<ijWK�}���f!�\߄�{��X��Loh�y��-��Ro���� [g���0裿�X���C�4�����%h�;��0f�<NR	ς1p?\���n�4�xx[O{��$AN}�`RE�\h������HҕK���]�g�SݐńP~0����`ރ=��5�����b$�����(�+O��6tٵ�DI�B�ec�U_α"u%8�����
��q0r�����aum��p-��SE�X������+	8볾)���]���DL�*���2�$$e���Rb�ц{}���b	R7=����Z�����7d�3����x�a�eL�K+����f�MTŔ���%M�������H�V8	���a�o�*S#D��i��
*��1V��s4��Y�0j�E��k:����T��0��^�P���� I:d�A �5w�����#����h��[�w^���-F�U-��#�Xk��K��3"v�VmF�t��+�N��J�
�r���;ĉ�.%�5����Z���lG���ӏ���(1Lx��F�f�N��.��x���Sąʒ�%��S�q��&���Vo�9���ͬ�����@����[�N>����no�����U�I�酀[�!�CM�.w�*r��M��z��cY��l�6/r��������$��\���B@_�ŧ��JMf�s��Ьf(�ݰ�G@
!��@���'�]��å�o%�\�`As"w�,�_�2��5�5?��_����g�3/KҀj*l\cf}���!���|3�:�����O�iO�] ]��viCNa�n�TR�s>ϩ��������
o\�?97�N�Wԟy��im5��:��F1���w�	�R�R�]�C��"����*�!�G�,F���B$�M?������
�-�-� .�Tl���*M�#$rR�<�������!��������$M�Rv�ļ�X�a��V]�r��OeTXgj�����i%:�r݆FL����}��4�,ٰ��0譵�,`z}�r��f����&�\����k�1x�eR׈��1e{�:��W����7�Dh.���Z3ݾ/�YZKQ��2�s��e;̐���H_z��T��>&a;�a'�����_�·j�e{%IB��N.@N�,>����)��d���A�T�'Ù�y#�����xwD�'݁@��,h��@�X�vP~ӠiK��.�IH��������������'e�L�Y�>o�"}n�y�`�r0ܤVl���k�	4}L���8U�qz�jt�+�r�FRy��q����a	��!b�]��P0���f$omJت�´.���C�=K�诱����u��>y�^��t'���ѵ�Yx�|�������dC`&N	Q��>���OVK����g}.�[!��%k��;������0.?��,�؅�̅�@�ǩ@ij�m�
J�TiF�z;�ʡ��?��><���B��(h���8����lP��i"}n�j�8~�E]�JB�?��R���_B��߭b�
����t���<\���_��&չ)H��	��؞|
�z|:���2�t�,���+��;��|eѢ΀X��Gaџs������ -8���'.����)p=��/��_Qa8žkN���`cM�";���V���8ZP�I6+�.ƅ5/e[J��n��H0�oE~+�V3��Ǉ���Y�O�l@Ԙ�N�s:�L�-LuT�܃�᭹�-[j�2�Dߛ�<�6smU��[��s.ԆV��b��D/�G���?�;с�z9W�ǩ����_fj���ds|�nT�S��.G�Yi���_�YBCzS�0��WU���'qW���6�̅�ey��lԲ͠�� �&�e�! ـ~�g���ft��	H��P��|d�*3QqPIӅ����+�������p�����':�b{h!�Z���	�g��C��C��S4f����snS���5�~�)h��*PH��vU�	s:���r�ل�d�9�Y��:��Iʣ6���������"�l
D�(Qx��%�^�rzSw܃/�d_�;4TscyN|
"g7��H�J>��ȵ�Mu� 2,G�J!Ɣ`�)�'p{�����b$'�H�u���`����Q���� �b���(q�h�6�M������0ynSz�,Q
�t���6Սj�5Df֛q�Xi��0�Z���J�XR�飊�5_3l�a;�%9#���c\���k�>�+��^ٙltCY��1�#K�.�����oĆ�A>8��#O�ؓ	�#�d��ָ�v~҂�� eRexi���)mA�x�Ž�ן�Kr?�Di���m��w���$�K�B]V�n��
�,�oz�q��tgn/C%�	�BM[2��`��o����on�t���[�j �1Ơ�z�!�^9[�s�D��Q?�2�z֨qE�����#��Kj�H�x�MRI~����#��B�US~��``/ud^��ؽ�v�%�
1Ert���\_J�TO$cS�����݀�ޟd@u[���mO^���HG�g�&��ƪ��pQ��N ,l��ym�f��q�/|Z����7v���0󎻔L?/�؄!����zhd�rHȯ	l8��e����	� 0�3��e�=�τ��v���0u�_��]���L/CJ߾d���0V��7���pX��w�����q�0�&Wv��:��2����f"��X���#�ߵ�����b����P�ǈå������{��d�Gꗴ;S��=���_�^7"��&2HR���P��Q���Np�JY�����ePE�T�s�7��^-�ۢ��8�2BߵWu�;������_�$BW�P��i*��t�4��P��^���0�����c��f��#L�辅�ؗ���,˦�: ����%�5���ϐج<����Z���Դ�f5�����ۺ�&8zF8ѵ��ʐ�z}�-�X�7t�@}���� ��zx�%aJƓ8�o��\j�XK��7C�; 5oH���%�Fq�	9y g$Q�]J��xD��C��V�Sޡs�#��ByZ�)�t��>�_�7c^�"~:z�g�a򗶥Z�����)��Pdփ}���ҟo�&%�zB���5���&b�jl�����s`�]�Č��]�>�@2�76A��΃��Ỽ*���P�$�>�EN��o��F�!�q����측Z)��V+�����9��7���р�J���7���@�� �ʘ?)|��}I�2zߙKT���[/nk��4g��?eg��S�v�S/״��a���H�J�k��F�0f����O��w-@o�{��<c�J"���R���/�N���'0u/QI|W������?�W��d-<?Na�A��� TxݖS#� 5�N%s�r��PE�51�J���?ёyڪ��e��xW�@�]o��Fo�|��sK��!R�6[y�:1�IY��R2��cנ3v�g+˒����m<m�Z�wqOQr��UŹ(�ʋ�wH�F��Ys>�H� �Ͷ�̅�'@F�"5����Ig~��|�~8��Ri����UaDI,V����<^��d=�mh���	Wm��mN�� ð���"Ҙ�vA�Q���`��tү��&��{����鷛*��ϭ+���	kD����Ut#��w'�z���o����yg=��N�G�b���5(�d=/�%�R�Vd����[%<��/mW�nIS��yO�e�Y�*o$D(�1�Ʋy���z,�%j��ï��js��ǅ�!���n~I�q@}�M}Yn�}�+I���L���)~w��K��{B�L�hs>˚�	��a˭��]#a�r<�����FEZ=�a	��hkd6M-E��5E�i�U���{v�f�H)�B�H�)�}dZ�}����pC�"w{���pL��҂������_��.�u	�������쳒]w�A	y�>zM�<al�)�b�/�~lXJ�,ny�J�Q=&�ZV��Jl;��AA��M0�<�'qpX�߭z�����X��	M^\�(�P`a"]�!�?nA0�=�K��>t��R�d!�p��4�.�����Tȳy�=t��͹N��"������|���[i�5�R�h0���(l�:�F�	n`���@�JySo�d�c�\X(KL\�鄹x�IOއRګ��R�������΋G後;��\R,�_����r��-�Q��/G+�"w�[��r��	�a�+���_U ��
���7��Q�T\���ai��,��(o�kԝ׻�F�`���A��8ʱ0w�Z�^���־���d��F0#���P��ɹ�[>�)L�	��zcA=�'�b}�:e��bi�E/�g�OK������Ś����AFz�E��nR�R����CAo�u:��N���TK1�/4�ꖫ��G+�Z�eM�_	S�.%�����g0�41~��P�#�>��o�͸� Y!ή�?z0�}e��6�4,�Z���p��GA@.�Wg(Tx;��̙� B�{t�'��8Tv��iۧ�\����{���z�?f�#���	gx0�l�#M�Kl�~d�Bwa-���:gQ͈�������;3`#�BAنᄖ�,
\�`�Ʀ�4B�����w�/3u�<���O���zz�{�%��q�ճƚ�sp
%A����������"" �W��]��
�]	S|Y(�XSdҮ�ڤ8�6��9�I#f�t��O��� z.W��)H��d�/gqƝ��J�fu����X�ి E�Y�攺)��c�����r&�0�r��nZB�H�c�G��V;�l���`�k������<m��1_�k�љ�q8�r�3��f���e�s{���Ι���&5l��գ���Z�����E5�+$-����
2��	R�>�W��ޡ7�1���:����)����H���H�6_�j8ӌ%��v�>O*���1�֠	g�zj&�eq	Z��������(b=FB|�D �(-Ɔ9sA���ZY�$6����9�<F	�
�R*j���L���eP��zv4~?�.<~��GB4�2>�rC�\n��]��7/fcqBG!s�>O�ZA�?��X��x��?����9�Z=��%o� xB����NhD1%�;�Qh�S��J0��g����T�{�o$�<��gk4�M�`ҕ���Ө��S�����#])T���+����������όD��K[<{�
��'�iaiV[`�:��7��P�3�Ja�4 �w����D�n��1�c,jP�qX��W�1�+$B$��
͍t7	'}�I�[Z1=���*���xs����n�03Y��oQ���s��
V��F����X@��NM��Ξ���e��
��a8�����)��⋯%h#���r���S���[�,Ue�Y����>�R=MVi��>.m�����C$��-7 ��]%��lݥ��J�?�d����d��,b.L}J Y��3�d$�}i�\ l4Z)��ce�[�{k6[�*�\�'�'+�S������
"Q��y�x��>UW�N�<,"��e�3��j)<O��7�3��Ej�S
�o��هhk��6ў$<5غ�}��&LT����@�#9e�4%��`�b��麐as?�fk�<��tC���t�蝿Θib���1�ڝ0����e�]j���$�&������r���������C ��7���m3R�P��B�:N��� �zr��[��}A�-�8)@p-�����u��}4�(��=%1���>� m���?
�1`���ȹ�`ϲ�}.�Ur{l,�ǰ���C�4��^	Ŧ�u�2�����p��O>
��w�nQ�X�qrK��<Xc���(�g']ъq�XcnL�7j��~x.^��w�{��|�.g�&�ExO��:ȎZ���d��hON���$h������7K��.��˵�[Ɛ�V��[w�k�H-��%��١�$�.�H���q���e�E��Z�x�ÄOm��ƲK#E�W���sU_Y�)�}?8_�â��4�����D��mZ�6�h[���1(t��u~7O1o�T(�j���f�u!�x�h����#e?� �¾=��/�^Ŵ��r�����|n.R\�p���̂I���7�cJ�dc|6�X���ID���W(k�z6��B�������W�q�X�cI�72����M��S#��Nn��VZ�t�ys� �I��B��V1�?�/O��Еa��We�^֒3`�M�Et�85�*n�12�^�r���@ X����x}�� �mQ�qAkqi�F�e߂Ŕi�-���v�\:���pP�cK�6��O��>dy]��cr��({e�c�Ĉ̷� +h�E\9���3��>d�4L�g�d'�m{�L�,��ʋC����Ix�W��F�����~�L��&�K��C��rJ�æˤ���h���j�Jh��D.�C}�ղ��r<�\��ޭܢ˜�x�oM��N��I����x�mmg����6�vt��h�LΒ�
Tb���2�Vd���� ���H�-a��R�x��q@��H#��Rݡա\T�p5�9߶�7�M�"�9����ݭRAC�[��_v0A��N��/����Ц�	�H��}��I�/(�����2c�T���&��0+�U��g�h5��7�H&p1�X���O��[?�U��q��.(dŔ�cn+��B��f��T>�h�PF;��PY����q�*&_Su�O+�ap&O�.𙤉Y	W�!�8��j���ƁՌ��r�%�8��� ��\!/+xwd�=K�S݆��Ck��j
�h��C��p��U^���n+�)e,�伤�l���dXZ���{�ι��B�[��|?��ePń>������S���:@��R���΍�^��H[�J��;�;����,��/1P2�͍.��@�V5Yþ�7
�2�9�D���S�0}F`ծ��_���1�%��U�"$C�_Uc�G����h��QjW��H�-�&��V[A�֡�j<��in��DiD���iv��7 ]ϛ3px3��N�?"ֹM<�T��3���<|� �CO�x�t�{n�ޘ�G��QI�pm��RfvAĸsy���[���n�}�V�8nP9�6���z�f�@b�������W?z�4���Ѵ���R�F{M��T����J��_�rd,�h#�G�vʆeư�-�^��ܺl�A��쏩��&�q�L\��k9%#69V�	�O[�OH�8ӎ/��am��0�Kr�������oH��Ʒ`���%�/�b��J�nZ�FN�Պj�˫г����	�/k�e�|�{������R45��u5�[��,p�D��?c6h�!�L}�D�8�,�h+r�)C��c\<��D�M5>ަ�R�ˣ�-שp�<�G���8�۽
������&�9�������oe˄�5<2>f�F�c�&F(�����"�N��ѣ�6�t/��=� d
i]]��v�͹M�~&s�qH��h�L�w�Uԋ�s��7݉OW����f�֛SjMا��}�w��u�z�����a�H-�Y�r �����=��)n����w�hv*c���da�}�����~�鄬���݄�̵�0���`�:{�G:�Y+4g���r��̧̀B̊(Y,�z���Ca���k��1�^=��wX��
v��i�A�-lӭ ������J���.��⡈ �f|x\?u,[�7��T��5�b��Ϧ���%�+�^���a�"]��ޒ�y�x#vw$�(o�2 '`����q`쩠��8.�!o����ꀩ�pj�2N�W��9�v�ppL��5
��\�+�U����Ⱦ1��Y�LU� *���In���UI��qBl⋔z�n3,�k������q�%mL�|P��	����;��@���Y�f�*�8�*�-|c�q�C��N+�N������+�O"�Y��U�5%�*0�!ʽBL�Ȥ+Z@{�'Eu��\���QG� ��P4���1:(�,>8̯��ɚ��5�c��JФ8g4����=��h}��Rgv�2�����˿��Y���o�%-��q��j�<����S`�-(
�X�埒��F�ϡ��~�-�*xF~�b��B�c�7:Z��Ytu$�''���G���J�<Fz����Q����,�3����1ZE�v'��2��@��Ө%n��F�uhx���6�):��Ǜ7�ܱY�+�[���������]_�bči�P�)������"��l��.!�M�W>�ʀ���g�`����?�L�W�n���qw�9��4��:��ճX$��VH�!���.R�2�a��W��։y�TŶ�E�p�HDú�����y�sM�&bzs$�`�G�"mw7n���x:���O��:/��Ɩ9�"
h���t�V�@��*g����T
�M3�s��l݃��J4�`����]ɭ.�V4"?ߎ|LE;0
B	��6�� �E.l���V�Px�JA��k}u5�L�0ܧ/�ǻd{.�L��2m�d�,m�c��b����=�vzv��።���gP�:m��	�
;�W�η��1W���Fh"���&�Jp^t?9�x-#�}^��z�j*M�6�̃�8������b+��.���bEe�_�0��%Ǆ�Q���aU���KkЊ�/&h���_�n����R�f�����(�F�J�}�i��*����@�����h<�=��Z慉���$$2]:܄�����2�ǭ��N�&�Ua��1���6obJM2{�J/AԂ3�9k �F��-�\l,H�v��d�z�.(X�u���I4x�~�T��mU;Łjf���Y��b_�w�Xf��*$^���jҲ z�����GF�;4�$^��U]iw=�����_T�N�V�F1y��L����X�`�	Y��\R��[�W�?�x��/3�ulR��Ƴ�uI���f�O[Ǡ�9�(l�)�����Of�M�F��J��q�d~�����iܽM*�0�SO��W��V������^}����R��E�7�TvD�v �l�]���r[G���4��r��[�^T�j�C��v��� ����=<_����/��J9�H�%�2Qߺt!�� �Y.��mQ�8�}�	�����P?�L^$���M�i"���O0��i���1���p�v��E!2�e����P�7�>~���f:*S�;��'R�;�vU�g�ͳU�{�7�@A�
"��b{�@�ə���C��w�CM��k�z�>�)��BL��nWC��rY6���d���L�b�s+0Ra�p!��lW���B�#!��^�о�NG���<-2���}[�Hm.~.��1u{�5�Ͳ��ܐ�?�=�=>P�~O��L�����)�%�$�0��=��������!��`��qa��<��6AľI��}�g�:�h}�D���Y���a͇]����|%��w�A����\���b�i��29��
�th�	Z#c�-����,�����c�JCBo�-�X/�2��3��^M��)��8[�PB�Oi۬�Aú���}��Q���y�1��xI�S	�6N(_��?�����C��7�r+�%3����?���q!�7��S�ѡ2k:J�꣬���n��v���Y��)�@Vt}��'�
�T�����sN�|	�/c4/W�:-,��wr)LP8��Y��������c���iě��b�"{��Ry{��S�#s��LC�$������kl�X�G�� ���w��%�S�Hz�kSh.�ae�g�¼ )�xF&��?MN����Q���R�;$/� ��S]iy�+
���7]�r��=����/7L�i�Z#Ǵ�iC��R�W��K��9}�"f0c�괧2)U�;ͦD��PT�g��匬)]ۯ�*��ł�h@��ç��fw��s��J{5�EAs���M��N�B����
}Ew����Ի�*�ť,ږ`��Y��AQ�w �`�9����SE�VN��eJ0�t�� ��&.NE$����?�R�Jۛ{��t�=��2�l�҄gU�t�2/'�sW-u��>c:3��Hd��� F�[�"����{�:}���D��~T��c,�`[X�%N� �2�#��j�:�˰S�e#�j 9�L��}=��s\��3qTU�c��7���K�����|[����.GJ��8�O��Ȝ5�
.),��%��gifz�`��Lj��5`y�:7�
�֍7��UX������e6w�Aəߦ��Ü��˪qР�t��܀"���ql�&��>���Z{�_yӿ1;��'9���,IL���s��Ӧ�~���Z�֕K����b/��Q�n�����F�j��5�ГI;�^d���X��F�Z~*=&���/FFU]��HB)7�jZ`3�0�q�ЯI#��aq��"���p��PeI���= ���� Y���b.o����1gM0U0	uOIW�@6>�����Al���a�U8J}�bYt�0�Pf�Tc�t�[�̓���y[IT��F�G&�76��c�rN#e�LP�Y��e5Cރ�;9��F
���Y�i�eQ,�I�1��.8,$�sŶ\�FQ;i��y��4�q��C�4;r��:�`�]���˵�Uv�W�c�������,f�=���C�\"��t��ϡc� �./4@�EU�M��̣>�_\�I~��>.��.�urO��ʇx��?W�SE�B5v�ɐߘ��^�D5��JE��S��-ꤞLr��zi_������f����-ٸö�5o^�`������C3�eعH���"ʄ�5�v��P��U�Q�#K���y��[%����H��#���Tm�M�zpIK`����e��_y�<���n�b�Y����m��$�f'uajo�#� ��_��?g�m��r,B4�|��"�	TQ�󯙿J^\2�Z�wZ�����+��i�"S�z,�O�L0"�����4���'g�E�4|jٚ�Z�85���������Bo��kc��7��6�P�J&G���m�h�~�Ӧ�MVn�������=��t��>�m���'�R�^J��>���� N^e�X>��/L��TQ�N�WN���F��P��:<�Ѧ\�)0���/���ܨk�舠�D?e�6Y衳�¦��bϱ_{-ܭ�saT�=|]M�<�+���FFF����7­_�"�iu�qK�JO����D�G}���ŗ�r�p���Z��?,"\Jr�p��Ľ#�Osw�V�x8Urۓ��
0kj��rIί^�5��2m�W�&�_t�P�)+�f$�vs��B֪��4�7�EC@�.������=Ն���i��P�	�-�)sWÄکvUD4=׭~��#?^M1�oA��}0Y���o4�0��̎��saF:d�&���[c���'Z=O�-�|�2����R�>�}1�/u<���_�3�n�:��S<�r�D�:Q0}
�l3� hTn	(��*u�a�������)\5ձ��n�4P֮�F�T�������Q
���P��Ǿc\�Iv٢�'i�Y 
����h嗵�V�_x�v@_�K��Q��E�FOH�/Y�
켻	���b=)��P�@�� �<qF�
�-[�v�����)�Ћ�����NG(�3^�WE���e�?�]�\�ن)A�!�g����f�1>1-���&B��1V.�Ԭ����s�[E֊N5��>D^���d�+Bf(�7`��0A�bV�n��n�h��`��':��2@������5-"�75ں����`��@����j*�~���������N?'���(��ܩ,q˩�8�#������I�Oݖ�c��p.����i%Ъ,Dn?L?��Sl �K�4]��g 1���e5kֽ�^�U�"1_��G����K?_2���_�ZX%i<Z��C3�HS�Nɰ���j�%��0e� ��ϖA�P̄,E	%���Pؘ��l�|쭆AX��`xWka�.G�����8���C�d�;�@�����ƭ��$Z�D��ñⱺR8����3�G2H��)<^^��N̙�8�Cm\��>�8�I��8&M�K[1&؊�fWi���?&P��g�Iu���Ayr@�9�EG̫3uu�+�2k�����\$�
�9��Ȩ�Y44㠈���`���ˬ��s�x�����xu�����H&Uמ� ?�qP��e�aY�=��ߞ�$8<��4���*�6���#��HS~�2�(�^�X2l�p&<��%׬x�:z3��sB�ʄ��L���ܽ#=>�Ƀ���uɼo^�L��� �4\&Bx�:=�)��U+��Y���8P�ыՒ���0�>�	�zmH�����p=�ãc��ƥ'�^��AZ+�k2o�Ò~�d��!�ٰ�,�(%4����M����G5��Ov� >u.��r��b꾺�6� N�-LGr�.	6F��&9�\KlO0��Ʌĳg@�>@E����`c�l^�J�� �e+����|��T�z�9�����Q���`�A�ph`pF�ԥr	3�Z6hSF�����t�	�nF��L��t!�k+ ��(���;�
���-;��r'lM<(��g4�GXՇ�e��δ�M�cuK�^Y��X��}�h�����ދ%���I,��^y�S�C�x�~d:��8��t@.l"����X�H�R��~N{Ω�������tMUJ�Am�nM}��Ʈz�GD]X?f�K�T�Ac@a��}yu����΄~�9�����$%<��5}:r��1b��i�j�����{#z8-W>e�u��=�fBZ����OU��E\��F�Pr(ƍD�Cˁ���zz�B��z��d��"�_���	���*�	c}�ZTГ�[ՙQ�$G~�;ש��*�YgA�ڧ�C��'\�HL���q}��<)���0��>�,�o�Ä�Y��H��~��ၡdޒ}z�S��!_�ze��gV��t���yH¨3`���d$���8��˄�x���Q�g,{��a�)�F�K]�w8Ąy�Rg��(=^+��\H��b��"4��������2\}ˮ�:1�4A��6�g���P��:�vT5nX��e.��I�l�rz�}Hh��YzYb��ܖ)�.�<��C����HMx�~��op!�?��hl쐩�I���������Q��(Y�}���؂�R_�<hIX;w:��@�6j�X���e�����i���T+��s>��3ƴZ��~YC�xG�32��� $.��L ������M']�H�f���� G� ��W�K׵aJ�3A�E�K��ghz���	*�l�DY7=��|��$�u[�4�w7�O�R*��u�PW;dV�t�$�x��-5Y0�l0�Q(&�|��gdh6�� �"����ǹ/�5�Huq�a��ps�kF u;<<�v��ދ4��;"���oD���|S��K��60��ۦb���2NX&.ɗ�`��=�:ÿ����%�#��(���{��rZ��.jΑn��53'������(\m����Z j�ν�
-���j�K�X�1 i�_.��Y9��G)�E�

�i�N�2�����~����*�n��y��.�zǊh��*@�� $�E��w����]�u�e������;��<���������ws=;.�r�Q�� �0]۝ #�o�!=�d�9C0U�ahGxn��@�1rqȻ�t%@��CB8]����^����P�l��
�ח9^�.`��`�<:㽚uvw�\����|�n ǿ!	��w~�aH��^e�s�Pn?�w ��b|��m�g�=���j����9�Y/����X|��:2�Q���	������"��ˡv���Aʆ�
��b�;r���:�h��Pc�H����G�b���\��Ѧ3g�Z����F�M��#-�Ï��s)�-�%
��h��A�[�{���a�c�/�-5<�=�>m�Lk�*�}V�Z�#߅�� �'ϲ��E:�.w*�Y������;����PgQ�у���=1=� $~YR#?U�J7� �uC�\!�X���l5����̓���b|��_�a���LH�O�8KZ/�k��� �£�@�ih	���?J�_�_��!�_�#T���⮰��n�y�
��%�Vw�������%d�уaB[6B��`��#���ʎ��<��(��*��H��h��������������%o�n0J�����W�� ֶ��)=��/��{"0s����`�u�e��q�fq>,)�.��=2��Yr"Oe�'<
k��-r��Ѐ5��1I�j2h@
ӵ�#�f�[ow̚%o����w��TӉ��D$O_�u��hTR����Y��Y���0I�J	�݉?�B���8�wը��Qԩi���-�rD޹1ś7�{N�kY������iqG�?31ki�,�|:,�]�3I?;b�a�%l��҈נr|��&�C/$�W�UP��C�-�xT�K,�Rļ��G?5&[˦�l���'	/H�8	� 7�jVg����|�aAf����N�D�ZYH�D�5YS
�i�$
��e�qV��ZH��e�f֠(��t�>A"�TWP�^�������~B8�5�x �U�9��g���uf�Z�2��ښ��yQ���#��N�%%�(�J!��'�s�Y�?�T����8�7y>K?wc�!�U�40�����$���1��#7��;��r���d�Nu���>(T��J5������Ļ���.0!h\6p��^q�8AqG�J����QY?�8������CLP��ѡ&��F߭;���t���z��$7��;��F���*F;�7z��{�өO;�^M�A��
�Nsu�<�4\���(�͏z�B��[��mv�FB�MD�8\TI0n17Ցv���lli��V�:�8���́%	ϥ������`��B���~�p�0>yD�b���:���6��W#�­��Q�o�ʆ��䵯ҕk��%�����x�y���чB����U���k�%�6�sɺhO����pZ�wB�y`f����7��*�Q`�ӯ0l��D�עW�N�UJq<�io�ف��{ht�����H��c�ޘp��ve�ܼᵎ.ZX�'a@�e#>���-�F��3%�Uv���d��R-t�	�� �E�!.�*|�%(
rl�����^��ZC��u&��`�8�r�aGƬ���q���v,����*�O	m�y�V�ɶ�9�W�"���<��/����g�"i^�u4��{z8y��H�m4��4b��'92�7�<c]�\1���v������#��7hFo��F�@��aL��j����m ,X6x�/����FX�9�=�tQ�J�/	���,	C���TL�k�{�q.̱��O2�3洜j�,s]���[���Pq>>��~1Q^��J����-K
��ad�OPq���j+�m�^

p���2�c���|Gz���MAR���d���2��{���L��D1c�ٯRX�d'{UoƠ�	}�������%¥�ǭ$iIb뗋�"��$�G�g�.��K����ڟ ~�j�d��9�J}�y�Ba*H�I�E�mu}�	!׽��<$���S�>]��b��S ��ߌ+�,|	Љ�M#cb
x��Cp��s$�*n��|��^���w�Z�!n�犽��T���
E=.��������* �[�̋��\�e���yTm�W�D݌|c���Ѝ���b��:��
4*Ͻ���xY�1�EG��:cU����KY����*�S��!�\��O�|�-�7�z�~L�sT�e�"0��p03\%h�D!�i���`f߳}?X9R��b}�����BVOYq:�9����p�b<�6�J����3L�U "���1n���fU�f&K�� ���&��h]�����3Ǘ��(Jor��5�Cz�a4GU���!z����p�w�B;�����Ǉ�wtD��������d����<�31��R�6q���j �Èj+��T�.���"S����ߦ����7��H�?~ %�-�֊>�m�7���V���L�Q~�V����Ge!�1�\W� ���"�%�C'����{(4K:�ζ�$ !��Z�>ۏ�/�Pb�v:C�KI �f3��������������7��#�r27�<�-�	�!��VSn3�
���?�<�@��,f�?̊�����'g+׿s긋�ME8����8P�ɖ�=��V<pfF.�)��?�zh %���;�[��[�:�Oa!v�mi Q� \���s�[_���b����p:`�[}������ox|sv�����Ro���=�j2bm����$8~
�>��R���*j]kJm������2�5zn�u��1���6ކ��AXd������M]�5�����z�YD�q��	���ot���K�u��&�I�/�g�*���_	�b��4Va�3�T����AKx����G�G��P|\,X�`�1���+��]s%�)��,It�rE�7C�
����+����Ǵ�=�%~�z7��{�vu���|h�8��/6�h-���V�?֦q��u ��x��.xǳ
�o��4��s-ԽWY���ҵ(�Ӻ3݉��	x+�Ǟ�PCYq�/c
�ƃ�Ꞓ �C���O���-�r�ο��k��SE�`������)�X+�eb��t��t����)�$��_�2&A�/[����5�Шm����_�Gq��h~O�V�^�~���3���z�Ҳ�SP���-W�5=�y~��\�7�EۋZ�}|��U��y\�@tL�9������%��% �����׭�������W����4y�~ͷ�{��������~�i@�g��MBY��H/Ӭ'��xc���7������a�J��ht�s|�B�������&T�.�SI(���![�<;��0'���\O���
5?�/n2��,��8��b������`��T�Y��c��[�#����35�W��O��rȹ�ɳ�=��2�����2��A�F�E���mT��<��y��g���-]���x�ù�.E:�	z���g5<� 0#�yQP$~����ƨ�U��U����D�� k�����?ů��:�����׽���U�$�����H�jҞ�1ؿ�EA�>=�q�˨���?Qo����;���>F�m�QY-r�yD?u�1�/��B���̏��Y�[4x0�v���I� ��@Fp�y@ԓ�Qs����W�eP���p?q�6�J}�X9�o�M�H�T�`T,��[���b(U/�LyB����i�@��ei��2�ɸ�S�d{�+|v~#;N��K�����Y�pP�;U�d��E9�[VW��z[�
q"��nh���!��M�;��`����Z�N)�O�Р���Uґ�f$R�(Q@z����_En�R?�P���4uwKKA�8x[J�
A'��T���Y~S��sG�X�?��_�m��p�1�=�[�E���	?M�[9��c{��g|����y���ipl.��@�>FG���������N�%w�l�>���	6�����Ȫ�Bk�����fpT}��i5n�.�P�xmI��E���H�_����^��t�mH�{�|���f��߉_��	�+���xĢ��`���[FF�-t֢D=�IK@ 5�f�z�3����:�~�뛙�P�DEI���"�<H��d�p�s$�*�^��_ߐ����hy9��F"[���V�Je~���%��2n�����@�e޹f���.��s��xh�P��Q1�S��2#�c:o�u�M(G/-�Fx�p�+����a�`h3�D_KȄ�b�1��y����e�x.�]`OU�:�t���T���&��W�EZ֮s��!�&田 ڣe{{�O��(��;S�R^*����oM���ǈ�v$Vl˥?o^��v���;�+ sS_����M�S6j�K��=hO�&�E~�νU�z��>�|�Ϲ����L��iƷ���6��3�->�3r����F�W�2ͩgUY�[�}zBsV�NU(�N�I�K�()��O�|����q�齃����,f�K����`�B^���2$��yn�	 ,����c;+�m��4�]H�||�v�ѧ�=�$�9���gn��92��JN(���r�Dq�3�
�#%B8�t]1؄��_�RUb�GOSV�b4�q*f�}�re��+��گO��?�t��4'�LN���n��Y��Hļ���(������ƿ����vh|�u�n��9����fO���1bݎl�,�qKwe2[ѽ��#r���m?��/ءJ��j�S�=䞷 O�3�ۘ�{�:�D�������h�4�5��8n;��;W��T��̤>���~#��#���4��4=V��3��	��`اi��n�	z�6�M��-�����R�a*p"�\��'Q��?���	�>�.h���=F�������]b�1W:�S[��=��|�����FtɟU}>�i�P.�tl\vĒ/T|�tDN湬������ҝ<����΄W�-[�Ă�E�?�E-�X^��rȯp5r�y/����{����aP��U���[Q��uC��mK
޽�	�G%����ᗖ�"��S����4��m2�gw�A��E�5�_���Z%���6�~FB�{ro�++ҟ]��bwQbx��/#���#��ǉ�bY�͙m�T�~�>�//��l����c���<�g�: ��ʆ&�3g�GE}�����A�6��Ѩ�K��б��~�fBH�&H�2-{G��J��Oj� x� �m�j�FԠ2m,� #���O�q�$��d�X�ȹ�[3SV1P�5�)��yt@L�=#����w4�����T��#�=�+�=6��4RytJ�IIW��*�c���̬�)Q�/�����x?��{E8u��re����k�I���1���>*+V�"Q\�Lol_pui��c����5�
'ْ�}j͢����I�囱�qnr�۷A���_}��9.8>�dq�5C�����Q�-��?�-.�F�e��n�@F�}��:�G�Թ����`� g]��*�X�bf%��vb\��d��*�r��j��v͟��)Y !z:=������r�c�VFx"�� ��p�\���Nl}��j��Q��,dU�������z������gAŧ`�`I[@�h
�{S�%���x����p��W=��<?N1Ha���h�O~�-	$��|V�N����)U���ƍ�ˋ �Y]B�xb�q�p��v��� BC��!�0�a��l�ڷ�k��ws���ƆLC��L�ᷥώ��N�n��c�(�<�x5����k�Z�� &!+�p8zPB�����ܖ*N�-�-Y�v�$Bug�qE���J,]��w_�uX����I`"����	2>~m��0X��j0�4��LM%�˯�ZI�@#u�G��KyL%q�ճPǲ��B;�b���r<�] W.�B�k��B���<)lta�>u/2'6%0;�O��#m�@��-ވ�.p$w�5+0L�j���k��o�%�4�	�G���54vĩ���\�yP~$�؊Z��Q�dM����/�$�&Y����N��)1���R�9�ٰ���7�:��`�1c��~�:��+�D��P��~}@�;(�N�EM�G��wd��A���~4P��g�n��5S_@�f�!+_A�W�ͣ�y.�{�ad��_����MZ@5�F�k���w�����q4�x��7��V�q�U� �{�C۟��yYd�į(�$^b�CK��6��zd�L�sy��F v����M�n�>��Y�|���%]��x�+���v���2��a����`�F��3���܉���ˋ1Zx�Rڝ*9��a������5��.�(��v���'<�P��P�.���/�q��n�|&l~�śf���g�_H��t��!�^�p��..�N�r��l2Ҹ�`��o�h��1�J���":V2yQ���vdV�&�+�:)��hE�֐���E��)�~u�
���c ����q�,�*�DbI�Q�%?��w?l� ���g[C�+� 8Z�W�q;@nR��nH�V�Uq�qsC.S����JBm���"c�����a*��ZUf�����/���n%{�t5�~W��KD�G��@�^�P�zf�ܖj����� ���뻡�� ���	_���+�r8e�B���M�3�ه��H,�)�ħc�@�@y]�x&3�""��xe�^�6�	�s��<�����*}:%�_Ge[�����q��ʅ��`%�C{E� ���J��h��Op'Oy��o@�W�Q#�j�4�4}�{�'���̲!�P��_�l�@����E��+w�	�����ok
��n�XzuM�X;3���g����޾����>�k�c�B��4�/UQ��r�4�����Z���c�#�8�Co	_4���3��Kݿ#���L]�=6h!"�n���Q��� ^���s�T ԰�RS{'j_��k�G�Ń��)�
)c���n+�$�&��>�	��`��Es{���!@��8�qMl�*�����$��Z��4~��@�8D*w��=4�k���WW�
��B+=��?U8M�9�,[8��c���J�TB$��Gj��Tq����#�b���T�'~�+&��I�kDX��@ȁ�03��R�/Tcɻ�p�sQ
r2����3�t��6��ͪY9�������w���\�<^���5B�n�J�Rrj�_���h�k�����M��w��_��%���L�K�R���M�P�����z��;*��h�����N$�
�¾����o�&�{4�] c�E��^���b�֒ ͑��Ұ$m���:j�\^	4����(0_���~^U��SY7 P�He�,��hln��Q���h1�.ޝ4�u���@lݳ���S����H���;pȞ� ��2)��G���=俥:���p�Y����6Hz����=k�ͅ�����y�K�H����1�؆%�@n����g�_.�PT��p��#�.7��l?���Z��tB�<"M�I���{zIǇr�sJ��/!Y���b%a��$-'
��plP�e#��<��]�'�¾)ױ��d�\f�gb	�� ���U�[�ߙG���#�M��"F� Tn��┲k�K���:����lTKt0�$���*	j�gȷӮ�)����\��;�{̔|�N
		�4iR�}�����3˚J�OO�Ѻ�߿����0(�\1f	�i�ւ\���O���Ȓ�qWfA<J�I9kǍ�ꏖ�qZ磁��>@�������%Z��w�Ηq�����-��x�2I'�j�Xjse��z��76�<���9F�@Ғ�/~����/��q�W����t��c����&=[0��������C���}�;�.�FǱ���P��~���t��$����v��#奈�-�Խ(A�W��;8�r�<�f������\��O���owL`��ʮ�>X�Ζ�A����Ԍ4)��G��NAiŽ+0����������n@��/LLM�i0�o�%��fP��϶�ׂFr6��t�,�������¯=�6�������v�e�oc�*��Y�Z��^�;�l�c7~צ 2��
�rr7o������r��h��8GJ�T��M��{)�N��'�iq�ū���9�Q:��糤M_1Y$�i����H�A�V��%��,���J�N����D�����*��}Fk���I�,��#� s`�N�;\J��
$ѼF�`��	/2B"8��&�3^�jc�Y8�v
�^\�n���+����C*���t���d�n1���Eբ�v,҄���k����T���p����Ȕ����E����H�d� ���+P��>p�R*4�>�q��p��*a����C�?7^�a�?�
��bX{��%*C�m���7�>&1�!s��ӲU��8���VCn���w@���5�G�o�`>-������Ҧ��!V�����j��`v�OL���
>���� �Ln��Xt#�9�W�t�[7f�#f-�/�tl{���KC�I�Pٔ�!m��%x/�3�O1:Y��@���?u��|�b.�斘�XLl���	)� ���RF��#V�ZQs��sD�{��<��'1���:=���58���I.�a��}�o��.:8#	\�a��{x<M\.A�@�TtWP����T,�#]L{Tɺu�i>X�2�ɍ72��Y��g�mh�U���UiM�Pu����#O�C��s;�������.�x��׭����b|�1���Ѧ牗�d��a��3@��{ X�uö+9�+7�֨oD$yiL!��|ʕ?�W,g���6������'��o�3cg"�	���f��~ �����m�����0��V/������Eۛ�5�����j�I'�I*����i+�W�=p��D>���ËR2m���ա����;ډ��jhp��~�B�w ��yp�TJ��'H�$P/�O��zQHB����<L�_ز{?�7[t����$�̆F7�\��:�fO�0+lw{X��R��
�����%F�V�ɟ�ܜ�1��>3;� ���~�d9�ۤ��J�I4�Qٯ�B�1d����Z]�4:��5әـb]�tapPN=�����RŴo^ �XF��㮄����e%J?@+�+@�t���^��X�D�-����&=2�*���vϒ׆�_Kd���,�- ���ςU���C���RI��
v��Y�qy��ʋ�X��z�=��e)����w����1]���d���(�<CXm&�_��#�εQ2a��8C��[����
��:�:��O��?Ę���w�&vz��ʏ���4�^F���aM��V-��i3���Vx ���M5*+����c�O�Ȭfl�2��qvYX�WŒT#��j.e�LBӒ��4�c�K0�j�l,76�ͱņ[c�yB">L4�2��nh�٭��Ҩ�F��\��f}�h=�B3%e��B�Tb���x SZ�������s2㘝uGk��⷏x'����6֌}m�����5K9�~eI�Q a��-`De���h�>�Qcp3�;���Pݙ��Q��Q8ͬ�+�4ud)�_ݤB����.g��_��=Ķ �����sS�`*�X���{�--{KHg-����4.�1�TS"�q�g��p�=�VR�H[_��C*�eÅc�ɩK�z�Z����g��/��Ͱ�A�u�u��-�I$��lG?�c�](BV�+ �I��ڥI�����������PQ�7�����a��5�KA<tT���-�"��
�y*���+E��},�&0{3��JDS= �q�0�]�j�|i�	}p���:��)�|��#o�e���%h3�N)C9���0��H?��2�����\�ǳ��"�&�+���'j��zj��մ���U�q��x�'BS�_�����u⽭����� +����C���ʾ m ����fƲ�1��懁�˦�E���3qݨ�+��Dk�Xv�CF~�_4^ �?Jm������ԙ�b�
�o�]5��H���&�c.q��hc3�P2ˍ!wWD�}𻱻�8d�kqH�����oM}_�,�����.�]��:�m� 19��^t+�E|����<nq�T�Q��V����S����� �����p�F�~"�QP+�
q�)����X�b�U���G�`�%�j��)`��R�U�
�����C���p�0�-�9\P���l����b��Z��qY7|^R!�Uǁ�W�78E1B{(�}�3?d�6�m~bʇ��1��PW����1�:3L��̸=Nd�sT��X΍�.����,Q�#�V��U#�s��	*��	k�T����)w��<����|�(N��7xo�^�:�t���M�)�e��{$0��x�Fdɑ8�Q���<KŲ�����G�pCo��)��$�Lϱ����fݏ��S27�8n��3�^H��aU��͘Vf�^���B�4O��\��:�("�%�|J��z��x�,$��t��]A\���Ř�O�v�����_�e_��[$)o����z瘧ȜUŃ����{���;�dNh�r^fiP/!&$?n�|nA�1��J����6z����A&{:�	:R��_�����,#�8I�B6ΪdH�x�S�e��+\���o175�!����a��n��?�:��tO�2η�Ř���a�AEn�?��3@������x���.�nxD�4�zz��^Y����Er$8n2G��8B"�F����z)1�M=a����W��5�LMl��n�	i�9��ڶ95�DFQ��ĂFʅ��������9Ү��5�U�H;�,�fđ�aA*y~��~��|���!�2���X�O"��m`�9�oK�)@<,��Xl��	؀�o���A<���oa0hfv�2�m�+"k�u5�ص�P<28l���?����Ч����^[�,��~;��1���/����(	v|M���tQ&�\%#qf�2q6��f����2G ��&�����S�G�3�t]�m���<����_z]]��k�h)���]�xc�q��o���3%o��!��TS��gf�.e����0�*wrM
�9�R�0�I���6
yZ�fȺ�QЏ�����I�&��B�3�v4t�	����s�h��8\[I;� �bsĠôRu�|D���Bl������=qGc�iW����Yrx��stڂ�� {M��\@K3�7I�I�N'�_~.$]�!���%��H1��?,�}����bq�G�8j�b�ùwv���pfd�N�/`��-���^�ﮅ�`�r"���e���_"]3��B%\	p�̘|^���B�
�u� F�D@�V5�+_�ژ��&&
�2Z��gg�yR�ߡΏC��eh�|����F����y'�T}g��©�\@'����j���s�*�� i	g��|��EG�ͪ�N�ݱ[���>M|���K���,�f�P��e�Y�'�;P��t�8x�e(;�J��>i`t�\��k�iR��Kc��-��Z r���9{��u��������cp���HYZ�pJ�i���=k�W���ʤJz"}؟ Z�$S���ޛҮw�~��h��PWƪ�*�l�Sy�6���*���ꥪ��� ���u��m]�n��A�W�p�E^ck���vi/[B��C�f|�����a�!1/�������!	1m�ߢ���wʫ4�aFN�Ye� �aH��9�Y��C�%r6����;����ua]X�w�	=�H۫<]��x��Bj��l*�kLco�gN���Pb����=��]�7�n�5���+��o�i��B�y,?�lWh�f�kM�(�c�sF:p����4���eV}T=�k<Qb��oK���l�D%VpY3�1�~֝�p�Y3CE�F��dk���UJ2�Rd6=��m۝�b��X��-cA����ni0�7Eݒ܌<f7��I�6����������ʷ�����]7��K�g�%�����-� �Cj�
�U�Sc��Y��cYU-�%C�K�^�uh���^O�Ƙ^-��x�ǳ=*�as{�� ��X�o`��؇������{J�B*��5�^����Y huo@�!@_BKeF�5����~U�C׍J���#�	�3X�w+���C���>-Xk'�$-�*����؍wTu�M����+WR�u����(3[حm"J�)!���l��;��U�y�v�#�<v+�3x���36�
-'ߵ���n�}7p��&0}B0��>���3*5ש���`����w����ƞe��$g�[*ڲ~=@�]?�x��u��p�#t�n�B���ng�+
8|���yi�SI+�3n�\��w6M��Owt�"��{�|
��A��wӣL٥\}���5Q���GS&%�H��-��ᮗߎ*-�dl�be�G1�GQJ(D.33�:>��`�������	@�wq�NR��7m�����U�#�Q/���Ϥ��!$u�Eݿ��wе�5q��b���"2�8�ۼw�w��YoC&����B���ڊ�i��A����H���^|�!�$��N J��FN��?���V��^�1.�ɶƪA·? ��Se�V�<�����?ܥa��}	\�ng{eJ gF16OJ\Fl��dr ���)OK�u���T���ALTK��=��W܁=��ڧz ���x�X��X��'�/*X�Ccb	A*�2��V,���y�3���&�*1<�3?�Rg�뾊��X��zw2f�=�x����`5M,�!25����ŞŽ�?X�d礓��'Y�[�
/���2d���􁭮��y�_�����fD�l�2s��C/�E���wu��I/�z�	��IІ��:��ڀ0YTM�yպ�Aa�j��V3�i�����:�Q6��I��'P��/w�ଅ+��Ir�?g):�f��D�iK�EQ?�����!�o�l���+t�S��A�@�%}_]2����J_������q)���FҎ)�6�� �?��A�����hz�����Ɂ�=`�8�.��BF���z��?4��G��~ s��m��vtB��d|0]s'��M_�;X�yg��N0{�W��̋�p�FӅ5�����h���.����T��B;yI�}�jΉI�2,I��#)kӯ��o���fޯq0��PRn�-�~��L(��N�.��fr���W=�co��HM�';~{�(�y#��V����X�4���:u�%��]Y&ݙ!e�X�� E/(����N(E{�Kތ�0��ү�����s>��0(m�=y�MGc��n~xk.'��6�Ǫ�I��^�Y!Oí�m%(�)�V��ϵ&��#w(yd�o<��;���b�����EN5�E-���h+g_h����Sm߀_j�}�G��p�kC9Oj�،�B��m��Z߬����t���'4��)}.�7w���[�)�HP-ۖ-���rE��e����!��C���>���a��IVK�溺zuCY�A�	b���_kys��ˬ�1�7��w�򃅧-
۬$K�&%aV �*�J��]���,EL�yQt��lPB��B�} ����P �/*���~�����d���B��s�Udz��(��̽��J����"������C��*�"C&&��ړ7 X*�������\m�__���?g�E'{�����=��z@�i��vb�{����'�4GQ�1�a�зE6���W6PJE�fDu;��'߹�]��Ʉ�5?n�4!-��������]�).�%t{1��"i���C�)��G,�U��-����j��5&���xA��p:9{�ݴ�:�~���upZ�h�\�U�_�=y��6����.8e/�^� �
O�ʪ�U�3�؈�S<���j�>���hK��C���Ė��u�C�xGjA���욉gxh�wb^4�R3�c�!td��=ւ@`�ì�D2���&��A�)��%H1������՝��zXTf��1��������rV�/���~u���$�W�o���8��i��ܕ��}����U�����"��j7W����O�p/�{G���M���e�j�i�+>V�6G�!�E�V�ْF�VB¤��H����	���!��}��a[Q�X�	�iD8<��_���'a�I�Lf�V8l�'<�^�)ܛ9S_Y��Bْ��p�'��L>@kD�ϒ�yj'�g�l6��xm��aΡ��W�h.u�#�xA����~p�5&ٚܨ���
[N����8|t<T�Q}Bs@�a/�%�f6"b���Pg���+��E[t���Tgd�Mr[dMn�u3�B���14�kZ��>�TR��*R��BF�����|l�m�"c�(;�����g.P��w%ԩ��4��Q���K�3&��\����7z`uT�Lÿ���v՛{� �l�� �1	c+�Œo]Y�i�
˶����;����kN/�G�A3mb��.�j��ա�/��R�qȶT^6r����|�a00����v���I��ֲ7�q	�w*B��7.��y�Z��H)N?�J�1+��q`z	�h7�r3�tlL���Kxh �꯷C��T�ñ��Z�O����D�ފ#i��奖��V#��]��3"���<�" ���d�>䠇l�3��د��(X�V��@�CoeTѨ���)��0���E�c��[��_/�t�	�����Q�����Xi�r��/#�IIa�Ǣ4E#�A9��׃I��#찉M�����t�2T5�̞ѝ�k�2��O%�@�K�}Zkl�j�ˬ���^b���u�c@�!���p�Z߂(��³qď�q�򚹂��m� ~�Z�OƉ*�����LD�z�b�'��e��3��.�	{����KMV��H�U,r*��EU���uw����eV����O�Ї��/4�G�}E����b��n�xb�mG��[�ͻg����EuM��l�]
7BWe��+��rK'�9�@�g���C☸ͽh���T���l}S���6u-�.��Z��9��SvXc�
2<jx�.�ć�k�SF�oaėa��Q=<��3�8�Z9( �k�Qt�37�y=��Kl;��t�-�r��x ��Ȳp<�}y�\{lq�dm�����l�ù��	C��$�a�hG�6$9b��;z�F6�|�**dR։HLH�Z�$��:�U�(��_/fh]<9�����H�w7R��TR�@���U�0�;�OB�c�O����C�7�%�(�v�i��wl�q:w���ުM\w�����OU͟rbx�&:�9`�{ٟ횖��2y�+�Jzi���d�?���C��#Q�䐳���?廎���l�����-�YZ���nMkf���+�:��;B6�A�ig���, 3���&��;X��M��.�����ݒ,�x��1��V�U$W��<f�1�d��y�-����N�%�m�d�L�{BS�HY�g�kR�
��2_2�衍黶�©0�UI�x>��,���^�9,�O*IN��qZy�묕�Qӫ��&_�:i�Z\��HU��h�DW���#�~��A2i�@U�1�=����t��
1բq��Si#��!eT;��pW%D%�ͧY('���bL}ȗb'k��Z����W�VQܷl��\0e��K�N���p�8�,.H�Vq�m���	b������/��������V,�F.�Z���ؠ���;��n�>�-EhE0�g�� ��g#Y"�������s͊�`.�
���t��s��E�?��1w�:ȝ��*�N|)���/�<aw��+�\���0�(?�
sω��F�٥��ep��urV���G��eq`m�ă���~�.b�l{FȹE!I���4���I��=-�,k��n�A��j$l9��v�m�F&�G��e�x	Ɯ�,��`�g��hk)���]G�(Y���AC<�uW�9��E�k������z۬��OX�Y)`��i�/�;����f�:����ˉ���2������R����z����!��F���f&G����8@&�)�?�����n��XJ�S��]A��'A,#�Y$mC���q(�bN��<�G�J	��CF� ��
�9�����K֓�[�+a�n�HRA������m޵I�ֿ��c���]�7�������]����9(Yczɑ$��mʘ;2��s��/$t�H|�ܩ���{�\?E�.�jB����C�tk>1
��`�	��.nE ��D��Ɔ�s����^�'z�o	u8ƅ�VD�|�$��/��*�?�^~�8�q�nXC����t�H�U ���8���Ms�Tpڝ������E'��8tѮ����9bHֶ�~���x�����n�� �+�/H5_���&�ď�.�:�r���H�<�J2�8	����^׷���a�ȡm>��!�ܩ�Ln����������Dߺ�V�g�<�W��.��sc��o��5$P�SMf5AA���M��0Ń��O�M���|�{�s�E�]܃��C.s��>�8bA �[,$i �;��:,��k��d*ϰT�1B?�'�t!f\�r�:���sT�[�DpiͲ�f���A�Nʯ�"~���;_�в �7M�u�Q�eUFR?d�X?oZp�a���ϐ���Z�PgM�(rvǨ��_Hm����*�c�ӝ�?'?ZD<&�	D�7���:�������8ol��-i�MY�3�:SL� ������\#.U��t�ٳ���Q�ר�s��4TK��~F�����b(���E
�������>L�\�<�ƹ�x��J�mҒm�r�-1��2���`��K�(v�IOMT1��+��`)�{6�ΓU� �2艖9�*���3f�0��"кK��#8���iGA�� ��>UF*m� ����A�������JD,Ο;L���U�m��[s[,�߱z��	��'R<*v������ШR4M��'_�<
�G�0�.�� ��<PJQ`��Xx��- QB_[�Q���v�o�a|���_	Q�1t�����dC�$[Mj��ߖ���Z��?�;�hnF��`�^x���nXd�d � ,����fO�.�J�f��>�a8{��O�s�Ѩ{�˖ +TJ��'Jz��#s����%߱xY��߫�~~����-()>�6��O"�s'�,p~�\��E��GI&Bl=����?�i���4�騉��^>d߽��O{Lx>�W:���$-7�� sH��]O����59ǩ�)�bl�k�#�j�$�L�.�-7�n��`�֝��S��p�p�22�:j��zS�;�,�����ڋcd��)�J�`�Z�7��\'ٕt�Ʈ��N^b��e�L]��I� Su!�u��&g��.�R��� ��k�UД|�X����3��e�\y5�7'ZI�AϳN'�U8�j��xm��Fw��1)c,m�B�Y�?�>�g�u(�B����Z�|�!d�~�4�	�I`�# �@�.پ�;x)�GLm
� ���[���z��E��w��Z^�1J7z=7N^�82Nc!7�C;D�sT���0�N���ŕL��l.^$�Y2?��g��KK�M�e��:�۟���!s1��&J��s�P�[��:�ŠpX�D�k-�9��!h�b�/���{&f�W�W�U#�q�ӿH����A�L�+%C-2Ƕ�1��2��I�<]6
�a�{i^_ث�@�S%!h=�� �w��(D����
�E@�NT?9I-|����W(���v�x�������G��^��%�C�m_��>������x=��aa��EBH�%��s2���b`��k5���;e�ј�IݎfK�S�y�d��9	<����s$��M,Ձ2)�_Z���o��`c��"�\�_v������O��h��[Klz��K_��R���7�#r����d��m7��0%��̫0����HW�ZD�����Oj�!�i�Q�m�Oْ
m(�m�-��օ0]�n�k'I+�J��v��'���}#����ذK�`��f`��J?�L;�SG_35�<���iiv�P#N7��Q�KkB0�{�o���W�7.K�V �knG�ֳ�8J��	eᅊ���K�x��R7����3�=6�9������ַc��(����Ȓ;@�����Hr4{���"p|��=^��wN���F�m�nT�'�l)Qrr�ܩ�$/��-��z�NɒK�~�%Wt�ɮ-���x�8�ۗ��0!��orD��K-�7Ƅ\�����K�ԛ�ύW��v�h�1;��PXl���x=���_4�\���"d�Z]���9ZbFQ�h�H���:.Fz.�,Y�\��mГSs��E#p��#�F�%2��}��gy���"�:l�4�-���OA��O]F���m��ha��?��E��ӊgNV|R�i�!����&MYխ������Ԉ)����`'ʅ�zlR��"nK���w"g{�\���Ò��9B��kt��ܸ����-7�?7���f�'Ɨ/�H��zK�Bgx1A��Q�Bq����b���x�ӈDhm��ė[UL�������Ϡ�/�I$��κ>M`�2(*�.�J�o��b#�&����]�˩2/1NZTcM�y��!��O���,q~�z��b�n�����!�j���96��ሤ�}��a�&�g�:���[�A�܀A y P���ji�Z�t��)�޺�>����
���T�<(�E/���8��qDޥt����{o�SA�K�)�W5$��r�k
�k���X��ъF*��0.5�,��m�Ǡ��Pʴu��e,r�QH�G7]�u#�}�Z �V��|j����E�e�Q���F�L��c��/Έ�1�
n¯=�����yѿ5[g���v���!�i�`���F\mN�;�(M�V�ω���3�\��h(rS�{���� �����fL<��!=��9�Pֿ�r���L��Q�<�H�
4Mg�+ٶUF�	�6d:~����)���o7G�c7�����uG2A���D#y
(w�&��ep�DKX�'�� ��5 �hD���?;�p��D���~jk3��� F����-���\�ûR��Y�[������������q?�(�(B�����fnQY&�"�\�2�<!6�mw�S��xJ�tS�[��N�q@�s,�/�gk��SB�v<�f�vT�a^�_D~w��h`o�BnL8C�㤕���"�,�D1Yر$9Py�������X�*i�Qb�i�]¼10���vN�F�c9�9	��D�?$���.*X��[�I��@���Y�����Ɗ+lL���5��g�1t��K�{��qg�?���~YF	~��^g��?w)���o��Âۘ(	��`x-#~�f�C��BR��!ۇ�Q�Z�p�s��J�o>z4ڹh�w����i�+p0�����2���P��r��]���,��%2>_��sWE���1	�t�ȝ�����/P�GCk���B���$l�2ݹ�T���Vn� ���b�z�0:��������l��F��N罍�7`{	�ʲ�ka���8�N_�"��v��=� ���xca�k�^Ҷ�9M�*u��\�v���d�L
���H>���cy-�'� �sJ%��IB���2�\�)�eO9�7�ٟ4���1�-�I�n�#̣W(qXC[O%��T'LOy9��&��7��i4��?���r:"��*� �hZ$����f�%2Q;�"5�L
����cJ�>BU:�t���]���p\2�M_f��-���ɽ��y�����ᩜ��\'} ��EWH���筮�a\�H�W�: s�����ꦵ��� ��|��B���(��S�^=��$��$��Ҁ�,�/̌Y������w�䇔˓~� ��U�:"���n>ZuP�������v�C�J�Y.^o�	���o�M��������R(�_;Eٻ���	,�9���!�V4�6=�g��^-�҆�f�ɭdK�#��i���#�؞��o8�BgNe�VC�Ai9Im%r�G�:W|�J������,��9��H��DZ�	ܓ5�U����	���?g�W��"�}�#��=}@���jp!�߀�3�$Jj�δ
�"[�.�|�&�G����Me`�J��hH�%dȍg��=����lBo����� �Y�����$ko_ۛB���7*�[3Q<��V��v���#	<�|~�"�[&|�t��`�n9$ڎS-g��UE'���˯+i9�ŕ|�D��M��ۅ���tҦ�¡mM/�#�I��;6.�?@�����T���%���5%�n%�΢���OI�ш����<����;��P1ȶ�?85BE1!�-���}[�r�I�¬��O���!�e�%�s��K��'�hb�)0h"Y|:"=@�/��7@��9��T�Zt�:��Eɡ~�`~~�b��}�#}�3�<{��ܠuwĵM�=�s��5�@3���b����5X��߯<!�g�;�W�e_>�Ȗ%í0���`�(�
����k�3����1-��������
��P̈��mq�b����E$�N�MJ�܀%�h�_!Ĕ��lÿ��\���k�A:��&x���s�p.�7�v���!���c��r��r�%"쁋0�!Y�+��ɩ>�k�<�^��'lrE�h����W=�s���z2��8��z�G���w�Z����8o����B���=��/���Wu���:��0+`"�&� ��5�S���ߪ���X[0L�&8����_㈅Ƒv��H�7�YX_�6R�0����Ls����[�akFӗ�����~�'G�
��1�1W��l��R�����̨�]�e}�q1+T�a�?ܒ�6��~����6�O�2��궇���y���M9��KzX��b���� �N�C��IW��]'\0��:�B����N-x:l�7������{�x&N����rf~�Z�O'�S���4��Ũ�@�G`����a�܏�M��+p��O3�~�TB2t_��L�p�L�j|�]���x5�Kw���O4����&^�+Yp��౏m��*o�=b�3��V��|��ĞJ(f�|�V��؊�H �6�/rZ��ٍ�,]�����0�~T��p�)�殄Ŋ��S�����X?Ul��� ����
xH�P1��)0� ���h�c�J?Ѥ�����W�"�[�R�K�kU]s�w�c֜2�G��\����Y���Sp�k��W�#:�K�+���D�mi�;L�L=���Ǯ�Ȑ��Q/_���!�m�9|*^ǒ[gnףjY���Q��r��u��f)z/g��|R\8�������U'�P�ZZ(�Z遬Gs��HaZE2�rR�E��HY�eը۲Q������)�L
|��ρڦ��]��x�����0�1�Q�*�r-�2�*W�e:�Υ�V>���<w�+�Nޡ��� ���{�m�A�\��c-=wrx���$���xΐ弱F���kT�2b��Ͱ�L���Y`E�g��,>g�5�0?�8 c��E*�=0q��f2��t�Ë�����|D�/��w�a@�{�d����B^� A@ؿ�/��yۣ��<�k���UfC)�	�-�u+����k�z�
>
�49"���ɤ���G�i������o� ���,�J
}:�9�6� �9k���#E�"��4䐐o%A��7d�λtU���zk_�텢`�{-���/��#������U��ҥ�V�F�/������n��t�jQ��{MbVdfY����
��1��99w��1����)"K����@w���,�7�l���vI
j��O�%l�J\�}�%�j?2$/x�+��U<6�>��*'%�b��?�}���>�k�B~?Pǡ+��v���,u0�c'RM�1��P�gqq�Nx0V�"��
��]��#�s�,�"%�Lջ�Ze̿{�9����nh��L�`��I����M���,/��E�"6�*��t�����&���&��P1�)��6��p���} ���f't����.�J|k�����O�Lv�v.��0pt���~�gVF6�|��g3�?+d@]~����Q3��^���f�[���2�=�f�r�����u2 ���RzS�cX��2ъ�Y$,z�ȣ��.�d����w���2�u�w{a-�3��ٱ!�_��&w�D�U��oA�|���=�t�Wѓ_��u�/���MR�Tα�>~wu:���'��y�*���ŧ���C�OHB�3���9N~���Z�`)��Di��W���q���!n%!�pG�a�-3�8>&1�?�>��u�KM��
�ѕ��K��,]��2�:I�>+�� Њ����yB$����������Z����& m��Ȁ�|=���g"� ;�]h�Ģ%W�.�f4:h]� <Ц2<�/��cl::I�0#�H��6��������RM�G,�X}�Z�[��ᒵ���5hd�$뗃�&�(����9���м�(�91�9����-l�l&�G�Q�,�Y�c�� ߻���z`�*�=�y�kD�����+�Z�S�2�gH(��#HzY�^RG2�:���ID����s/��U�`ȓm�3�#A�7��H�嵨�ң����*����5\��z9E!�	ʝFt$���z�C�Ť���� �4��\��:�a�}�qG�����i֜�E}_	���z�U�;����ű$Ă��
�BՐ���	Ժ��0�~�\]]�v�_D�U�E@3�!��ޮ�cК�,���ߨ���B�w�*#S��&ݻ�w����ʫc��+V��U2H��K�/S�	^�"���@�skwu���ޡ`���Ҳ�i���>�����;,���d�h,C�>�Z޲^�p��OQ{d���H|7�s����)$�I6�B���Mˇ�B�"[�[b�8�.B�٢)~o��d��1�M�C�Ɂ5���R��aL��K_ �?g��|/!�Y��y	����'FW�EM=����rozF�H3��bҒm��j ��d�VzZ��)z�3�����,ٟ>���?뚅�q:�����JM�w�q���N�I9+�7�ǎ�uK�{�8����z�?(�ȘK����Zi�}\���� d���zS밡��
��o���N��a�� ����@�v�^
\qR;�t�?"����7�O���c��_a:��y�)3`ǻ���l��Y�m��*|n�u�U��>��!������UƘ������#x7uӳ������*�H]=7@�
Ā&�T�-�eV-f���}�O��mu����tЗ����]��u�i~���~��'%�"*���/�@m�?��N�:����G%��3�c�kJ��`ﳭ��o�5-�j���w_�B�2Hos��7\�M��B'���	��kӈ7S�R��<��Եr�;�$A�Z����yb\Xnx�'R�j}c�J^���^����C�R��Y@��|����=�Z�|�%���$u��JH�u�%�oՆ�"Q�B�18'j'���o����r����#�i' �����ؽm��3�v�U%�
�h����g}�-��s�H ��}�5�t��k�m�XNor+�NR����F�$��KŻ[ւ{���H�����ҽ*�R{P��w�m��=�ЬP��.F�ڶ}��t�Yd��d��t�y׽�)H袮b�E���q�v^�(��О�Z��%�mY-#�>�	%KW�h��CJ��CqZ��G zY�_@�o�����ul\ ����'�[u����v���g%ˉ�A�$b;$��m�� Z=��&�Ϙ�+����F� WZh?f�~t,I>{��9� ��D��!��y[� �+�V�#���!�DcPf7�Fˎ���c3��I���1�Nݨ���]�������^ݖZ��hm@ӈ�k �OX�hM���J��N�pC����xu��[h�z�W0��o�W���
E��Od����H0�֝������B�PO}�_`��D�� E�9o�Y�a��i��fa**(:�M1��"�h�*�Z�SwV�x�>p�4��b��H W7J��+V^$o�S�ԃ��;%��=�f�gգ*65�^�� +������dt�|"���n�4_j�X��*Ҭ��mO�q�vV9S�����_�a+��5Bα�{�b,C�6e������y��Y��7F�����'�r�Q������Z����cl���`�{��O�L��k��aT����[�fY ���1�f�&�A[��^��	#?���RJT��q)�F���T�Ք�s�ߙ/�		�	y�#v��W:��Ԉ�QKκ�LRg<>]���e�����"�xާ BO`?�}�e&���x$���T������=W�m��]7"H������3?X��PW!M�R��y��OO��5vZ�T�O�M+�c�n�"�_� � ���G��=+mT�s�u���~M{���\
�}�VBh_�)��� ˷7$i�#1k����~A}��s� U�,jӱ��99�`>;,@y���<kj�Z:�b�eZ�2Wʇq.�U@�Gc#�4��V*P�-�PB�R��|�uh��ր����}����˛K�ȕ�oj��,5Z�7%ž��8����U	X���[8u�b*�m����[��{Z�iS��#�WG��QN]vI0�^��H��X�W��/Cb$�F~B,*7n���"�v���8i��z��x��\ｄ{��&�ٕX��S�y�Ť��gdx�����8�G�{��mI��ju;d3Z����Ə�n��𾟠�}����j5��J�{�~�0pͭ#�?��r�����4������m��9z�oK��k虋���ʄ	�-�3_�C+��/YL\��s�F�����+*~c-H���AX�>�d��E~��U�Z@�<v�U8<��9iX[� �MIaTu��6f�Ew!>�Qϣڗ~�ʅ1t ��6�o�Ж���8�|��i�f�#����9��C��a��Y��+��q���y�`�e��`��ܥ���V&�Z-̚�F�_+*� ���e�Ez����oO�N�t����M��{�ԥB#8f�]�h􅔇����LF���	T!0��>4hXci�- �8���kֶ:.���Z���n�&!�12֙"�]5�g�tݢ������9�I�ycC8[�O�"�M��)·����� AEb�RsGg����G�D��Xc5r�k"�����^����.?�����B�� ғ�_�ϪƔ�a݂�@�;|b�yM�-+�7��D�u�9C�Zd�Di�����Ɨ|Rw�����i���U�d������il�1l���Us��g7%4�z١���D1#�;���#J����<��(�W�+���@�ҭ��7|����(Rp{�?o��[K/̊Oi�A��΋���E��c��������XH.��0�AΎ��}Y�� D80���������Nj��;� ��W޳	�? B�8���f��!\rS��7t��u>"?(�� 1JA�v�!:1; Ƽc����~7���U�N\������,S>�V�e���DǙ�؂�}�0�-�=#3Ђ^�ᷲ.�j4��n�ʟ������QЉ�����6fty�)�,u����3"=���=�/��Bqb%=$��w=0���#����@���Iz�Wz�0�,�]�&�,V�dDw3�'��	5����22f	�3!� uJr�5��m��W��oO ������W7�|�C|1h�I�HݝڐA�}vc�6'�q��a��zD:�Ό�%y8	i�ЄQ�K���k1����x�$��ή��.c���cF���,p�/�[V��}Nܕ�����L��T�#(Y����|N������c��Ŵ)Q���v8G�s�)=�M����8�# PnڹhJ���'=/��G�e�������;N�����|QǺz��&n��9����ڄ��>���<3F�-]=4��#r���0;��D:��5$�?���y4��9p+��u�=�	�t�t�͡�L�^B���l��Ϡ���oK;�����6��<p���eNIL;Ww-�.ld%I�HU�8�Թo��L�9�~�j���$1�O��0
am.v��Sb��w���,{�!���dy*���&�\̩Dn�HA�Rk���MN��C��̮��P�<ÖC�.	�@xw�:ğ��������O܇?�[��ÊL����M���ӇYH�b=�7�t�T�_s�W?[����pk��0/q:c`�p��bC��4�1VG�uY��`nOr��)���]��x�ʹ��&�|���� !��?-���g��}`��2���5���[�a�Q�"���^�4�]����iR����S�06��>�,��;\{Q�j*r���X[�Ǵ܂>OyB�&V� H�U�J��U�,O7�*�D��vr��m�m\�[tM3^�M(��D�"�b�r��!���U K����/���P֞Z#�M)��pe���F7��O~Ғ�FH��d��r���LI��Ո$��ߒ?!�
��F��#%a<�.3���R:_}Y�94e+����f���ǐ���Ja�	�'�S�`<���������}�Cɣ�H�B�������LJ�/8������4�����pq�jg�j��0-]��7mJ�d%�0p��E(�_�;�M�n�"�t}�y���
�X���Hk� Vh�:�k�%��~(�_M�G}e�\|u�?����D�kc�Fݬ?9�KS���!=P�||����!P��P,k��;��8[+�2t/E��}��$���*|Xo�/$=Ƌ"�27:%)
�xȓ��X^�� ���d�k���T����%��,���9�}��$�s�i$�N�O��#9�]��Y0٫ö�ȝ���l}z)Ey�v�F�q�z>��]�7�q�Y�~[@[٭f1��^vs�&�b��]�|v�"t�8'R�D���:M�a'�Y��ʜw"�	�'�$����i��#$݈�x�r&-�e=��:��^��N�碌H�::S�\)�*�T���Š>(BcXB d� $�$�܈��LN` ��"8'�J��]�n����+p����妤�����P�U�r��:2����Aʭ��h��Y�0.�$��/V�N����8�۠'�}�@(����p0�3����c�|��#,�{ޕ�H�Iu�m���1���X��8��",�CS_�G?ʥݶ�,*�Ђ�/er:j�3uw�h#6�߶Ң3���N@�(t�|�g��)��֯ (Vt[J��S��#�i��]dw��� 6lhvɚt��o��8��ɊS��~X`���@�Z_U�N��9ߍ�y�hK�kϦ5I望�|��P�n�>��|�}�w�;C���c��'~�,vO&yE���G:xt�}R�Ċv}=D�L�u�����޹[�}?�E�;�6+&gRx�>�-.Q�R2��X�x��z�p���!��W{j�)m�8���Hަ�=����ȍЗ�,�Z=Y�r�������V�[ۖЌ�������z��U���v��v�Y'u�$�������=r�l#g�Eh(}3�c��_�^���QyF=��,�U
6l�[�L0�a����APg�Lm���'�9��J#��i�YK*H{�G\@*�l$�k������.n�,[7e���z�ݤ����Q��5r��'O�(�-�$����D����d�ڈI-�K#r�R��~��}(�R���Ƌ�`c�>���ەY�>���[����Y+@�@����\���S����-D�VOQ�a��"��ϴڰ���I/	6Q����U."x�e�{�Fl��;yJ��	E�_�PDĉ��ڸ-������6Q��wt�7V_��%n����x��D�-/u�\i�8 aU�0�+���i7�G��|JAJ�J_��-��-�H�W�5�1�ɢ8}U	m&x�8=~�rw����N�&n�ܙ����%0�(6��������_������~���W�p� ie�]+���(���}V�n�����K���("FL��A�Sd�J�F�m#rp��,��9���~���d�}��ӭ4�6�38�P�L����k�d��O7t+>*wf����:�S�8��������#�V�"�Za'�|l�	%�� M���RQ8�_�1���23�fwQ�9�W\xq9��Q��9(�Ծ�XB�c��\<����謥.��D]!��J{YVO[>�ƥ.ErGJ�y�M�������U����:;|H�O�.F�e`�_&�7��=����#����3>�&�L�Dg*E�Cw�����m"IA_�(���o��+����0腕���q�2mg���:7���A
aY�#9���c�b�~O�F}�N,��vK(�d8)^m��&v�FL�<�`�u@�S1J^��/��Rdp��to�Y��ݼ� ���f���2x�*�yV=����_{o�u��՚��2�e`K�+�����ع~Kp��ڢ��C�gXa[��'	3F�c�\�B�{Uo�<��<�2{��n1��A�Y�C���m�w�!���<��k�crIpƝM��Ы���.�'���5��A]tg��U�M�������?�=n�;���FP�'/��&"gk��K:0��6�.4��,���4�%;3ŞA�������'v<7�]�`K�4��c���Fe�5J�_p�2OyY7�B���⥑oQ��o^ql�zl�w����pa�r,	̼x���7�7~�����K�n�v���34���f�?�"�	!�	m��a�ύu/>�f��RxEF-�_4� �d	5[��$��j�^�p���z�Дm^^�p���V�D��ړ�m��'���O4i�Օ��<���v�K܍�C�$W�T��o�2�4��G�]e?cw4��Wgo<���"Y���s2�/�s� �]&`r_�2
�l �g7���[C���q�h�:�&*g����r��h�jRxhw��Aw���3:z�>�4 L͵���wЗ*+�n��3oх�v1>	m��NF0v^��!&�:�BJ�<Q������?p��ڂ����dm�(n}.�"i;o�L������mp�����b?�=�Bt����7;�%p��Ǵ�wyQ�J�nϸ�/��d �|:�U|��Et|lv�#��:+nN;���1���p�ne��W�����&+ÓmǢ'�Br���?������t���g')&z�9uBJ������ui�Y�X�X}@�%�{�~X��|�ƫ�4��W��r���;�oY9j>��B�֊�e2S�?�J38�t�G
��B���v��	k@b�U�PY>n���9���ܫ��p֞IJ����j�JG%�-�F��	� �O�3A�q�q(� ����~I�{V�Ć�P+e�ݰ�q�K�q�"h�No�XA�ج��Ĭ:֐�8�P���l�a�R}�?��+T��rH�մ4�gFɢ�f<`�q@�F���,XD�&;��^�H+���F��ԝ!v��ݞ�O">�tB��ſ�M�.Mp�B��3H5"���2��h�*�3��E�d�Y��0X����V5ʒ������L�v
�n�i~�n���4�b҆�^���<~�_-��v�ĝa��&e���'LPB!n4����V�֌Izӏ폳Z�<\i�s3/��������'�һ����Q��UċSK%:S��ob�
�!��lH��9=Q|�;�=��'�l�>��%�|b'b�=�EO�t��a�=��t�+��U0E����REZw�?��Z�O;J�������v��K����r'�`0Z>W�T�����9������'UU+v���5�y8c��
��A���$4���oM�PR�Mq�d�<�")�c ���3����<�K-�>��~��;,=�����6*6�NC����&*#UrS�^_&�&w�4G�_�0s!XZM ��I6�A���B�zK;�k9��J���`Fҳ�LFXea8Z�[�z�65If�����9.y9��M��]%�b��}�Dʆ]��p���*��V�<%�� 6�- -Q�ok)��Q����2&����g��TB�S�֙J/�Y��_�VZ�,t�ԣ��H;���Y#��|��[��g"����L�G��x��e�;�.�Ѷ�	/5U8�������t��� �I�s��.��4-�7Fo,�Q
-4�٫`����{85�T*r�1�c�E��Zx!Zm��ƌ�ձGѽ�:�ϡ���s�����Y�%�Nі�N���F��"��'����}�4p~u�t:b�E�Z�(����A���t���1��IlI5����
���l%�h�`��E�f�������Z��u��3�e��zPo&9������/%�Ws�*x�"|p>���"5� :���n�p�DR�;�<ۛ�����?^2���:�c���{C/��\�Kj��k$��Qe� h��~V��Z�[X�WyA\�Ef�"*u���R�CjZ 3��ڝ�g���q*��l��/��h�@���G���!�'��z�s��߼�^��ף�[�H��d3펻9t*P�!8�-��y��EJ����L���Xmn`��{[��r��k1���[Y�\
ϥ9hX���Qw����ʇ�xG��t{�9<OJ�Em�DN5Ԥ?�Vlμ'���H�H���|�g<�ĵby�╧�a����A2m�[�6N�&C�;'�r�&r�zͥQ���^`����Q�i��ힻX:�аy� ���zM���_ȟ��&�V��y�$i�b?"a.\�fM%�8��8@����U�{�dmu�Zm�_���S|�>N 'q��LU.�RY�4�GNX4�7�Et@y,O��IE7�Ϫgm���/�2,�Rt}�{ֹBcS�=k8L@͏��mB�V��Z�XJ�sI��Ɖ��rF�B�U�Ue��`�M�>��q��Z�0�5���5u{�^`4 |�,��*>�$⮄A.���āݣ0�g����ݮ�*�����F��j�7�_�<M���Q��Uo���/)0�I�aC�¼��l���Q������ 9So�/�1Kv�;��N��u3(�]�s֑���f0i��p�~G���W�>��/u�P.��t3`d����+x�[��w�|e�nݤ�Q־F�?j������x�>��;�e���C�v�Zb}L{�� �Ě���~��Г�f�uɒ.5�F��B�?��|3��]'w��
�b�\�t�,z=aWI<�e�Q?�.y�1_�rMR����*yB�������'�����M'{q�TX�g,)*"^x�k|79jM�P���#��6C߬�o��i�k~�Y�j�\��Du��Y�}�D��_6o�P�`� ��F5}dx��*��;�Kx썍��'��L>�AI I
�Jj0����`J����t�X�|:�����m~l�^�B�0�����=�(S�=���"��Bf^���JɯPS�	;�)P�0��skͤ[�������c�
7�+�`XO�9�n3���WĮ�P6�1��I�>�N��&���K5erD�P���r%��F��
����6���'F�}�z�pl�5N���~N��g�M�
8�!�eD�R\�3����6��v�i�"FE�+�s<�$fq�0���8qڰi%���n7�| �y?/�Ȗ�j�X�B�(��F�|��BmҬ�ͬ�a˨�D�l��ˢ����z�)Lf�3����Cr5�Z��F"�J�'���	�fE1��6�RX�'�!�]Wϳ�d�~XSЀ���w�?���? 3v�Pr`ηfh0�(�mvռ���U,�F����P�-��vFgJ�V���k&���MP6�ܬ�[o��[?�1-�=T�_�4�����CP�)rpH��6��sn���>�_˱4?�D	a��ϖ�x��	"٣/�&�
�L�����ӊgsl��r��c�Y4��=��*>�~�*h�/��x<�Ȩ�?�Tܖ�Ƙ�'BB4���\0w�\�x{⌊tT?�!�[+��MR��"�o�:���%�fܹ׆�j!�%�a{I9S9�sا7��a���B}����.@�w[u��r�N��b�!�j��\������	ymBNdj��fKΝ��Ɲ'C�v��B���fΙT.w"���c���G��:�;(�QxN ��q�������aN�Y�h��9=?ٛ���o�8���]s}�عG���(?��&���j!�J
��ѫ�D�l��I��E�:��fC���H���� ������F@���ѹ���������e���ߐG�|��5������>��1��Y��m��}��ʶh�#j`4����R+��F*�ʆg���8TY&�c1�98Z�F�X܈�w�����M�<��� �5ɖ�m~�)/%]r�~�᫊,��6J9���ΖK��mR�	2 �3�NJ=�S5"a�C�S+{��7T�b¸��A��߼��zj�qq���v�eǿ�����-I��I����c�Ћ�*Z �S;ts�+:*w���A]or͔q8��)�͑U��B��9NX:P`2Q�����9�0��Y�q�j����!w9Z:Ν[���S�fN�/����%'�B�1����s�J˂��x��XQ�8����IZ>�ء*T��y(�#M�	�5�"�N�״�DxO�����o�nh/�"�[�1%F��4�\:�by�^��7
�lh�d��G�գ��/�tWVi��L����z��A���n�\J't�<s��~������ڔ��I�>���a"E�ɠ�K���Few���n�t�b����}hN�O�u����a2��Ęy��~�X�,Э5B��?6g�'�l��e���[��'vmP�)R�ۮ�+ �/JHYȯ�BK�ښ&k4��57���u����^�H8�Dl�p�p���D�9�h&❄��t�p��]�\Ȋ^W%�/�G~�ħ4�� ��7GY����OG�9�(/�.��������R!w%̷E�F��M�V9�}��N�	�����'���5hZ�i���X�r�}��A8��
u�Tp�V'�d«w��\��J��n/��)떜}����G^�~����5�J�L�!R��sT�����0�M:�,�X�Mv�Rl�5y�����+��{�K�Y���4���cogr�{߲����J;�n0N��MlD�&[�
���^X���|Lt.*�	�}�����w*�3<a�������B�E	�м��N_DM����B�^n~���_�W7�x[�����JЖ��SX;��LPiܭ�W5*�E�._Xh���!��BGջ
�\�Tpl���M\7�Ro��ޮ!ǟ\�k�1�	� $��z�+��|!�p�4�)C� �����'�A���Q+��v���W���I<$Ʋ֛�.Ɯ|��F�!�: ���P�4�)��y� 볩EU>e7e�,
����\rHOi=�����;��и*�#)�bv���VIgB*V��0��i��܏�L'�\��Č�h� �ӽ��s�VW�N�X����	ld�l�&�ۃ�*\oCӃ��4��6[�����dI��~���@g"n�,s�φ����f�4E!h�5�`ҭiC��mY���g|��+�K�������w�d�\e_&��%}6$����Y-�H��O�Q�"p7�R�ǲ�ذ�c&�
����0�����S%�d�N�n���Y�Ntة0v�˛��2<��u��.��%��d�[��i]f���̟�Q�̡) ګ�]igoM�J�O�?���~�u��}~m5�bt��i��M\��R�42|�^g*h�?�`��˕�����x~�'�j�?�Nͻ�o%�*q=c��<@S�ݕ��M��f�<�w�fޔ@��[Ѷݓ,�%���9`�.谍���U���y���[9b�ۉ{��&����{��L�Ϣb���JZQHm�1;U�%p�ygv�~B`]r���i^B�Gh/_���@�(E0:7�͵P��l�����k ϵ͹6N�MHP+�af/�n�����A��q;�0Z���q�h$j�dX���h0�6�H��]HG3�T�����E��΀%�+�����Ͳ�57�K;ޔ��?g�S򶜖|9ϱ�Q�x^����ݾ�~)S����ݏh���Ӝ�=z&p&���.Y ��y�	�Ī���Q��6]	�~�3�j�vc��U;M�2�r�����߂��g�-Y�|�(��;I�`�� gY���*Q�/�״��\��+�!�;o(��3�N����͉��i��]���Ր3� LA}�u rc�	�-��N2;�is���p�nR�̡�o&��'`G.�b
U�,�v�f�G��T�s�LsJ�#����2w��F���A�����<i�����m� �M����ԂP��kY�'P��ZL"J#��N��v˜��̸��
{��>�z����6(�n	�����M��q�Fc�X��Dx�n�	tӻy\&E_FU��I��-X���Z�d�;^ ��|������;6ި�7l��#tJYs�P�E��pO9t��K[�l�}Fv���@K������ ����g�	w�wx5j�& �#��~(��#�?(�ɾ�����j� [G�aJ�tr
��ϻ�"�}����_~0�?@��˥���7Ԭ5J��2�uc�GX�^��۹4�W���j ��T<y�c���^�\��K��TL�c���U߂?��'��������,YF�T�˝��b[f5���I�|�]��0{�� 4�v��^Y���T�c����'je�r����8���zˀ��CIyN����b�*�W��erA�a�-gh���3�QN/<rG]��ϣ�2�ʔ�/_�<�Kg��n8�n��������`o74r;���G	�6���X����-r���[�^��8KI���R}&��(���s�n-��b����=�sl��A���}�?.����/�Q뗶VK����V��x��+����?�����e��'@n'~��~T���he.p�1?�bC;�>���2�}$�>�.;#�c�7���~�G�dnuK4&˲ק�9��f��R[��φ6�H��͑o�A��mK��?y����f^�?p�:�*}	��y�޷-)H�d����@E�����F��.��'�0�h���D�����!<����<�+��l ku�]6�!���rH�8w� ��T��_�ܲd��th{�,!N���]j���b��j�d�5@�<F���{�,���0_Q�4�ch���"���+F�B����,�!�q����;��EKWI�����ml�6�RA��ٯ|�U�0��n�}곐�{�"p���S���1��T.j�G�2Eq�!9�n�k̭y-<�gL�
��bݫElH��?%�a^)K��C��x�V�~�O �ۋ&)���.9��`Jۯ�R!I��jf[	�܄�R��f�U�ď�
�v����P���K�,J>��l���/���!���zqP����zZI���W��כɱ���34ׯ�ϰ9�Eȕ[Y�x6��Fn�f7�]?I�z��P]�̙��o�����c�&
�������<�!��7'�I�Fa�����Y�jl�Ѵ��A>K�����������s#� �[�L��^vsV�w�?��ٚ-���Χ�'����^�׎�������{8�QwD����P�f!,����n���B|8�B�����[��s�>������!%�; 1R]��L��T���$�%(�3yM3���,&�]#����"̶@�ܢ0�ޝA����Vl��Sڭ����+��4U���T�̈́k���w, }\�d�:�80�(��y��e7y��
D�����VR53�WÚk���\��Lh��|��6�w�\c������d��r=��5c����1�ҷl2�0�����x�sc�)u��E�on��ă�$N�D���f�k�es0�!k�wE�kE;zb�Oݽ���ь�x�&�團Es�m���H����o/��Mձ���8V[e���%��j{bl�]P�>`j�u�r�����ь9����_�voHJ��h����o�ou4�����?f��M�`t�$Ҩ.�����S��u��� �	V�?����^Pv�|i�UZ?�����0H�e1���KYz8r�*Ʈ8מ�s�n'�km*\5���nð;hC��e���.}0+�sSa��=�����g�T;���ӤSE�����n��+eΊ�w��(��!�{Q��C%�˷��#3� �0Ai���b����7�?' yBh܃qL�,b�0��{dw!���3a>�<L��� JvU����#�l�
<���rٚ�V��m԰O[�j�?��$�|E��$��
}����*�:��r�B�nq������|��bOX{���!��~�Ѵ�7�S���߳U=�	�5d~9)'�ŝ����.���h��t�J���H?)*�v�\z��U+U��]��֫Qp0��}U׬��*� ��(�Է`���n�]�Y��m!1o[� VlBQ���}������7 ��{�ń
�"�f�p`o���7�"Q��� (������[�xP� =���z�h���c��<����K�c;�&L�{��ew�>���e2���Pf�'�ܘhu~��~,�oI��V�n�ښ@g,�\�U �K��+��N�3� !�M�^"�(E���\ Ng[�������n�zs~���^�j��?{c�CVc(0JL�/��=���Z���&���6�Q�����hwB
k�w�LE���{�?��ǣ\�<���Vϫ�l�m�_Qǁ���~qi�i�c٘�%�L>�z#T)��e�����;��;��*�����6�_��c����,v�5��R�ڻ�}C�������T�M�xwv��_���o�X�t��<�}������O;�!������"r�>G��79�'#A>e�Uxe��W��'T�*<It�&ZO��1&d�;CwZ`���& ��݃�{�)�W�g�
�@~���I�n�9K�]�`�PN�M#kT�lf�=��G
0f���k�}��bw��Vʱ9ü$�/V,���0Y�/�ߌ���-��)GrO��
�
�k��J����:���=5�3HxI7К����P�UY]�@{�Z�ܼ:~Y0r\���GP�f��$Q��UD�t��]j~�Cp�� z��ھE��q��@�kjh�A��]��N�O���-�y��4�T��C�D��ִ��SHc;QR�WT<ǁH����YC�?"���|@#���Q<ߖ���#�D���,�z�d�q�3���WBp�Q�ȁ�9d�z�5dL�KF�E8�F��1��J5QQZ��v+�sH�~]��&z���n5gU���jc���I�4�Є5���lw�O���j�=�8�#�J�y5��a�C���q���$�!��Sϑ� ~]�čR6�'H�xJtм�-���}��N*N:_ 2)S+m��Owm��[���n�T���ZU�1����z�_����N�c�Ɗ�D&��7?ze��*U><���o�
(6���B�b��-��tQ\�NЌ���:5��TG�c�� �bA�BI��v�~&�M#/*�G��=�����5�ƿ���>>�h��b,p�)����eT
�U�&U���3��J�d���^���k6e��j�9k���@r�����3.�j�S4�������o�;�U���s�M@�tE�����ev����u�q�
�4�'
��]gp�O�*	A�5{�������Z�m�G������d�(О)�PE��|
��N���9�$�<�|Wߏ֊����ߊ����e�q��zczI?��f)w]�(��s��l�À�NP|�h��V���c~N��D���B�N5/o<�X�86�C2�dP<j����c�0�,P�ɘ(G���2�)I�F�u ��"�۽?Z�l�4[.T�n�����t�<u���6|��B
��ڐ$?+e�|4��z���K,{�٫T���(n�k]��
#Fg�DϺ�1\T^(�����S�A�Ì4D�<�"i����v����$�v���������� B��v�e6��2@�
%�@��B}kp�N�զ�R*��U�,�&�ۡ�;�Դ���_i֓�<�} ��E�W�z8�)�f�
v��H4RGK�=�l��׼��R�!�I&bJ�1�7���Ckl�	蜀��+q��F���;A�]�e;�����W��<L�N3Ԯ="3���a/i�O��L�_�K4�g�s!��uK"~>�CK@{�Yp��u�� ��ܐ���*?���j8��H�zI�� .�❍* �f�Ο֤-��;8+�ԍ/ Z��g��3Ј� I�N
�e:>�O��!G��uY��`ذ�3��a`�I/�F�����D�N�q��A��O�k`�jl����C�zb�o��ߚU���8��+��V�F� �)�����ū��-��`�o'��o�+"Gɣ�ĉ�B^�\�f,��z�L�m��l��K�R�޽\Ԥ|�d����
$�A����5�da��9��3]�<����}ɽ����]�귆OE�s�0|hpI�f��f�+Y G�8�t2ޘ���X>I0b�F.s�Dꀼ�ٔ����ݛ�T�{�����Z,���	`>L�`�?�@Y�S�'�f��"l�Y���=��}����<��fJ�4�`(�Q52�(���l���t�p�FD�����+м EY�D�
�:�Qf��]uF������i�a��J���'���]�����	��yR^b4y��q917��?spѩ�L$�y9�X~��?rH~�h��q��I�͗pHޜ�.v5�&�1]f�ŝ�R�kf�P���+�ۡr���qu�֤ē�`W^�S��x��y�����-����Jw@%F��sS��NP��'-YD�\d�N��W4@[{���O�h��(��M�J+��������)��=1����2Q/�K��9?L)k��K3�@u�+F)txv�'�M��R�W��@2�4˖�X��:Mރ�=,���.�t��M��e��\&��:K@L��iH,�L���{�\�Em��
���hb�d��)�=�+�_')�*+i�ElT��h'/�g�,�G���P�6l�A�q��������O�/�s����e�����%KJ�H�7-[������Y����̅h��ۀ�'�
��f�N�j{��%���9?�%���)L�i��/�%{�x���a��������H�g؋��skĖ��"�Q/�zD�@�݇4ʱV_�JI��H��&)�@��O�2s�ũ~���3�����Vf�e�����F_ΨTǎ0�URl'|�� !L�{�)����:>�PH2j`%~�~�$�׉4���K�_����dF8���]9��5��ر�
����[!O$d>���ۯp��s�Y��b�]AR���E>�I��\���ځ3$d�A.��n�P@+Vꛢ����5S���k�u��T�
-$��0�^3	*4��X�Rm,4�"�ߧ�� �wق'���w�E���À�FM��y�<RM�W����T�8$�3�d��9�k$�h��*�]Oi�B�D>�D��c�I�>"&fm%���Gw�B/ۚ~����6q�\�o!�X�X�(�لFS^��]����/�`9���F��ኬ��0۩L�S�z#.О�E�}9���i#	@b$���-�֦��g���� ��=\��-�nZX8צ}8�m4~q������z͌�]W��0!��h�ӞU��h+������|������%���~��'��X�;)�ʒ��Cp'ގ<�A	S����I�'Q�9�+_e
P�PZdP����k��L�"�vio�bH%h�d���k�����7����Ըs�o6[�I�p�� ���Q1<���&�c^�j���J�?�v�@o��2�;����P�*8�whF�<�C�=����I��U�:�|���-��(�L7"�
!�QZ��s�s?���Ò,w�-ҰX�H������
� ��h�S����f��4�S���l�XE��W�}���Ÿ���:��9j)�����	y����ʬ襩C����u�����b�4R�KU���bS�Cth�>��Y�,��To�,-ˎNY$(rޑ���ǎ5i���FQi�+r^ V=�1�+N��XrN��=��y�.A�s�{x�Z�>�u:Q��bAP6N������\NIP�~�q͸��:�ۦj{4pJ���א7��l#������6�|X�gJ���[g�����+R���o*�m��S�b'S6D#�� �$v�lM�Oa󸧮V�����y6)!�v���NL��'X�r��vU��.����x�[ko
l ��W�c+�.�6l_��ba�%���Y�V+S�{np�I#��Zm���х�rHNb�K/�ZSM���M��\��Re�sJ�݈V�4�r�	�ҥ(��+DU#P�� H��,�wʬ`��롇NK��㯆GlJ�X0���ӎf"��?�1B���4�/��2���D��/�=�J�$�P�y�υe�眄Ǭ�b1"�7�_t��ߡ��HP��u'��~��K;,�и�-��/0櫖y� $4Tz����);����%������bކ��P�`A,��Qu��L����=����4��Qދ�]`�+�L��S.I�܍�VN�����-n��i$E��x�k"���v�5� U,b!���i�!�z�ߣ�K�-:����'E~iT�5�ƒ}~L���3��̷_q"%��W�K?���8srm.��xc3��TJE#�V�rI�P�r�.e98`}8��4���Oq�����+���_�z,x(� d^'x�	�@T��� O3~w�������
�@`��15�&�������oV��?ZG�t��O��晭(�����e��*+ ����*�wAAO�Y�kC]c�@�S��-g��ɑ~+��|o���� �#KV0���`�S��K��ZD%@������*���[��C�G	��#���ݑM?	���)���&�U���0 �Y憴c��˗=Hpg�_OW�ȩ�v�{hu=y�Y[rh�/����|����Ż�����U�?�2ԝhp���ҩ��I�O9M`O���j��2�`�a�~�;HF�ʖ�\�W�R���H��8���Ɲى����U;S��wn���-��H�͊u�g)�*K�s����[7�&w��q�%[�괋���R�eIE��U�1bS�d5�@ֽ�n>��>���/%�N����樆���F�.�U�\mf�w��:�ڢ \!�����~�P�N,w�#y5���&��7]7�_�@��"�O�>$��#�[�F�x~���4w1?Up+˂b�@�j#Ls{DhO-�nX����\����k��&��OФH?>opwKugU�����T����0�̘��?�.*k���D���Z�'|�&W�]���5/�h^�J��Bz>Z��z6���Rc��x�Q�[�w��l��������|�:O�dOoi�wO�->��lKDlj�KA�N0��:�.�X�SJH��$����'��qn>�
�#�D�����Z:����j>�6r�Rf���G;$��M�)�Y��.��fz(�QC���&�w��ٵ�(K������e>S��4��hĀ��-l���Fm�0�����U��$ҳv��2�E��0|J�����e��ʽ��z8
�k��!�)��o,c�`9�Ȧ��7������-n>J(%�aVYp�ֆ;�(�X��R�ݝe,�K<H4	Ƅkٷӽ��{ ��⻩�(�ş1���6q�{q�i��ǔ3g�x���"I�w���0��-��kd̑���
�R�B��MW��Dp��Gy7�*�ƈ�-��JҺ�j/��[����z���@��ޙ��}��/�v�rp��=s��gT_�/4t�о�#�λ���#���.����W|i�n����� �2�t�m[��	�'�VL4�����cAk�b�l�
�$�z$�K��Ʉ�����ѹ~ �}�LC�f�y,a�m����ف��̣�1��|���YF���$Qj�`�X�W[�����D���ᓽ�zf������F:C%^�B���P�ԝ�>�-�C?R�2����=Hz,���F��E����N9�j7���e�`�ڿ���|?�8*�9K�\���s�Y�Y$o�.g�N��A��]f+ɿ`G���`U�u�Á�&���Nh��,�o]�)x��"d��!hA�5X7��Y.I�Э- Q��S�T1�䵐���=��FН̓�2��O��o(3�l~I)íJ�u�﹑M������n"͹>��
t
~[�͍����T�fb��x֒%:�0�ƴh~��a�n��_4[3{_���OIRaHk7G�O6���{�M����_��~v���yg�� t�!3a4�G�g�r
,e�Z�����t(�1���Ԧ͏r�,T�+���	~��+���С& �)0�~Q�U�Y��aa@�*�j�
u�˧��i��=�B�-������6��%�����T��m��IJ��z�-�;yt۔�<R������
�C ��
r}�M�9��e�����ǵ��@#LAǳcM��߮�����K*�>p����;�m�oބ����6vFHm/��s�kC��v�Ϙ�iV��̪S]iO}@�ʳ6�BBJ���s� �����srX��*�48�E��--㴡>�_����;�S~d0�]��9T��J�k�ZbuX~m/	��µ�����ȍ癋`�Vݟ��8߯�=�)����e׾ʈ9m�,2����U�l�m�8L&7Ԥ��%�a����K{�r���1zN�K̝t[`�����W�BO�2��<)�_)i�0=�l
n�� ���0��L-�v"{m���6�Q�<�����O�|�x��N�S�h[?��q��"�3[����]J��-�_��D�Kհ� ���]���w��(��k����ܙJ�ұ+�V�(��Y�x�]av�<:E���x�&@A���)&�3'�:	_�K��=��𦈻�6E_Oފ�ݿ~���Y�٧�&(���@�