��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|̪��q[�d�x�%O�ٵMro(�t��),����z�}�ٱFq{y�����f�y�gM��0��ߐ�䉽�<P|]]�ϘO��S�s�u��$[X���ޕ���2b|9+ gC��*��ve�9�	�`��2G2iV@�"���w����Yk�^.S@h�5t�`���D�V�d�k��_!+�ʬ����@�UD�Эr�>�� c�[>��A}m%�f~���i��{��&�uN+�����6�lI���d	9$���&k�,?Y����v.�����O�Nx�iz��C(b�9E;,�g9n������Ve��b 8c7J!�)a?�a��Bf�%P���}�o|��V�h�kdQa�ݶT����{^ww�Y�d˟��9��͔,Ǌ��!�~����t���?ȴ�!���a���'jQ���9(�
\�L���!*VC���,�,���*g[LR��t��l)f;&��02�eB7׍��Mʦ�z9�h���"A]�@�Zzi�S��]���U���Ӟ��<�rY���g�H��� �$�k�X���ȯ:^p�9�Ï��-Q��Cg����-��҉B,ek �K�suЧ�W�8�_��U�9�WY-�(�CQ�-����8�ڱ����s�I�
R�l{�Cv���2Z�����w���Ŷ�/��,W�:�zt�V��_�����W�i[�ߢ���cA�!�w��yFSs����/���2LYQث������2>xfy&�^�/{�iS��v��3a�
��g��NՔ��V����@�?���3��%������K��f�9}�Q	ƂW�"���;f��4mAjt�:��w������ۓ��Y�Z����>��<�Bћ�,�Q�I���FO��}f >�'c7<�WqPk��l�F���:}@ߩ*�2!���T����N��d�6y��ة
�|�0>R��|�ƺRǚj�^��M�(���/^��3Mh��M1���6jKBSS(�5V���ᵡA�䄽�&ڙs��9l/��8����9�R��� 3�x��ؾ�U)��{�����}�]�?qzDٯO��V/�t�4��\H���!��h3��{���z���8}Y����Ղ��E��A��49w�&��V�4j�f�/<��V��v�����y�u/��	�n�d^OF���9�F�հH�j`j�]8<��r��&vV�Xf���*޼wp�r�� �CB�:�v��O=w[���%2�ZF�NE��N�!�})���2�(�H���&�Bu�M�����mF��_:t �S<��:~���Թ��>�f�5��r�� �A��cK��u���<��Nξl�0o:�<�����y�V��=l�M��7�� ����Ѝ$��#�o�-w�ذ'���~\ ���x���c��0Q��I��c���$F ���U���2��IS�k>$���� -FО��_� �e�e]&�j{q~�<��B
�lz��~�eD>��$S1��y[�����h�=oF>�ϭ#[ɲ �I����΁�=B��a�0G�AP��ΥdH�|��َ���{,��O��Y��� f����b)�c���d�-�e��0"�~�����8�(8�$��1�\J��@��LZ'.�^L��L�Ɨ� ��hB<�p�E���N�6o��n��(½F�F����Tӭ�;��<�ƕ����;R��L-�#z���%��F"]�s�$V�.S�<�>4C��Ꞻ��]P���:�����?�A�')K(í�h��,����p!練�hu���֪xlLr0$�S�*����n76D����zs��g1�S*�?gx��2���V�o� +n��A[3*X�7l�BeK4bd�(�	v�'=��Js�^��}�~�5��ЄV�� ��^mE���ׇ��.�|G^��w,����Hh~�_��>��a��Bإ��x�OJAm�n�!~.Ǘ�ش��U�J��)S*�� ��y0Q��x>���Z�t���B2�q▭J��;�{�f�[�o�Ǧ��+�Ye�'�^H���!9�g!��&>
�t+�Ҟ���]����#9k���v��[?�w�k�B9�A3��H�8�h� ~ff�7��<�ue֚s�����)��lq����`=j���;��m��k��r�O�G�|g&MH�;�y��Z�ۮ5��dFހL���5p�7 V�|	���/��p�嚺�R�|0JZ�bϤ�ف2�,4JV�"<�x��.��2C\����x�n��~x8c�	1&-��ؔ	�6ͦ>��h�'�6ߒ��386-�q*�4J�	8�.uu�2
�o��<����G<��&�~NJ�Q�����y�Z��4H �?��ۚL�����0�-1��G3����l��p���G���+���^�o��%��rҷ��T�xt����C�sq�0"�^o�Ӷ��'k�c���Iq�sZ�N�p��aݲ��Jp�Mn�Y8=����B�V=�ʹ{A�en���?��P����L6����ow[+����,�m�;?lY�Z�BS���d\ �~k�����JX��ig^]�}/A_bq��L�Rf�x#B�2v��	�; �o�.�AE�
���6e��9��r���I��c�ۗ}�W�݁�N��Xm�r�]���j��o��v)����
��y�	X��	�>�Ɠ�ڃ`ʌM5�ؔ��x�^�Q�=Un���`^U	lc�4$y��
<0����[rk�ŉo���s�d�*Y�W?Q�ť�i>�[�!c꠸6#ج*A~"��?[�1��9�v��L�[��N. x5��b1��������b��a������-�b��|�g����E#���R�/�ҟ��y����E6m�x�m:�G�$�q)��\1����e�ԯ�X�6w���&�S%8Ry��Ov��k��k���M]�q�m ۘ���t,�ke�i����$	�k�C�(|�}���d*{�ڔ�A�~
���=�s��D��R�D*������Ж���ε��w��<���H�0��!�Z�睃?/h�5�G�L���d�J!&�Eg7���{	|�z���В���c9�+�09`��9��� 󚣥��^�Wy���D�?���x����5��������)��ڹt��IRԝUB�`=�2矉�ǣ��9��i����_���5=ZB�B��mN�*�V��xk�K>N�"�B�ͨ�DZ˖fk� B�,�Qo rE�U�g���] ���c��nG�`0z>��y��d�]U��bH�j5),��~ d�6Y�H)��ӈ�t�y�}�C��9�1��i�ƻ��L��^9�*�W���QHo �~i�G~u��M��G�:L��n�+�E�UΌ����X� �]����!G':�_1����6�w��£�}뗅�73��ĕ`�2�f��w|�z�N�"���~P���e�0���< �|���E��8��qw�L1���ez��\p1�J g�B'v�d������& a d�|u�𠉻Slw�9X�ǽ�F	�=�Z��O�N�q��
�9t�hyǎ�XGɧ���kk٩p߾����0f�_7_Gr�T9Ast�)��Ȃs�W���b�u\��=h%��`������б#zXo�R�>Rl�bg��=�k�Nԛ�m��.��%@[��8y���I��Z����V��	�/կ�T�o?`͡.���|�\��t�fN��R��e߭߄!�m[Jb)1��y����ܤ����U���9$��tQg���QZt\Di�2��V 2�2Z�=��R�1�$^�kx��0��5�J@�z(��/�μ.��2�������E���l_��I~�<�+~��c�v--m�i���{�����]����%Id|�ܐ\	���
����2�nȐ
���-�:���+'��p�Q�`�GK�F)ŀ���'�G�ؙP8�b�
x���\��0�� �JJG4kM�7���:3p;_�6�J�3��O耜�2���Z�������o}/���)߈a�.K`�z�%���*.Xq	묞��X+�.m�JâtW��0��3}�Z�7;W����y8U_�U�و������(���	���z�S�ﭷK�a�f����R�8ԛ�$1�b�B�΂���L�5�$�g7����p��к�R�]�		ɲϐ|Rk�9ލ�M�/T��M�d���n;����#Y�R���E%ӓ��~+\�N�}�h�d���@��t��ёaK�7Bm�]�3q���bu�J��n%X�+�iK/���b����*�������U���P*L^ ��z($�V)�М�x,>��;���J��tA���B��f��"����}��$��1L��Tc�v_E2��\ۼ��^u(�2Ѓ�pG��rS'���4�P��l����Uտ��V���V�VXx��9p�Gu��d��?�5��deJ��{�U��⦵��c�<���<�$����`$�Nmo9��0\d�`&�}��8�*��횶 �Ʃ����Č#:HJ�z�}%��g�l
نP��Yj4=}�+�]@y��+����:.�h���[vS�)0�'oZ�	�&*��*���K���B�Ci����6I[,4?�z��k/C���f��
s��pK�zy�-���N˄�d����hX�[E�5N�-��=Q��*��)L�DO����������>Wl�Xc߬y|.B�)�����_]KՖ��}�Dke#��� �R����m�� B��t~6\��H�<"O��b
`�1o���+`7x��<�5��g娦��0Fw}eU�Qr�8 �/���)��o�[�Y�Bi�N�H��^RF]�1�( ��.Uj�;�5��=� ���k�7Ifa��!�.>>����H��u��YȮK�.����s��-8dwꃿ��3�i��J�Z}o�����M/���؃+��p�^@4k�Ò���"�e��^X�6|��oAcX��j;�>�_�U�Kj��k(5�mđ^()e�Rљ�8[��e�����␬�'�l5}p>憓2߯�O��Y�>��唵�����?�L�����lq��xc�~���#A���c+�����q�)�D��b |K������E ����s�'���L
A��:z��V��bK+9���jhY��}D������7U�r�I����n��kK�0p����\<�t��d��3T&P�s�T$t�Ⰺ�zt��7$�D�U�W�ߛ�53�bI� ��Ġ�Ni{7�o