��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��XMXl�M�����}^3H����5哖B��E���d��`�~��u�W���p�n���mg��O.%�zn/��2�k=g`l���6aT�E��r�!�����.kw��Zx����;��(�! ����f���(�9-N]ow�����Y���:B���f#�Et�W�Q��h�������1q2���ǿ	�@@KJaX�5J����������\"1m.��"�@��a6��gצ��h�$3��=C���YK���s�J�G�6�����$)�#76��OtZ��Y�P�
Y�ʮw�|�MF	�z���ey��L��H<g& Sk�*]Zn��j|	r���Cw3��q��=��O�=���6��WT?)M��^��'�����.��;��*v��S��0����ںř�\�Ś�J's]����n ��c�F�G�����;�C���	�K?�yn��O���-����!4R#.a�����l�\f�?��s�ͨ�Ap�1����?k1�;� ��r.� �|�TE�!�!�����̔h�.P���"	g؞���DQskT̀0u-�x7^sH�j�Ӑ@�Ymذd����>���A���n)�tI�5�qk�Ȥ0Жkږ8; r���V�υ�c�9�c���40��UieiT��λ��0���w#F�S}+.
�0$�6̲�lM%��	���Xi�[��@�M9��N��~�`�+����DV�rt����������������l�)�z��&XF�|F����.���f��S����\��p'��#]��C�(Y�בP��QC��n�n7���r���z�苫[=��Swk �Ʊ-G��lJ��wޣe��G��s��D��v�5-��,�lS�;���Ҁ���ռP�慕 �K4��H�9�('�W$�6��㯝�(z@R����r�ô���A2�M�Q>��<Vc�ǁҜ��*~ �f��*�J��ۙ�T;�,?�*�J�o�_���$P]Y�x��&1��Aj{�M�T����rK��<:�d�G饖��Ml���H	�rۏ�/�xC�7o}l���W Yg����.��3�ǲӁjK~��(�o�SGUv��"��ď(t�e1��/k��f�d�C��}Ο�F�}B� �R�C`��LA���k"�⿰��9��v9�~FD8��5�`��O٬������*�|��l�H��k��^X��93�B6�95Ӷ���v��lgs�C�p̄A:����y�{�*1���0b�wţ�0:lrf����E�,
��Qw?���Q3�A-�F:`��'JU� ��e�M�63	֯K�=���w�.�{��*�,{1��A� ���o*�Z�B��3��<B"G����n�gr���Xl��у�	������v��Dƥ����m~Lؖ
7Q����CYVP��-s�B��u��~3 Q�ga���O*xI)��Hx㷱Ć���hv����ܐ�����8C@kW臹�vA�]~�L�cn��u����8��}׷T��y[\-�wD'�66ו���(�b_i�~z��w��Eɻ�oZnQE�	�0.k���q��r�u��N�5�<�t��84t�fpWP��4{櫕��A����ɧ$��<���Q&)�^��Ҷ����3��,Hz�ju�9�E����=�[g^~)��^�?T�_?�[�"�;X��|}��
��=����_�y_��3�>�ްk�&�ׄ��A�˯��E`�)A�jk#���|<9��o)�t�%�n$=ޒ+���*��/��΍��Z@'��2<Lkga�	�C�b�������+�,rU'�h�f��J�ĺ��N�퀰��a_!�G�e#�z��N�pAI�qꊜ�(�`d�j,>���q`����dJŜ�$̊�|B�H�3[��6��<�Z�D�����:�Y8j<䆩�)S;sncq��"�����i{ �:�V�/�fQ�uP�m�؆��&F�C����{/g��v��[�ߏځ�'��{,L�?N������x�-)0�b=C�\��A$��l摳�v6K!�a�3k�9]a`�@b�O�����z���O}��w4�=�HC�6=!'�|i��	�U�+(�C�����o��,����ږ���"���|��L�Z�]ј�Ĳ�g|5W��P�s�d��`��&��*
vh�-�6�����$$3��H�,�OX���6�C Skrl�?�,�萆�4��>���iKe��W�K	,A}��Մ����qV%���ѐ�:޸X��:�������j���A���AD{ǦrD����$!���e�C���w!%��X�m�=��0ɏ����O�p4�p3_�B�����#�eȈ�N�:ƹ!5�f�.C변�(��gf�MC�s�l�=9�[q�)?��o<�
=��06���L�6�
2��V�#�t�F�!�*�_�U�fW��t�ο�,|��5]�G11/��t6�쿪���£`���V���~SI���}Ͽ}5�	'G�	�Y�&��LB��q�`/�`��ۉ��R�-֪2�	/�d�Xٮ$�(�V�91E��c��Ӥe	o���[��*�\���{ ��$�� �����������b��J`��i��wj��N���>�hL��tzk�|������XC�<��M�Ȕ�c[�%0AT��y�4* ���7�ωq`7f<lՄo�PC߲Q���O��\r�'�x4�q:�����f�z����{c$�2����P%�Oҩ�h�}�Ao���G[g�� a|����e5�?'<��b�<ޗd��|��o7����9�=�V'���7���p�&k�Οf>�օ��i�8�rՖA�n��?����*>�C�h��?[������/�̼o'HM�RLZJ�l��۔Ψq�.�w��տ�}�V�'�xa��Ϝf��0�_+V�j�h�	�G��j��� ��Q�Ģ�u��串[}M��Ȇgezzj���~����=�C͝��z)�Y��� e ��2�}x��� ��i��5��^t��=U@2���hZ��s0u�[��q��V�^�9]�G}Rr׵Bo�W-�>���a1��p�r�4	�k�����z.�R�C9��`�r�L,}���,+iϺ����
Bv�X57~�Sc�
���6f�"B�&�m�/��F;�?8�)����J�����n��7��ƴgm����}��s����p]��=�(�ۘ,n�cPc�+-�����/����"L~�c�긥��ٞk�R�2��s�v}��%o��9Ӧ��"����5N�Q������x��N ��)D^&����������/j<�C!�rz{�7҆�,���S�&M��hx����>_�1�C�)�y��ɖO�0@����� ��6��s憼��N$��?���L��6]�%���e97ƫ=߶����<;G�@j��t��h 3�*�C�]���[����c}�h�YDYΙ�+=}���DM/��#�)�P���#w���"SJ�a��:�ݙS�ZT�ΒZ�����z���z�lL���z(W��d��C+KYV3��X�NW����Aa��q�7-�\��K�%�Í\j�<7��i�F4[)�a�\���m:F����__�?�`�Ǽ�["��ڄ �.�(4k�	 ����i��M���B�������P�I"���}��u����1T)��eBSu�'�+�؊��&����{}�t�B�)ۘ�1���
=cX Ď���d�����;I]]�_#4m�I���o�	��S�V?}=��'_i�Tə�8{J|v0SΜ�I��=ޡ�ף�K���P��vn�.�2+c��gg����Q�RZ@5�u����㆕�S~R� \�PyJ�r{����N�`�f���=oE�ҸU6LQܒ��H�İ�����lG*�7T'����i�c�8�����a��2����GGO�W�x��Լ
^�O�:�(�t6-�¥f�Hc�#����Q{|�Z�rO�L�����=�)�<^@���Ke�v(� (hd%'����$f�(��4q�iY;pEY4V�E���K K%3�I)�l��nt�M�;�V	r�|�AD��؊��X�X�NY�a����SII'�a�x��zn�`c���>�C"��l��d�|�єVR�^a!S��@�u|C!i[�������uJ$�+ �F}�Z�b�ϨV�ޤ���FCkF��Մ�]hԯb���j��|�#J��e�hjs@f݊}r�M X��*��2�m�� ��Z[kl��+)��Z�$�E�Vҧ5���Wf�&m�^�ܪ?�?1kg�dc3�� e�$��X��\p�c���WM�t����73K�];F�w�믺s$Hw��4���)["�K���`DD9��k�8�N�B-�ה�]��S��Cu^�$�br��e!�7M���~Uͅ��������D{:�s�y�>�,�4@5�I���	"8�n�ׁH�ق�uF�3��� ���g�p�L$�p2�'$D�K�1�W��}5Q�yj�u@7�5�,}7��I�W�H�,�y}K��(d[��.�>�]��Ul�.SqT��K� W���?�V��re�GR�F�����hq��p �75�<o�҆O���纰�s��@��B�3f���ev��j!�j�rq�k"���q�3�Ǎ|@0�Q��9>���6�m�ͽ��]���ʗ�\4��8S!��^~��E53޼;�:��mTݖ�/��S�H�@	�������W�4�U���Y.�9�Y�u<k����y�cy~�C> 	��l �Ẉ>7��%�fR_uou((Fs]59�|֤�����3�
s�x��ܮ���ҏ��ɳI��A*ko,�)O���.���J�?P�b��/7'S��T�ҁ<���4��v�H)tj���^-�!Xw}���N�`�M/ғ��aK�g8�&dСu�U���c�y�P�y�)�oZ�Pd�1�9҃=������P�6��dh�<
�'y�p�
�y� c(�l�c���]�"�{k �������߼�N�	^c�S�f2u��θ�U��LH�&���7�$MO����d����o�YK�}�t��p���v�<�þ�h1�Г1Ph���|���.R6�U���,���>y{rP_�ch�Fg��W�?b5�����i�ԓ5�p#�7��{(�L�������cE���Z��%�t�1�hO'�![}J#�k[��i\��[kKp�+�~���e8X<6��u��ǥ�"���M��V���9Ŝ�$�t�
�8YX��wW���Jd��FW?�?l�7���F�춋��v[�	�����Պ�gډgf�Lһ�^���A�>�H�|⁊��*��N<���"��M���)�b��U��܉	AW�R�V��oS�a��D����D'�\.�)�? )6�*���o��wN}���K�Y�CbAk+�.#C/�,���.�?����6��gw����`�Qy%s.���d��.�e̻��g�o����.����Va5(�f�ݫH��Ф�X���жԹ�A�R�L�L�̹igX7A�����]?�u�z��_wD�@3��J�k-��S�������}�s���V}?G��C�߽�@�I�;Ā7hu��6oӼ��`#|օ[�wɵ3�%�v�;�Ưwٕz�����Z'k�R���-k2�X�X�"AT���Ɍ�E!�(\J^ǃ~n�����&-H.]z�,�����U!�kv��zQ��vվ�2�/�Fs"�@t3[�X��p!V<�����hi��4��Q?��>�����P�Ҋ����B���j��J�۵���"+ ۝W5�(����5�`�}�Ҵ�%�_�$�»�e��zz%Y>���C����D��~�=��ᕧ��H�*G��y�!�t��@T멷��r/�ɸ��v�U`��]��-���&���Ab����\�3o�4"��Q+$�y������m���[��~��bq�-�	|�����qA������B���%|�#�� 1�K�U�	���{MKk���uF1��n!�(IE5�4���8Mb���Z0~��}������ˮE�E����y�2�GQ��Zj	Ӧ鐀ԖA�����-�L���뺁|���E�U����*[�枫�V���Id����"�"����r��E
� ��gc����0P�7�A�}=LM��y%xx7���@��3���7�X�I���	ţ�K'qT��5��������D]��/R��9Fn�K}���&���cVxW���­��$�(��"�>@�eT.�Cb��ka7<<��D���ˑ��@��������f��V3�o]Y+9i�1�ȂaBZ�����O5���W֭�N��WyB	cGP囐�U�x$�˓�w.���LB%�_��VV�*v6�����O�PIt��f���n[��~�?r!Wg�:����m���D�7i|qn�[?�����Q��龿�$j���<�g�1����p�v���M�~����v؇
���S`�2��h4h	����ld�,����h�q/	��b�׸�.Wܦ�=����U��_��x��x�j�g2������|�)����݊3!��>�#>"ъ��PB��۫��-��/��X�d��lD���>�˺�:)o>� �vԧ��H�P��X�xy������?�*@S��<��:w�&�MdW�q* hK��lM�Jo,C�z�C4�)m�A���)� �O����������Ɵ�g�e�O˙�,��L�d�K�߮��g#�W����/��H��ٚ��N�^�*�]6/��4�{��ק��P���j�6�<S�����f�'�Ks=��z	Ŀ���!i���˽ �!PŌ=Wu5.��Д���/�#s����O~yx�-��ܼ��V�[h�)1��ʊ�$���,@�[���c&�S}?e c����,�O�Ѷ�X>�冗C��Y]�6ׂ@�ϷV��L�jf/`Rcˡ�bkn�l������ @�ĸ�8��%'�"������)R���x9�RNc&(�c��5�5��# +�J>Au�z'EXj/��	"H8�a���
���hlq�8Vf��=��(C]5���C����_U�2c�n`TN>�J���`Z�c[��T$L�E�i~�>�̣�Zڢq�>B�|0/XǷ?�g��(����A����,#�K|X�=����~�f詒�� ���>�Î/G�Θ5��cm��'��G�9}���5��#AS��m�zO����N����Xe��_�s]��tYz��u�Xs�)�ʿ�n"B�`�<w��_.�9s�,�.� !(v���-B��c��
;m-��-�j��\��l7q�KV�h� ��'�����P�9�`W��n� |��[-R�|�j2���u2����O�`�8�a��}�f�@4o����̓��)��=!LUB+�(b�R�a��	ȶnAPz�umT�!�d���ma���yy���4�ϕi��w$����D&�G�a�]���;�!�مINk�¬�R�r���`���%bibu�N��\O2?�mo���f���13�\w4�}�����b�Z�F&Ԁ��mL����ܦ1j�,���xe$9��6�r>��f���`�r�u����T!�.Gȇ58-�b_R��с�z�V�K�t|��S�y������������.f��.�� ����r�lD���2
��j�s��X��)tB����aa3��������躞�3{�	(��1<����>"y��wd�z���U~0�ҒD#(��E�T����G�ۥb���t
4�z%\}�%�^�O	��bx�a�B���f>h�@%��ӻgv�l�[$�
�˰f�E��Å��[ׇ��v�P���c�d���f_Ez�XѵG���
ۇv��dA���n���w��)�y%��H�j�[�vz�ˈC&���hZK�+i"A]���5�|��!��1��F���:�E`lUYD(3r<�!�AC���$�U�Nօ�1��˖b���]�����>�C!Hw�+��D����`���t2��LT,A�,���ꗩu`^���,�%�Ky���5];eUBK�c��n�MG6�Nm�=e��q�-��#}��,7��u!� ^�l}1