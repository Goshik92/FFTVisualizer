��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�fL���2��>F���ĉ�ĴnkL"ǡ�oP~���s2�o>S=�ė��1�b�fN���'��G������1@��\[�x���c�8<6Z~Ө��"�������N��Н0(���>*�V܁�������4�c��W��A�Q��L�|��$��'��%��A�c��9V���g5��' �t��O.�Ѕ=��E���#����a2����������o8��K��ǮMt�����Y�3�ۊ��vE�~���Lߓ�P�p�d	*����)���\���q#ͪS4+2��V�y�`��ϧaA��uN%a�j0!��Qߊ�4�d� ���`��q-�+���0*���_ZPV�d�̚P~��k���)��WL7������H*�n߸7s144�DmL���K�_g(�瘧�M�E���qO�4AiE��~�qK4N�t�ۻ<��%��މ�_Cr��M�'ע�/B�Fȶ�Ä��_.���b�ȁM6���G��8pU��72w�'u��N�-0S��m�A����-�$�A�����w�5MD�B~���`Ԓ(F[^���,�f(;�^"�N�թM{���*YP�R��[@95Ɔv��j S���v͢�)^&�"���?���D��T����u�M8����/g���{'T>����@��G����*<P�]��X�_�L��L<a�s6�����a#&���>�*�����\��O��X�,q���¿��f�Rx����uh;�,�&�
�{JV��S���ђlgƈ�/� ��	�&	+ \�L�$�IJP<�~HZ,7%�a�	�	��ʿ�f��N<�\��*��j[��p`��O����`4�!b�p�$�΄d(!���%M�B�cGJg���[��&�̰�sg�u|NX�)r�$VbdkOQD~6�D�jO��� ���M2юH�m��z\l�܁o�-2b�*�^,�>�LI@?l��R�#���vx5cb�������rч-�$���}��륊�.�Q���΢[(��=�@I���ܽj;Wi���{{��kr{�pY�:5�O��0~�?�2_�P��˼H*��`�] o��Y'I7�Dtγ%J��&:3�Ə�\x|��C��.�0s�-J!5T�g��]��;���@��G���J#��%+���F�+:Y�SP�Ȯ"���/܍^\�"7�g������{z���z~� ?䣄�1e��J���K.�C��RI��Fő{alBo/+=\�!�RDMLk��2�AZQ�>#&���	V/5�bq�|Z����|�,���0Kњ{� ��2�!�ʭW��A����M1��|=�V�ol�����_d@�}��Pw�y}����C�UK�~l��#7�G��꭛�g�3�̹0�3�2.�X�O
�'ې�*� KY !���Ȝ뽚�mkh4��!G�\�Ƭ�_"#Er��r!ĘE���>�,0�~S�Y�!nj�rb��d��E�^\��ޡ �� o{��:4'�4W�S[�j�2�پ���-��"��3���>�_뵟N�-���cr!��
�;��?ɸ1�b��~ăF����4/	��U���>1��je��Ềy��j�o׎�s'�3��I�l�$�rq��Z��uNU���^Lo���C$���Q��,j�6�%lf�FH�k��R9ai�Xq�R-�(�����qN�o���*gGX>E"��<j�Q���8T���j>)�ܸ�@��F��E-����K�1�[ӽӚ�,��h���
��I�:.�hԁ�=������>)��'�j����zi�k��<��r}՞�K���2O�ܔ���^�#��Ԛ-])����W!�Ծ`�k�ݬ�Ert�9�q�:�i�/�dW(���>Q2�o��+a�P\u�idTX�����{Aղ�F���Pl�v�g#,X	yB��}�u)&@&[Bl���=tE���V;�p�(�AeB9 [����kï�^3P�m���<%
97@R�����|��Ɠ�PT�9�K:�ZGN���\er���2���fA��N9�d{�p�a�rR�Ky��J�(�n��I���5$o���� )s��@ODBl;��7�'���N��o@&b��о8}d<&*U��#7�����TVPl��������B��y=�3�b��8B�z��Φ�:+��G�������d�w;�듚R��}q68�2�����E��q]�4\�s%,?)���|���7,|�D�P}g���] �����%פ�/`4nv����b�j4IHᆒ�~���S�:�t`\O����]�E��٪�t���0f�	���T�-F�2�n+ ��C�����A����~��(�oJ_�F�#,�5�q��8`���0�?0w���wG\���&�w�ӌ���`��ʺo絫_LV�7�U	�#�I&S,$ǧ[K�����
�,�7�Xͯ�0-.��`��ѓExk�x��TV��)���$�0-m(����_pcĠ��C�i�N�Ԕ���2zH�Jo�_�K��������(��]����\
 Mj6?����%/�y�<(�DgL3$�	���M�H�O��� >/����������g-�ڮ4N~Cq�z�+O��w�y%�p�>v�17�h�3��f/�t�j%��Bb��*�&��C2�}F���W+�-A��C�R^ "��ۀg)6����Рq$��+v��37Á="��a���Wm$/�{+�W5��*�Tb�AX���q�~AҼ⹡����կ~st����շ�e��W��������ٻS}�5�s!K�G
R��5=�M+�G[�"b��Z�pv��~�]4E[����T�y��t�L�q�L�$x]{<B��C�<�~��Ɖ5�ω�;3��R��<���Z a�J�7��-��ҢEX��'|��{�sy�_�<P�km��}T��U�l6k��`�����
a��]/U�J�PӒ���w-]�o|�{N�YY	%�K���̬V�XZ�X��y��*�eGE�){v2��yLS���<<�G� �$�i�g�yl�j<A ��pEu����i�M�x�[�n%n��/������^W�ת I^�ʉ�);(���׍f@V�g���S��Z���0�����I�(M|=2��]�g<+���[K=w��8"|���� �0�Bf��B07-�VWYmp���5;&_�c��P�Ϗ�R0'��ǌ�$�Ӡ��p2c�&��x2�|���y����/{OiGd��.�1�|mn��e8 fO�kw����5+��V�)��z易+���zϙ7��Tm@o)��⼻���J��ʰ��.1(B��Pe4��S����
>��&�cz�F�%j/`rx��
7���x�i��v���5���il��T�XF�#�͕E$8
!�{����'ժ%���Eq�jF�cX�| "G$�Js�r�f}Z��n\���݇p�
m��������ߙ��o�?ء1ۅ�����ۯC�M,@[���|o@�G�`PEawGSWnjE\����?;^f����7���(��b��/JC.���T^~��_U���f��4���j*x��N�uM�[E/hxC��7t*?�����$�+���^�d�Li��6��9�j������꺬��7;�-��ޗ�"O�2s�9�=��x�sy�V�b r3��Ff�	�q���������ۦ��8^��(�pr�7r��鸓8�2*���?�|	C�=��s��,�{�H���K�˹��t�t<��T���Qݬ�nソ�?#o(���~` �1E�%$�6�-�_���vY�I�.ng���\d!��ӝ����-0�%��k��^���?�sh��g�V�e�!��ޥ��OrNb�NΖ�A�����n���ok4ް��FRI݆N��D�
CTf�TO���r߶�-X1��c�ɠ��u/�AH���A=@/s��DOnW��m�fY������J���2����<r3�L�a�/��m�����P�ټg�:cy�VP����0�\�����9j@)��H��q�`�����3҉A�NED@��_wJ8�}SD�!�����}��:čA�;�0ΰ0����diYŀͬ@%2,UH�";�5ψAu��S'|ٱ�����*�s�=�lb9�oȇ"�<�l�0.�.���l�d�0�F�y/|e׿�٭T>��'��#b����ȕ����y�)��%EQ٭""Q�i� 0;LO���9��(
R�0����:�j��;�K���u���:�l�}�L��ռY�+�ۋ7ʟ���d��<����k��@~��y���Й������=�2��U�h���� {V8�������Έ��I���Y�bU�f�*�hŝ�p�[��v!j�ܦN܅�+g󄗀������i��QWa��	3"��Q����?��*��V&�?�bu�s�`F����\1�������QY&ڑ�$��6� ��%�R,�|�����X��@hdWB�A��=��FG?"-�E�J2���;&����U�S3ޓS�ԗQ/^g+۽�o���|q���`�1��q�Y�t<>W�s ���֎[�h��3��TR�#���d���7�U����˧$i�%�
�g�oLTּ�,c���VP��~U�#��+��?sO`�*���3��s���vl+G+'l�}�.}�,`/p�W��K;p=#a0�/޻z徐�{�bsw�����w,ܐ@���t�u�}���������и�ÜH�3C�E.2��u�4]��der̥����fC5�i�O�5��M4?Ǖ�B?���l�)=��:zR�]�^�=�n��J��?����3�s�R��eb�D5�B��4������+�x����� ¬p^��!�Q�? {��f�Ȕ�zk�7:	�������B�L-LQ�oY|5"I������J�}��h�����1�@��\�gx��1��k%���l�Ǜ��%�q�}6�l�t�c� P7�F<ߜ'7�>>����oU0=�H�"�����E�)���P*���A����$ȧ��79I�3�qo]CfP~-���X�>"�2V�h��w}g��3�
)�},?��2�G_Dଆ����e�T0�׶�E/G�nO{�+J��q{��4�JvC=F�;���k]�M�r,^�-���A�W�KI�}+g��{��-�JN�Ϯz�ӑ�v&k��T��w�`[s*��E��0 Rw]��ٱ���*kd��*A�m��dI�&�w��{�N �1Q��� �٠�MV�dk�R ����?!�)��;���N\+�!=�ė��!�:86'Q�-�/q�]=(�tL�u���Z�V�dfM�W0�:�<�=�ۑ��1<߿�"�B�>p��W��f�U�b!Ub^z�?��=	ʇ8�����sz�g2y��E�"�)׮H�(.�R:;��eٶ��3�p��[��2��$ۡ����,{��p]X#P����w��%��Ӎ,M1���/�x?�Ӣ)�P;���BI�8ѳ�p�j��h��N�i����w����:a����=�m�)�d)C���*i�Bd1=/eWh<9J��)��u�m�{9Aq���y���>�H��g7��x-
Ҡ{@ޘ��[rt|Y2_�F �ئl���Z�e�;r`�gQ=L$C,�n�'1o%����:sEȁ3�|�s{ �uM��fR�anj*/}�	�J{[��W�^��RJ�5�"0����q��W�t;�HX��'#�&x1�	�]�m&׉�J��������Jd��C3!��f!n�kC���`�x(�R`�#��.?��Y'����Rl G�b�K�ea'���I��xG.��F	�K�nS��Ιa8��e#k�@"�,�՘���:�%�m�ӃoH�5�\���O�R�`O�
n�l������M���1�@y��Jy�ӹ��s/�^��c�9Y棅Za��y�jz�Fn���0E���k	�� |�~�&�Hp�jW�J��͋��U~+ N����6�b�:���ֺ�W�F��d���m�� �H���~1�����-MY���4���貙bb
,����������N�U�9���{�\ٗ�RP�׀�Iw���/��8�m��oY(��GRI2J�S��P����0(S���7�K]+��A���m�=�Z���ѷp;��B�M@�"�z�������Ôp���wr�_�<by,�H�e�=#���dX���axO�\h��J�{߃��ےS��2��2�Q��/�d��[��
ة"B���	Ԏ��\0%�X����+L���?(�ǖ�u:�f��C%߼�� �oC	F�Xs(��≠ �B�k	q���ȴ޹]�z��H�׏n�|����cP+,��7�Q֨�-���ڏ&�*`r&�>
��:�j蘭F�t'l@�^X�+�����#���*4�my�y�wCe�ř��O#�mW�@�S" �U�5����T]&���@�G�Cʿ<8���~�.���!�(�6|�ȁ1S8ps7I5aU"�^(:�(-Oz���=)��e�F��M��gKJm�c$Փ�C��]|�:Fc�RY�38���H�����\���X�J���l�<�;���?z{$����J�M�zߋ=�r~�'��|�N}%>��w�U/x6c�D=��?� ��fRRx��1>�C��Ǔq�g���T�:��pLY�Y4����yDW͞����_��$-%M��C�WA����7�N���˓|��ohf#>�#9U��j޳s%�oٞ��]�=���>˱�G7���~p�t63@j��M?U�T#�4AFk}Ĭ�_!����Yn����e��ڻJ!j��}�p�:(� �����0¬���%�~�u��Q��=u�LC��O��hd���N��u�)�P2�7׋��y����B1�]�� %�g��M�Z�d�z ��^���Z��0 ��ԟ�bY����#�ց�fQޏ�oj<_�Q��?g����jw}�C��#ߨo�b!�GĀR��hPd�G+A�ᒯ��hO;dJ��6�ZٳB-���H0�o� �g�Kbj�2 �T��vy��x������x=��X�E�p�;d)���ZK�G�����Bs# 3�B�
���/�q7�[���&~�O�D!��<�'>�bFO�83��,��]�����o���yGk�G�� �����R����[PH(U-�i���M����8 #����b��� |-���C�W̆x��#�3c��C������PZ�}����3�Z�`b��*.���ܚ��������Wf0}��B��K�Z	*�uDε�5�V��:��l5��ng�2��oM�%3��^F��(�TI��Eqr���`|�+B�W���Q1�E���A�I#}c|�N4��P v��G����X����N��l!�S�Ml���>�`H�
�A境��U߲�/�,� e��<?�L�2��8�h���DׇZ�n����<+U:��U�����\Dc݁��������`��Q���R���r�ʒ�~σ����~�g8��>Lv��5D4�t�~c} O'.���Ժ n�	:Rf,�L����S6�4��f�Z����"�zCA��e&��)�XZ��[�s��/\������4 �K'�������V:�η:^�f>���$�O��R���ӾE=�e.,P��.P�B-���,�rW�w�Y����&��R�h��2-4�����n+�kKE�	�m�bSE���9,�� ���%̐��Ρ���f̤Yg��#"5sp�hdQu3q�!�j�l�_�Ĭ�����:5��ע�q_Z�C�wG�����1� 1�58@l���wسf�Jc�xF"����^`Qrd_Q9$���4��FE3���c�@I�<:7J�aO'�^mBsN�͙�DԢ����]?͠�k�^����Hy�Hѣ1%INA�P�W��-���dK�������!|K����Kj��+vRd|�A�ɫg�2x������+Y�W�Y:I���+�X�-mR�����O~����e�����Q⋞�9�[���o{�IO�ku9���CK�rX�?_gT������L����T�/�1���O�<14���)X
}����wݜS��A'yF�)�P�⾀�0�Ks�ǫ�L�OU����3{��&�y� {�_���W���z�����8�q0T����<D�Qr��	��ISn�b�뽡|P����~����c|����\�E�c��La��O�M�^a�2�Z � 2���Y��=���d��ч��;�v"<�~�]��O�u��v����%KS�9�M໋��B �+`��u[d�O��+����,$�m/�_dZ���u���7�A
����z'��������K��m�� t6��k#�8�>�U8������H��0m�˞����7�� :�DDߌ���b �j>*1�X���Ē)�����T�"}��L,G���,�4j*P�Q�0��뷹�*i��g�!���w�
�C��SFI�~)'"�*B��A#0�i=���)U��1$*ݤ���3v��˴��8�ʞ|H�E7�@��O>��N��2;dA���h'Y�85s�䜈J�t0��^d���J�j@O�XPO�D�*�ި�G`�C��<�޲7�^��J���[����3�x(j�8
.C��YX�T:(���0��¹5�^=C[>Rt��^-�эL��IX��Z>{+�\�"s�ې�:��]�6����eh��݌�wu�E�Jd�z�]�g̤������u[&_iz�T^MoZF�v�?��!zp�>ĝ� 78!#�⑵D����-(�