��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>%��}w�K�.�TfxJ<ȒEb�����X����E}'RN�ݜ?���B(*fP��g�n��(wn���`NO-�v��&ŉ�G��|�n��s+1�z��0�!��|(��� �Q$	�sT��:�+=Y�i�g�z{kҨ��
�$U
s�SQ�Ɓ�jO�aEZ�/��Z�h�VP�ʟPD%�%Ο��L�i?W�8&".�J.̛�ΛpZ�࠯Oc��7t�-Œ�/h3ݏa燯Mkx"s~2�ڄ�Ӟ� �C��y��SP������l[�N���9�4�#7��HB�-�vo��b#V��9��Q�|�8v���i�v�6Xn-<�+D6W��@��PH�M��,��4Wdv�ԉ�F֧���(~k/�@N�:�Á�L�9"d�e��Q�ɗ����3o�w�ڛs�9���)o��X�Z�O?>Ju����ٱ� e�.���+/$bb.#a�A��E.,&����J�f�� XQ@6�z
c�ɻ~$�∤G��e1�79[I�H�}5�!�5�h�m,/���^S#e�9v@D(y�{D�rP��Zi��X�}�:iM���Õ"�Bܐ0�R͕��pt�Y�}\�z�����ߞ=�u�,��]����HQ���O�n���ËN+�z�;݊��w@X�������;8w��	k&��(2�Q��}����m1�o���q���GY�~��,��?�B7��q�_�!�I+�����8mD>rC`��Đj���h�/hn2�-��O�|y�f�i�V���.�Ӱ�`9K�t������r|-�Ӻ��
N����y�\��Q�	���Ӷ��H<��v*S�Г�4�P]���k�ue?���	C���^�c�KJ�y�ǌ����I�f޿��{�%��Q�fQj�>p[�<8���򟟡l������9�ð#�*߄���^�{Ϫ��L�u���E�O�#$�ߠ�#��4� �'R��t�P���V�n?�l�-�!y� w	��lb���v@�Xo��7�Y/t]*;y�"
�dR�뢈(0��W[dqF�'!Q�Ñ�`D{�d����l�<q��T�����'�*��Yl7�,���l�`#�jPG��h"��iќ}�5��|Q�a�i���"E��,�� *����k�4Z�l���k8��I�|t`�ݲN��
՝�2����t�J�S�
���%�3�!����76���ü�&SS��w��b4_p{��O�<&aL����YU��G*�j�®OU$��xD8��FA�)�	�ҁ풓6{y�i-�9 �7�"0��3���.��v}�7�.֐����:��B��_�!T�-��#m�!���ϒܓ���| �?�ѥM��c��y�
m�F=Ǚķ��ZS�e)AUWq����}�A���D��,T�6�TVv&��f�p� �>�D~*̕�P��h,Q��w�Vs�w�.��JGc��v�٧9�!Px�B*�s�޾���ѥ�6+�חhg�?"׺�].�!рF�����#� �6S��=�aZ93?*�����i]�bI�<�R����ŷU(�BEV�V�bT^/�����_N8
���}����ҒX�DP����˓jF[�E�$�Qb����G�*�S��;�+�7�)��e,T��ɣ*Ioئ����]���(�R��k�M�!�h�h.��ʤ���
�X���~7YE�f��E�A� �Ų-��Х���#"���Y8��E�����W���J�k�c5��H��A��1������q�L���v!�a	V��\f�_|��2����`щ%R���h�Ҭ|1]�E?��i��cȚ�`��n쓺�Lt�#n�CT�0�[5_����`�:�MK6�W�f<�����2�ө��DN��%�ςJ��r�n�W�[w�Ph.<��s������%@V,��Y�`�tB�\8>�臱���r�<�+�mE!|��XF��*/�8��V��\���2��D�����w"O��~@�Gpm$��m>�}�p)���'����!�a'��mtdK��!��N���Y�D�>�\�&�Ve���(̩�����n�U=�a�v�T{mD�s,���C<|D��c�2Kn���8�FҤOEV@ć����y�fč6fQV�(�s۔C��qn�)��e��F&i6�Q(5R!˪���k��a�K��6晥�@�ĩmՈ]�sR�����A�����ޤ��	g�J��Y�� /|�Cd�I�n���B��=Z�j�wi�ݛ�L@�xU)d	UBwn�U*	��v5�/��6kߨ��b����#t��lT�xԼ��e˄�m��-��G�T�|ܦH�{�>���`X��t���]�vy힮c��aS���z���3��G���U���?�
�����n9��[�os��d�z�3����(@��]�rz;U������Kg���i�D$kw��yPT��mA�gp��(���v�D����"�hԯ�N֖����z�����m46,G_�`٦l��EVy�m�F�rS�o�͵�� ���:��v]w�0 �a�>�C��&�ZFm	��a�+4 E(	��*F,�g���k�s͈��1ͺ
{����<۹ ��Z:�V�����z$E����gBX�P��JGD��e�'��N�aⵥ/x�3:�6W�a��Yy�v�8R%��u�t�hSFw� k\ǝ�c�ڍiF��Y� ��sv�ݠ��ԉ�s�4 �1�*j��HLj���UVA���h� ��o}����4W-8�N�\���֏ѪV+�����|xl��a��^��ˬ�zgZ�V@��<b�t������TK�y�-�iVN,&j�BuV��2�{D�*���|y�����x".��",���)���"� ��N�����,:]�h�Ex�=0#��'W����c���k�D���dk߭�w�8��x��9��map�����������D���22��2߆��v���<8��/	`�Uʰ�w���)W�b���]֕ӎmг���$w��*�;��G��nb�2ɠ���/��"h-cC:����M1�`��#hL{�Ybqz�a?���D�\���L���l>~���R&W�*��K=����՘�v��?�w��!��3���'h�+�h�M<�>�],���wA�PF@݈N��S��3�}������ߥ�D^��D�H+��<H����zCޜ��2�)5���G���S�̀��o��S_���{���"m��=�xǃH��V$���
��c��Wc��~�� �.��y�]���_�f���{�������������;YoG��E�Ͽ.��m{����:��ކ(�f�Gk��T��Nb�XD�,�'d��VM(#]�0�8��|�b���FFE��	�=�t����"_Eֹ�����$6����!������w*��������]6W�����$�h�x��jRU���On�Px����p�o]��Su�\)/���B#B[u�I��=�
����iZ�zW`���WV +��Ǳ�9����B����cJ���8�~��'i![<�p1|G��,K�_2�[V�߫�ӄ�>)�|������/�PH�K|�N��sFo5_�0wn	k��E�Fͨ�?0H��ȷ֌p؄d_�����a�}�ynuب��[eq�:��Zr��]�A
�ǳH�YZ2��U�N���	PV28]P��; _[)	!��\�/��A�?�7D3�Ql�����0���a���������~�R}�R
(�0�bmt��t�cw�2R���Yv<E�z2�۸��!�/�]�����Kc�Y$�:�Nu�Ӳ\ؒ���}���s~�;�v�ܵ�O��䌇D���I�+o~΢�����,�*/�Z�
`;Y��j�n�����]QL����^J�dE����n���X����~3Y9X�I�׭�C�чZ�82#�[h+�!0Т�Έ5G�]����0�rms��B'��mk�u㸯|�X�է̅�`(��|@pa�x/�-�%q�5V�,�F�o��	���(��2+�$T�sq�`��!n�g�O|��šI���􋁂I�c�C�����[A|'�� 7����f;|Ȅ�[<�$A��Z����j^�:���K�:6"�3v&_sjԠJ�k]�U5��t]&v��3p��8����Q-��1���<��d+$�Q�Թ��_�6Y��S��7Ҟ�m�*I����V��p���h3:�c�M�9�Q�I�Z<t��3��-�i&��6&�i�ﰕJ����zd>��T?v��Vz�p�x��{i�>�4��l�۝������Ҙ6K��Xj��3~ɂ�)9��4�^|��X'.S_~����n���B�?�*C��wь��=4"���t��p��lX4�L:z-�Y��FU�}!�B �>���kbE��8���|!����Jv�f-�))p���>	�[��c�5��bL�2�yew�t�؆�/��>��6#=�qi�75:�0bh:f�4���<�~8C��1�q\���a�Olq75]Җ@N�"]x@D!�R�:�Pp��@���k���D;r�#5�R0���m�h���_�]�hv���)G�\"a��fW�����D�����[�řH��e���:+�"nx~�e$�Jpz33!����@�i"7o��W�K��Z�;L���qdx���&��c�;A��
pjBn���~�����T�����{P��<�'�t��g�\�?�2T��F�EEؖψh� �X��
��`����.>h����P^p ��t��_�(Kx�q����U�����2�ц%H�E<���rŭ�;��U��
~��HL����KiFy����!1wF�}Wk��i�/����-h�ݙ~��X�'��~dF4yl�`�[��QDՂ��P����;0[���G�M��U\�5�fè�U�S�U�N�C���_��}]�kF�R��F}�鯕�u�"�Ũ�K��dYc�xݓyN�#�hS) >��~���B��(3J���a������[��	{�vd0ʐ?H�S�,�QG�;F����#��Q�$Q[1���ig4�2��(
��^O�P���n!d0x�	�FF����t����d$�J�Vv(�HKY���2l҇�KYE@��-f)%��y���Ω1�؇:�/6�f�h����}�C�0�>MK�?��+]��q�_euexA�_&�����#|�z�n��N��&�H�D`��[7�� -L9���Ch�:u^~�e��Bq���+WW�hE"1�|�\1?��Z}��S;U�:�2˶�-���Dd��6=��\kc�R�\s��:3��͸c䢏5쇯���:C�����o`D���4��!�̡-L�O[��XP��g�����NW{o�z���m�1�7�`T�.��F��M����(P�<}�|��M�;^�[����ΔY���l�`�a�n,�yFs�=��U�o)ja�����y��xZ���f�cG�y�2!ܖ�|��׼3 B�/��$��dC>o���Ge�fW8��w�����t)���U��S�Tu���iZ�c,���^~�h�crm���Ʀ8_���S�6x~��s��)���5��.G�ؽ�}խ�yd�[R�2��ߨ�{UM�!ƫb<,�?H����j�랕-�������@v�J*��-��E��ps� *�ؽ��M��_��we	�FK�������8(��j��^���5`���G�zi�O.6���.�`����o�,`&Cj
Sc�Ҁ��w�1n�G���4"�ʶ�r4�ݤ�2x"e��>A�'������ii���YP�L�B&p���R��"cך�(�+��-�HQң7;R��s\��}+��K�b�S�x���{<�@G�%&+퀊v|����RkWzys�ɝ��?�z)�P����ۈ��69�!�qX���3������U��v\���o��(b��Z������ިҬ�d����]>d6���B�e!�~���Y�-�Z�4nҭVG?�]郶/�VԸ�x��$�ύ�f�o����*�����ܝz��q'�{��m�f3[f�Z�n�?���o��f��E�:sP@�'"f�!�FDٷ�P	���|��,�~ߦc��W!k? �j���S��)����4㈴��zG��;)S!����0����Dg����87kzV��ת�QP�2ޭW��Y�7���7�g` \:2�*�t�-Q�'w[��\�]袋�8�i�!�X�y�f��l[��o?^�3��A��tht���a`�
ljf7W��/`�����ċ}I.D�����X��k�\�F�.cbj;���Ԋ��mv/I"�x���l��,�7�/�\��H���fM�DT#ڃ$:dR謿QЧ�V́t$	�����Nb��	�b8�h+��� G��P���^)�����O�dK[n��	h٘Nd������_�Zb�lx0I�,R�,C����j�ۂD��u��y�? �GA�M�����6\W0�J,L_�c�����޺��>\ �/8e!���7��embr>!�;n#��4[��� ��ɉȬf�DDy`U>^�֤���8�D�V��^2Q��B��.~q�C�krѥ(u�	�>/.*��ht�i�w	՟��}7�C�bo�O�*�G�#�PC��W@�J��S�ueҎ�wU³)꿆��d/
b�X4Z��@��^��l��]��w�q�<R��>�B.�:��J�� ݉^�b��p�2?���S�i9�4������}�|a�{�PP��i����*�("[����c��	���Tl���w��NOB�2>�t�[Cd]�+/X>}ŕ�8��^o��:t�ui����1�M{�vj;Q%)g��(�Wg}E�K��%��=r���k�v�Mn��1Q�DYu�M���zh����)P�5�O_���,�iM��֫r6�X����<���_"�E!�y�:Ƥ�^�$7�W�T.$	95A`� I��O��Yn�Y�[�������a�b�mHů5�[\zs����h�)�'*/���%�
��W7\b����?I(!vl�<����R�r�	!)g'�rBj��]��`ȱ� ;J�6��8�����ٙG� �+˟:Q?}����nx�VI'a>DW����u�Z�P�'Äs����\f>=��tW���4��K�|gS����Y~�)���x�d�rq��@fפ��,�@�v�ǥ��N�IJ��bW��O)��N�y@&Pނ	{+���������� �
�r�z�9��6�{U�������sd����B Ƽ�7���\���D�|�S��mī�l=���.��sR�誺v@z�g�Z�H���
T@���;�n�����*z�`��7�u�{��M�1�N�&J��M�|��5�w�r�)>�I:�#$�}�a�����Z&������B�S7�H5�	)���.�x�3]��y���n�'"��N�L�{����U2�ލױ�e���'G��l�B���l��l��$ :��5����ʡ�5�������%�<9k����r=�H�}Wo��#iM�~v���~�׾�h��h��+ȠK��cJ������m�a�!ruZ˲SS�`�&�DӀ -m��=9h�H�w�.�ƣ5���$���T"M}<!��Ԭ'���_ϰ��l����0�p�$-L�-�λ �v��L�� ��u�	-�|~�&QK~lqX��_� �:.���o$�ڢ>�����V�<2��yƀ�2�]:��\(F*X�~�G��4�.����y8��f�Xꢚ>=7�a ��~E����`�����q�m�d�~і���c�=2�}A�?��YH��کԪb�������/t��G���f	�i}�ߩ���ٌ����4�����;�U'j�58I.�_�j�Cu l\��\����k����9s�`�R�;D�$BxL��O���<��⎪��l�{�y8���و_�%o~4W#'�Jw����&�H&�l�qnǾ��x&�Jx��50�� ���I%���cr�K�X����*ĉ���J��1���.Vm�=m|6e.ĺ�C/!�C��2� �e8��\¤{̑0�J��]�u1C��_�ŌԦQ񇏤�NHq������ ���8��r�,��e�,d�-. y�#�uz�E���-J���ժ6,���C*V"�r=�3�4��T����(S儊Vq#F��+m��K"���b��T�V�$�vg�n�
?�6hnG?�e&�mo�"�hBDS�"��D��HU�&�e��;N���L�y��O4�-��� ��̲��OxZ�W��u<d�^j�- ���qy"���W�FzC��]ZY���z?����sf�-�����e�7�jH�_I4�O�|�G�����y�s�>Ͽ��٠�qR�����g�{f��S�%V�_,�2��@7=�Z!��ܣ'#H��qqlH24��\�|��i�?i�tl-��N�]�� �E9�k�����_��C�wig�랋1���"�9���μ4�K������ͫ����g�g��{����Uٝf�3Xf,݈�����e�N	�,�ڣ��LX�ƧM7ډs{%�J<7*��D�F"3l�<�w ������/�#[ţ����I"��l�B�'�j])�w�%B�d։�/p�L.�L*���J���m�*OG��XG�X+�3=���\���Sz9i'9�Wۂ���|��^�u�fJ�i� ���*�[��%�^/�bt��E�|<D6�h�TQ��@�쮪\���ph��u#G���?���4�b��TY�ܨOO�/-	2�Ӛkd��7�Vt¸�2����ꇉ�2A+k���Y,�g�C4e�����R�۴�Q4�25Gȡ�����'�9qj�j�,c�6QM$ɔ�!�et����MGzN�er5�ik��� j��`��#l��OY�����:1�M7���kX��J~�F[�5(�1�m�:�W�H��3���v	(�r����N"�rCL8�w��J��[V���q�n�Y�gB�;g4fl��R�:j���#�򎅗�V�3j~�"ä�r��/���w�q�L�E��?��P�/p8��� ��h:N5����T���J'�cŅ����34��Jԇ8޺?��~0�}*rn��"���io*�����YjY��0�l��4�ÚU�@�gQ}��^v^�H�3t��¥K�q�Z�!�r�)�xmҧZa�P��W�%V=O��K��sB�1�6��JHc؆����L��䝳���xE���Ŋb{a{��.���ΈM{���������H}����'S�SP�BI®�l�rz&��&>u�[�� �<�ɟ�
glϹ�b��]u+e��3��?�ڤ��J:;�QU��6�����=Q(�cv�a��u���Ju�1 G�s^,-�~��qMy���!���[������U,�э�.�|��~�<-�zm{Sl&�`�E����;�;b/@���R#H͜�W�Y����yf43'���YZk�)���p�0+�~��qHOW�(�\h2������3�w;�����|�,n�����հ��q��������=���^|43�K禾�-�	��CÅ�����n>��\ѱ��������ྦ���k`�v	���/��{�x�}P��`�Bsʄ� ����.�O<��X�;m̝^��BB:YL)��ŕ�G�7���P*�����z$zX���E�-����V�.�	�%�`��o}ٛ4����Γ�����L+�q�D;��\ȶ�������u����osF(�����=@JY��F;hk g�ɕ���n�آ�����	>��m��΋i(��*�}F����}x��ҩ��kB�5�rF&�TWo# �p�<M~��7�Y9�V|=�%+T)�Gn/ʦ�u���wY�ݾ�Od4���3��լ�`�`�p�����6o�j�ҍ��g.���c�t��F:���ꨞ`fj'�C�7/㓚�?�r�P!�8O�Lઆ\٬�Q���+h��+�/����済�H��x�-�2����Ç��5!�E��4}��ﮱo���~Ǡ���<���G�~@�|!j��9�ёPj����vl#)m��uز��-(:y�ߣM�dv*c�(/�*��Cq#dk��2N�"�1�_3(����QX�yl9�h��(�Q��ԛ�x������sq�����A�38�1ΥШ�����hgX<>$)q�\ȣ�\qb1S��>�)}�{��4A�&g�L��	^{FZ?xIةR�؇GE�:�����j�N��nW�|�5����]X��}Y0	�9�b�\�GH?Q�{��}f�q��ݏ%�^0C$��{.�ѫ0Ba�M�X0�me���Y
o�B�����d�v����X��~;��$a�J*�Y���;xJnP�%���/�O���A	|�Iz�����à�O�0M�V�>���İ�3�g`5<yDߞ�������>Eb��'�;��4�:��+���@|R�R�|�G�����g:Vn�!�`��ɺ_��^-�;���
��)���FjP���@�j_�����0�>@��d·�	 ��̫�P���αW��I6�Q��L�v��Z��(����L*���W��O��#N5��^���K�_���c� ����]���jd�&�դ�nb�ಶB�i�}4  ߷l_{�6d�IF	���峕�g,�h�&�B�o'fds@�Fl1E|��)u1��U!���׺r�@=���:���j5A�4�{a:�e"��#���2��#�dqܥ�f�މ���E�rp�@����*k1�zc�k
$��$.={ �j_��е6[�i�;�ȫ��~#����2�1�'/p'z<�b�YZ �@p��GxDz��?��s�L�d���������VG���9��!��\�^M���C:�h�ٰE�n�1��'2?O�����1�ﵠ�+�,?��'�e+�覤���- �*a"��-��R�>�>E��Q�!���R�m�U����Tް_��}�ܫ�]�� �qr���f����d��	8���ӧ+E$�L�?⻜�ޙ���i_��<O:*��2;��-��l��q�t�P$w����[��G`�a�D�}�5t��m�q�I˺Ȼ.7�c�i�b����|c��e��,̰/yp_������H+t_;��2V<,:km��[������8��t�Ɗ�Bo&,K�	[Qʑ�^��Rg`��!K9�I��z�7�n���L�W�Ԓ�+��zU#�p7���g�ȏM�U����Ѓ�uP&�u��A%���,ƿӵz?�G���Rb�Tr��4B��֏�{��C��>���D��$����B!�Mt����zQC��o��S���Q�س�֡q���7�P�5~����/����Viꋴ�5��d