��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]���i#���&6�_Bq+Vr�Ⱥ�,����P��#�pa�G;��w��Ϸ#�̖=V�(�������y�&^�oO4z�6��;^�	��?��܅dg��N�CU�&ڻ���%��h��t�P]W)6�ro=:��Ⱥf�R�%��s�ry|��#��<H��\o_�zӼ�5�����Ӟ��w�)�k�I�5����`�3���4�1��z�����Z\�� �a~J�����ܰ=@��8�7�9����Z�n&�]	zv��5�7�R|��*]�*�����&'E�5B��!b2k����eӭ*��ݧ^V�;k��G���l)#~PS�$x�3Lf�Pm)��f�;;>z�J�La��|��߾������q�1��h�ACI���Y��fOD3�3��TG>a̴m�瓁��d�l����Jal�`��jG�� �FQ�TH����Q<���܅�Y���#�(hc�"�l�J��%URm�׷\��aa�st�&��z��`�,�D���i-Iٔ*�+��ϺyN��A��̧�\�RHϠ%Wr��Pv�6 �w%ok9�xD^k��:<��t��<t2E6D �N�c*�ø�X�@�X�E(R���)��N�9���`��{\�Y�Q�J]z*���\ia�;����Եݤ֘rh�
B���'�j�O�&zl��5����wӫ4
�%$;� ���5O�H	c03c�h^�BD�%I%�>�\C�$R	es�?�8f�V��vӉ�������}\�ex�k`�)�	�k�t��aBb���Z�y���C�M�0���_X?=��MՖ�8\:2CWf88~,�_�%�o.y�I�����^v�=�AD���lА����Ǌ����G�Z��m�˩Tī8�>�ޤ��W� V�B�!�+��.md-͐�.Uj�,���|��;Ć(In�������}S���k�̞xu`�V�-���Y�ؠv۪H�	v�x�
���*��Ф�Ʊ<�>�j��66Nr��y�ՀG�^��特3����ύhy-��7w�}z�4� L$��d5'uW�8�@���p�ԕ�N��+�]{�w/�����Y��o�`�x���7%�q�qHM�
@Q�I����[M�'��"uٺ�͂�y����fstr��v��W�ԯ1���kt1
xE��ɿ��s�rp��$�<.J�6�i��ފP�)Ӻ��e|ޕͿ�~ymլ��P�Ի��*dY�oߊ��9��Bo��U�e�q�ŧ�.t�^�9�9A'���o=>2rBP�Ё������2�����)uM�x7�*�ag�Yv9����
����M�+��H��bө
g��z��!��Q��B��"Od��pjA�
��ǃ#�%�qI���F�F��r;�����/�����,�p4� �C�Ӧ��v��-l:���M�fjcB�Ɏ�3�P)^ӈ������Y(���K�æ
�Q�j�!� ���2���7�p�h�(�%&��9�VFكmOX���#)A-)�,b��D)=a�}����Hw�9B��#��>�$k���$�����J���0��+1���Y��EH��u7�u=W��[WS���)&h.�3�lpZ�� �X�3�✰Gyyzqm���`k`,���k<*�>�I���>(O�v�OI���lR�u �'O�Eҋ2Zw~��d�=��/�V�S���<٪�U	������L��;�ۉP\��%q�ٙ��y ���?�d	��<�E���r�eޢ���Z��8c
�/�t�����[ߦ��	�THܹ6E��p���ZP�د<P8+�޻N�� ���v�5Zz�<����M_��*��8�?�4��r���Y�ݵ"	6��y��>����Rt�լ~���t���d9K�
O{�~���Y�Q��:����7���/��"z��B:f��,�w2tW[����TV�lV��[i\l@w�_W��2��r� �h(�p���Җ!XX^l��V�ֵ쯡	�Ÿ�,�*��!M}T\%�Aj�;��%�j��b&4��l�
GGq�+@��E��=�L�����F[����C�y	�0��������TR5N띐��M��L������ʽ�@(�7�d�T���u0h�]���g���n�Rvwd��%+��FQ��V�kn�I�d�nm/�͸�<A�{Gr	0%��*�r����Ʈ0���U�n�z�VaY�F�<��O0�o��I*� v��{#f�c)�p	��� }|/�1���O��{����6=C�Q�o�:���F&|縰�>���Q�%f�*����F�hFc)�.�%t �Yb,�l�`��Y)�uۆ�(����S����dvm��K"�#��z`s/���2i9B�� ��J���&D�xS���̥�z�3�sYXp􋸔ׅ�D�]��9������f`k-�	K���X��u��A�����`$!��?u�6��>h&�����+݊~��_�����j2o�Z�Gd�I���s���O�9(���Ҟ��:زf=&yYr憁8���\��|Te}��'��Q�}t��>�ĕ�,��p��[��M��!Ր�#��j��o��`�e1�wdG�τ���[��b,>t����jZ��V��c7`K�q谈�[9��vBo�~�=m1q��h��ӹ�j���d���&+�  9Z�n��_�]�c^�_Ǥ�Nn#�\�����ǜyR�{�q!�N���K����A�E���'w�0_:n��߬Ji�F�Y�/��ڏ� ��O���{�1 r�05��_�� n�\9.�SR�lRf��˶�#��N�P;,0Z���W��.��q�Xr��&���2��u�7F�Ԝ�(��6vm�E�Dl�(1р0P��&�ʮє�aK=@�M� ��hR�-�W�S(�ve�%�H�M��4n~n*<�Cz=�P�]ΛO�b\�ڮ�J+�d�7�zW���@i�5"�Ya�H �k�p/WF��l/�x��N���BF���R�p�[��0��K��;�n����-g:Č���|�ˬ]o��Х�@�������UU���)������ I}��~�	-��%�7x�`r�LNl5R30��W�w�M-;[���>�7�L��8TĐ��56,/Ut�X�ܥtF����	�atdQ��V�k��ͪ�p����J#�蜹��8wtY�|!��Z<ɥ�-Yme������*�g�X
	�Ɖ�M���]�[0o�ϋD~E�'cpaƣH���K�<��]Fh/�,)�K݂�� ؠ����z���"�f��w�t�&�Y�p$���\�q��_�I���.����R��Lz� �m]&�L�μȯy�K��`�e4�љ�����TFr�ý�����C�1����6�V��%x�.��$�'[�WV4MOd�Ƶl�l�α�rSRt��ë�����|�P	��~V�����i�7S�V!��V;0��5a!�q|�b'>��N��1��ڭD�
���ܱ X��"�sO`�O?���R<W�O�x"������m�_|�Kkf���\t����8qyo�8��d�*�~X\X���0��bX?��-��R;!��]=��-W��gāP���6�c�`z�Tq�*	(9�����K�`*4W��U*=S��n��p�.����Ci�\�͂\B,�('!M���<t5c�v H���q���~`:�o� �d+ ݶ��@\%0*����W��{��49�<d�����R23��7�u[�J|��)i�*�����#x;z@.���`��3��J�e�@�B���7�~v5��1��PB�߻�`�1��vvi��Z"{P�/}��C��B9F�����x�o�����7���Y�yMjFŚ���J�x�fN���_�#��R;X��Bc`x�C�|]�N�T )?Kɬ�XF���ҲXP�5��#�QU�Z�8�W�]$9t!jlEƂ��:c��E"��~����o�� ����Q�|�=*׶�$Xs��z�[��|�(��M�n���6kEj��1V]�������[��`{�M����$�:���$��2�6��4�VD;[��7��4����>��+����v�ᩑ3��J��+L�Γ����{z�.��dx9E�N��<֙&��O߄�圝!�5����Om�_��I�ʯ�tc鉼�A��k)k�����Ç����(�e6�Vdl�Pj��?\���4i�A܄�꫞���|"=h�g�3�V5H>