��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�Nn.��kg�g�"�
������I�f�T3@�ͼ���x�6]����)Id��U����n>I0O�����[ _	�E l�Һ����6�+�'C��/���ڻئY��y�@�qF���kd_WM�X��z.�s�'��o���hg%��j@��2e����L�1��l�`�����nv8/�``^Cr�T�����ў1���%�-��|Ū�E]���ag�l��	�8�j��v����x�&�}���@Ȍ��U�I�Q��<����4�J.��*����0���f�HT�K{5AmZ�#1�w>���X�}xo����9 �rt��:�3������A���-�s?Y��R�?H����&��!��_|��]Ĝ\����@N��ɳQm��^y��n�.������A�`����5 ����K�Ą��vI��Ua�k�[ݠY�pVQ��+:!ҷU"��N��8g	�儬�w����?x^�)��B[o��)��V�6C^W%3\;3�,���433�(��1.�_Eϯ�!�����5�<����`fF�,O �*_f5(6����$��F���E<�����v�����>D�2�Z�����4\�=O�E�rT�R$� ���S3��h[k/T���Ȇp�`�K u��衹�k9�h*���`�LLQ��n��I�����<�ڱGVP����@�̋{��x���7G$�����ZrqT�_%j�|	}ܟTȊ����#+g�� �>��ވ�J�;~�|d>~^�mX�0%k�\<
`�kI�:��E_4� �L�h��ӓc��D��ASf��+��/���B��g�
T���Iw�x>���}E��Li@-l
S��Ώ닾��G.���{�J�$��S6q��Q|�_Er�G�E3�9/�B�.V�)��揋�V��ܭ�=�5$gy��k�`���w�������A-���ԣ���.\�k���m?���N��׏ �%��)<�B����t?|�'�Q��HEl{GAױY`����X���v�g���u��
�����80��N�A�!���X��3쿠�GR�����~p/@GЕyl��P�"ك�f|��c�"�!�Lqm���Mm�&��$Ð����R�	>:�0c�OFҴh>��q_���$�Zc$o)R�xYg�(`�dRc���U��RȆ�v����6qR�x_4^'�aj��|q�����n�w�s��yw����UB�cEo��<�*��/��naT{�'�.p�ý?aqJD�Q-�_��D8��Ӓꞈ��X���}���|�^��:z.^w�ٜ��M>T��ة�X'��gl쌡`�����I��|�@ �;�uU}m8xW~7�����S#����4j��5ja����0�� ��u3��j�r?��Q_s&��#��Nn�"C�p��m��9���c	�w��D۶�'��j�6�@h��c��窠`��S̡۷��[���s�[݌����_�ϑ����n��"�8������6���W�S�8�;7��O��N�tRWxp����v+T���@X8ۇd��r�fan̢�ߥ����\<~rW2n}z;�-�n���D܏�X��]�j�����N���f��U�c����tɱ�u	�Vo��� {����*���[�*��7�O]���j��yll7F2��R'k�
�Qd;�����醮0���y!�ll��}Ϧ���7I*z��MI�9��z;
@���b�Z������4��s����@�L�}��
�W�Q�=z�-�έ�����Z�����;��x	��i�)���%�B�K�:��QA8��
�Wr�~C!)�g硬o�ΡF������s����hŉ�֫Az���O�J��cBr���aC���5KB�9T��$^��r��KKK;iM�p���n�^�ԅ��
 %�^��,�@*@͈�r�Yj*��@�&�|R+�#�5D�^�:z�b	ߨ�O�8�%5�l�wҗ��s�ɳ ���H�х�`����4����`gk�p�O�_��_�wV���e� -���MqС[$�m�̀%H䲦�rh�t�
���!��+��Z�s��Y�)w.�n�
�#� �S(��BD�(y]�>��?��#Qޜ;,��k��ݮ?C����0�|9�!����v�n�� �40��ϫ�\/!��l���
�R7�[w"c��s�V�8.���!��]�h�O�/O~����z�2�ů������S����4���XS�����c���P���}@���6�z8�6#����}�"�\�Wj��K�2�^�3g^u�p�-�Zh%2�9ɥ0�$�Sit�p�M�D/qp8}�#��כ��J�q�;Hd\`A���.fa�$F���8��Ğ$����N��b�P&c-%A��+���J��6@�Ҭ;G�)X���� �+���nAߵ��݆f�(~�U��?��;��9�Jl'��Dk�
����� C�k _�ۇC��Ts�ƃ���X��)5B�TtCn��X~i�P<ҁ9ܶ⓻RW��e��B�C�K�o�%�Q�#��=�7��E9�Bvw1���"�fv#ggypd���23�{���Y-�O�m�d[��!�KE��代Ť�l2�N�	�u�}	A�+���9�n�0<��hW��ڊ�����:{�%�32�<s�Q7�j����y�U�dkή��*i��"�A�4�W���}��S�������8y&`XK�����|��n�XY_�����+n��:-μ����!�֣����6��I���*�YBv(�tx���⋏0%P�YUٖ�p��Y(<V�����{>�&�r��)���~�ף�ۙ�2$a��%�k	��܊c1D�G�⥷�� �=F2��)+�Y"��+��L�Kqi�X���▘�W���9��|���u��{-s%V�g��Or]�l�#��9a�����8.�ZL��s�Sd@�����&KVBv�2_��	<nm)��#ف?{�nWX:�x�/�..d����
�} �Q�fʣ�[�<�.n�䰠(���{�2�d��ϒG	��]�E�� �a�k�V�uT�N�l���|�5��N�~g�Ȋ�ɣ�!�Mqv�z��0!�'�s2�8��Pq�(�q�B���Uce��/T9��g��~��Gl>��S��/:�&[���p?�t��+v���Q=[��ˬ7S��GU�Q�D�;Oc�<_�.�#D���LV��݈�'�y]tpY�F�J�0v�\�'�,�J�rvLe��%�&��k��$����a/��>AF�̈́��I6�>�x���~߻3 n3����Ct�'<ϙ�E0Y�c��	�����LH��>�q��L0j���Fo��K�s�)V�����s�\�~�ʈ3p��{��o���*�sXlF�8���!?lH�|�F?S��������&��VޝI�\$�4	�fCk8�__|o����ٝ����g�.�f�=|��Ɂu��KO�D�C��d�/@T[�=P&�ܯB�2�3w�9A���,r�4g��hc��~�ˣ%},:C������-vPZ7�+R9J!��p��^�3����N��9��k�m�5��<�.Bi�"z��B�[�}�d�D��]� V��-2��z<ύu�}D�E��	���Ee��x��Ԯ���&���ɵ�ʂ�*�5�� ����r+����UqإR2k�v��y;���&��+j9�U����;�2s��Cg���E�-�M�n2��B���}��~��}z���mi
��gi�L�fo���.,I���
�j�����::�1w�jV%�r��������D�7���T~��_Q�[0�IBcuH��{�F�\B�~xoP�;�u)�1�|���2����jng\�:�m�|��H\[
���ō1� ��΀�>�{�Ý,���@�A�4c�[/�0�X��J�.����q%ӊ���P�+d{O����<al�[�N��ܿ. ����a��s�M��u�M7;��_w� #�+�����7n�"58R�mu]���`ݳ�_�$��������8��~Y�Ӑ} ?hn;�%$VsO�փ`����w`�r���\� v�Ѯ�*�ؼ��@\K�v���ƪ@��n쩩���p����p��jΊ����#�7S�o�	2�������1�&������?/а�� �*gղ!���P� `�᧗��G�Y�|�;J��v^�>��;�e%�\Q����Q�J�[�{��n^+�]�jP��� �H���������\��h\� X��������so{��P�n��q���*���c�U�g�¬�[H .�3�ݝ'
���W�raW���\�%$�6���K�)��䪻s���e�kF����]�-$��-7�U���_���u��Q����i7���06B�=i�?��ø�NݔŲ��)E�\g%�)��NŲfJ��v�VӅ�[m�3R���g�m���O������lF���v
ޙ RL���d���1��3>D[hŏ��T��������E������o�� ��y@��%����'���x&��m�s��M�,�C��d D�@����D[�O녠%c�����.��� ��%���\~]�l�cwF<�X�E��v�>��iİn��5����zZӷ.��_0��X��%S�_eSK�7ԟBUP���uv��?D�k&�-Uf�Dw*�����6ۀh����k?�ÃUN�qǬJ+py3x�/��4�hE�z��_�@*b��:Sqږ�'�~g�;��s#%��y���,�Ɣ�����l�(\����|Z��VV�%A�KB�ܠ�
.t%eZi��P@���Qn�*�F\�U���`�W��s�s9��Q��`L#����,O��d���$nB��� K*�&��e8�TT���KE�k��`�#������l?�ꋲA�������N�; 8z��)�!�稬�i��ǩ����_d��WR���J>	��h��z0O�
������k����NJ�O�S���t��#t�DI�,��S��j@�0ouӐ�����{�����y)S{u���u�ҋ��;Y�������S1?{��pkw��߬��'s6�9����`;�*�/H
e	�.�
��c]�X~�Y�{��x��ґQ��y�r��I���!\sW/n�D��|-c�( �T���p�Ox|L�<{�� O ��l��g���F�{��+��n�������b8�V�d�j�'k%���Un���h��Ǫ��}��$��h�}���-.�>����v�l�4�_~�X�Ɛy4Y�%���vV���<=�r�Ral0�t�Ëއ�CB�V�%Y���0��x���cG�- 	�(��� ��`�V�l�_�T��2�;Q�(Ҏ��-�鉳!�#��t�J�:	�U�\�O�.s�5�9��{�`ln�&ӋLy���l��x.�p&�)̧����d(�}��3lé�Xf�/����h�7�H23����r���*?����z1�k����MPt�-\f��D��0S͠����ym^����:��a����(�� "�soI����$������\'���W/��1U�����|�T��.�]���B��h�^�\���E�P^��C�XN}������>�����A���˄~V ֵ��8.?��(I~O�`�>D�)�F'_��z n^������y�9`��[�Lx��b�8�,������u�@�	E{d���y����7���i��[
f?瓰��K���Z=�s����2G�ɉ^uv��h��_�
�N���DzU"	_V�T1W�C����w���f"����5�B%x�8�(��Q�BE*ʧ���w�<?PS����Vq��9$EBL�2�)I�>��I��7�O_�����OޏĹ��='���XNP/y6��Q��PEak��f�ɼ����c'�Z��������X�BB{jI7DK#!�f6�{��8��~N�`��~��缷�2��n �rٜK��EWb��O�Z$k���&�`++?�x���Ɛ���^����Q֭$�}"��K)�)H6����/���ٶ���<�bK�U=�U��{�2�/��E����w���9f�1�t�Ǹa���T�ԫ�{{.|2	_�1�N[y<ARzm��5�=Qo�V �+�te$�%�@�����4v����	�$.������*Tg�Av�I�U��.Q���ܕ���-)�YɄ�G���s0|_�5��4����%��fy*K4k�Lq���JW��N��l�:;�����͚� !�!\��|��D�M�ڲW�Mqe4����f���d����`��s��>3e���;���l�a�x5n���V�������B�8��ɺƈ8�H��PQG��Q���_�r�m?Y��̼Kp�}V�)�)eg�w({�@���P���@׉���wYS�K��æā�;ư����0��!�f֊��&o߮q��>:�"<��D`���b.�%��Xl��\���n3��_���%5&u��Q��8� �;�Ѱ�)	Po"ܺL�Z4��˛�����2�EO8�a0[[y���|T}y����c�0�9�EB�8��l:�]���=���\�nm���R�O�� � z��w<V �����{Y�HH�R�c!��P
?�tDQ�������O?��N�3��^u�&�]�¾"c���J�u�Ϳ��/�i{�inV�p����`�\��
�C�P�j�a�ˎ��ij���`�}�8,�W�P|��QI�l}$뵔�-��U��(rz,�p?506/�c�#w~D��������-_s�VY��D�=[�H+ׅ�	3�n��ϛ����([&2�윌.���l�A�g�v��D�d���������Y�fw�;�22�x/��5�Q���.�T[h,E�L��Xy1կ��9g��mZ?�Q\1ӏ!�����O� ��������u�4ʽ�,�E�S&,NhP_�G�/NI}2>�A�E�A�rZ���F�Ps�)�充�.��EN��G�����d�3���J#�䡺 `�@u.���;;���¢I���i2��]eB���$�Q�Pנ��m�O,;��u���S�%=o�QQކ�;�����I�d0�����b|<�~Pm������tu���?(єr�K�#���ި��6<��ǽ�'���?�hx��n k�h�F�ی*�D��",ym-0K�*�nQ;��iv��N8��A��q���`�0���}s�@����ۋیٵ���Ԛ�9����u068cPt��5b��L���"}p-n�8s^��Hx�R�;_�d0PltU�.�([�#-������ծ��5+T��i��Ħ�`2UQ��u+���N���w��-w��ya$̆�w xU�D��kc���k�����[�a�X��3ݨ�� !!<�%뵨[�R���nb\F<��R��sӠ?v���G������	��H@�3=�f�Bz6�� ;8ƃ}�  ���ZNꎺ�x�~[rU���V����U�E�C�|`�!��ґ�N"rI����]�0K쉂�6����K��s��EF��*���5;JԞ�\열��)���6��e8=�]��A�a�~ՠޛ}�B��e�eJu�ȹDn6&�G�U1����IL������e��S�0k�b�?#��4j����k�~${}��y`���}��!}{0j��<)����G{�DS�aL�i�:jQ���)��:&��)Zپo��x�r��bKv��'�g�$��~����/���c���/Mf�Nغ��z����s�F�n�'c��=�aFM�K�PWHqӫ����^©�Z~6v<�/�y���A{�z;��E��˥���������-�T	�Z�u�G�Ӎ�ŋ�7(NiyS6\<xn�-"��E��(hؗ�j]��ᙙH�k��$:�7
T�.vw�Ԇ�RĤ�1^���f�$�����PK�Ҏf"�x�j��籯Ma`���pIhH��Й>Ȑ�#�ȅsVw䱼cܚZj#n�ѰL��dɶ�B��+�c�ciL"{����q7�[}!���aD��$�I�u��
��`[�{�K�C��9�۷F�����蠑���y�n�=���;�:�l--�~��$6�U�:j�}�ɿ�%�u?�9ٲshc���#�-��OV�>����)���9���n��v��B0�m��{J�UJ�m\��w�W;�� ���]����W��;�P�scvYA.NG<-��>Iͻ������xW�1��>�5o�����>OU�1+���P��_�����ε�����zq���8�w���MBED��!"�Ē̍�.x�cX�ߩD��z�0"��W����{�[W6���,O4mM4
�nZm�����)���&��k����3�xQ�t�;�&�l���E�B`�O_?cJ��s�	���?��c�'��*#g���xN�^`�s�w����IW���*J�̩���@�"ʮ��b2`�9O�o.��(5��$���O�����������zִ�� ,�($,.��z�P��9N��rH�I�Tq�0���A�~u����jֻBn&`uͅ�����IWH���`����1��$]����"F��D˔�~����@�UDi���[Fz	�
�b�,	<!�ߏ4��g:��tl����X�P?C�"K�o��V_�2�PEaն��X�J��AH��EKY���`\�@;m���މ��].ΜROT��xK�2�Ԓ)��5�ss�O��������\tM@S���k4(蛖����'��Z�
GS� -*,^��ĺж���;|^�}D�u�0LL����jE�K`���b��U�U��~G�9d�ЮW�+��مO�F8\����	���1�5脲�� �/��q�'�t<��Wf�=�D��0��6�"���^��3��v7{o
_�1u�#�{�U,p�DS2(aަ�"Bτ
�^h =����@WU���#��