��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHnRN�h�\��%�P'^�|K�G�ݡ	��b���p@���=���ծ��t�f��s��%r�$�409��,���ɗ���35Ct�c�Vp��	)�>h
g�x��+{�/��B(�VQOpO�7���Fp�h�~�F/��f�	�	w�]�4 �y�F�ӊ��0pv��T=��p�aL�ٽZ=LX0���Nu7� ir�/��< ���UqR�n���B����\G���{f_���>�H�O"��Hb�����aܥ!s��F�S���qL�<[^��n�ȏ�>�
=h'����ϑ�p8�xo]dl7����Mt|U�#��K;F_�AD��qK��$(���B���k��}�b��m��L����>��6���Hh�x�@@�ge�3�>�/��>	�7/�vjr�f�h�m�맆ax\�	�K"�t��}眶'BI�������b��\%
;p�!M ���ln��:��(}�p������G���������E{���r�)a� ͐�)�Db3 ��MFfq�,D��T
�_l�36:0����9E�90���7(��rj-���L2oD�މ��� /aZ�GH��<�-��Ȇ0,��t�/NH��jV緡Qq��s"�4�vhM
���Hʭ0}=q�M������%B�K*����cY���~#M��$qҔf�6Kp�XՕ;vw��~��pp�����Fu�e�a�
��$�о#ɀ�#[J0q3������fw�lI�2���P����4���x��%jEX|�R�L��U���H���H�|�J��4�퇵��t!�t�rV6�����`��Ƙ�2�Gy�X�hJF��-1r��o��0m7Hq����"�
�f�.�>��-�B���f��y��j�E����52Eo�@��v�-'�����[fl��zg\a�G�$0j�X����߲��%�������V]�8!����,.:�x]9�a��U�׺�׸w-�
*%�i`n���]�al�h��̸���!�(�tS���7�0��;���4%Y��l��!���%3d쾕y�ڄ1�s�*\G���.c�Ǆ.@��/���(����ђ��g�>r�\��J�(�(n��r�fF7s�nu���J��%jrc_!)�;P�x��������󈎴��*[�`I���?�BU�[�K��e��:E�K�Ͱ���pf���b�5Z��h�C��7W�6[%�$0����)Z���F��m� v����߬�#Ĩ��{۹�!~+�*S�<����)tp�%/�#�:��!n�M�*3]�8Ui�z���c�ކ��(��Q��N!�):=�����B|1���}a+��"HJ~j�wG�M�J_;$(���n�	��"�{��m^�
$Ճ�ǜ5�۶�S0<�Q�9�$���[E���
�"��񍈛'�̈́e){�mTѮG�
��N������*
Bք��!�S�Lm���wi2�z�MR]m�cX��}n���K��*���J���a;�����AX٢Ou<��/��	�3��$�Iף����,K�x�y~*�E,}��|����=*@�}[Gu�7��jJB
Xb�>p�ߠC�oۈ�Ơ�v����;uB���)��}���0��7c�0t+Wӿ!�Pj�s�m� 9��5a������l��<�3du�.m��Fr�d)(�����r鴗7��}N��!����{d�?�Z�M��j@�;�i�����yw$�%�zcr�����3��2l
c4>��0�Jv{j�	���Y��b�$Փ��?G���+Ү�3�H��P���nf��.�Ɲ��D��QՏi��}n}Z#�n�,����?f���,_��Ω~͊�oJM��/��E:�̒q,� ��V�h�.6m�+'#F��1��L����
���4��W�1��*'����g����	�T�L����~�,�҄�R|]e:)�ߴ4�izSu����1�|�#��F+��+�0�g�Jy{o$h�H����f�^�����i�䗍�¹���K����x��ܝV�)����L+�Țs'c���;A�]�H�j��H0���%	�oh
�\��sXFH��#b:E]5�j�Wڑk��Q��HQ��u:��8�P�VQ[cz*=l=iIW�#���(�R�e\����ݝ4U���n�aB0��4��Mj�{�_;�L/P)����Xn�ϛ��G_�]2�
F�%��1z�o9"a_+�4�q@.�<��=1��Z	�Є\��y���������f�������&J�zO�!*r_�R�.k>�1ǚ�����#(�LS��^�S�ȕ��X3�AH�B����:��a�#۲�[��P��]�WLbs��vV� ��Ip���^7�`����= �v������-�d}?���	d��Q�rĭY���L�U�,�YSfw��Z}R�dŵ��zbJ������&·%�Ռ�S%���ě���u�Z��ێl7�=�H@x*�ں�P#��Hi^y��'l����h��eɿ{��'���D�>�����ܸ�@���}3��i2-/�87���]W��|�޶���Ĭ�&������}}�7�s�@ocy�1/b�4���&&����E�J���MJ�j\���
�xV�m��w6Ѹs]��@�C��	c��\Uȉ�}!�z��1M��=	ޯ�IM��诎+��Q]� ˹#���(��:w�{3��4"&F��_���H>S���4>�c��/8�>`�{>�=f�jO�&����S�9R�hasb�C��H��;7���C�#�{�e{|�e���0t�G֎�V�,}/ʩ���@<L=�������TG���{��2B[4\vt��~0t�n]�t�Xi���o:"V�\����
5��~5�{W�����E�\I��y+��䴝H�*2�؋��+���ShOgI���<V�)�p9���C���-�B�٥ź��?�{q	�)]<�G������(�?�u[�)�,�Jc����솁�^�L^I������F&�M�ڽ�����	o�K�f;�dS����������,�������
�0�8Gᇣ� �M��Mo��]�n��Բ+	���]�[�.��,�Z���J3UF��3���L�z(Z�[��	��B6��=�E�"H<ގͅB ))�f��ޙ$u������9/��(�4�Et�)�y�,��i:� �(��DE�J�ԋk4iu U�F�f=�\[��e
��k�a�>bs��D܋״S\Qy���+����a��]��R��~�h����03ЍS�a�wJ� L��H_��|�E
�C,&�فv�>g u�]�L�����L]nL����d����:�x���;hOQ�'�|���(Yf���4���+�?�gv��>�x�ǣ;f}���<I{5#��*�*8�R����8���"`��P����`c$�.H)N�-؏@C�(M'�0��������v�aY�rU��b �Ԑw;w���%����v��8�$�1���e������5tb�[��>�om+!U�W��`�����:jL�mA��Z�ӻ���=��c�1OTؚ�E=���o��k�TYi�֜	�n��<�G`�I6��Y����:�Q'b&9x�f2Q�T��v�����g�@]O�������:U���G�Q�Vb��(��D<��7��sN5Q���cg���&䢨$��T'*Ѹ��c��Q6~��:��P��A����IF�@�l��g ��[Or>'��2d	�Ban�,��v�f�"����v��Ak3S �2/l-��$�¹�u�JV �
�ŖM��'U�2�~�x PY�V�df"h8¶A��.�m����|P�����S�pL2i��#%W�[HPG�%h�8�������E:�Q5㵧�8ˎ����w�DQd(�Q���	���%��7L��4�S1�����1���m�_�eT0���d�i�a���pZ��3��"B��W�%&��x��I�֐�t-�_��s�k'�����a�/�p\ϲ��"��9��{��+k���������P���\�>�hJs�pN�5yr�����.f�e�@�����!<��&(�c��_ݟ��k���F����amIE~ �U�fX��B��Q-彅�l�w|4�����ӝI\F�	�jDπ�STU���%�`! }��`Y&<�\�e�]m���}�^�w�1#��<�y��gaoSԯ�r:{���gVj�iH�|Y��K��Lc����uJu��o�2�c	��N�E��Z��)RP3���
�J��,:�F;�I��r1/\+���h�IӨDr[%�-�$�	�=烾�x7��k�+b�C�}���j��U�!Y"�7�X����Q�@m-�z6�a�e�N����fc���/�ݙnM��F��w��y[�}�RnN�ĬT���2�p���m ܟ���ؚ�ҙ'I�{�c���yhؐ��o�Knp�->�T5~�@���jKͼ�c =>��~�����-��F�0&֋�큎�a���5�h��u�T4�b����u��֓@��BU��%�:Ei�n�8�ܖʟ0��D��S�^���TpΌ`�n���m2�x�R=�|`}^�jI�����>��'��R�f?�p���չ�W��m��� F�*jd��O��6ԕ�C]k�f=k9%�����8��(�$��N&�A�Z%ڇ�t�g)�\�(3��/(s9��s$�3��	���	�R*z	���(=�_��Ar���; �m�c��&�>�O��XX��yM m�toOoq�)��48W���8�PT�~����%�8Z���FpT���Sֆ΀�0a5����f��Dg[�����KF��!��z�VG����F{���3Q��
S�MږE҂Ȇ�Ȁ��#��e��|��G�]m�pw3���ã��o��;0�Nە��i�������j4a��\�p����9��i�:�k������e��"{a����m`�U,���D�&�����E���o�Ro�I��N�$������@f�u i�T��۬%�%b�NAo�"R(b��M��o0kN[�b�������'y��B�)������#� Fɣ�Z�g�Q>���ݱ�
9�|�d,@�CQ��ve�����Α�8ׅ5�Kڈ9/&��E�R�"9JK,�F��ā�����#��*�(��q^l$���K�l~�Q�y�����8�P�8tr�I���0���{T��<��Tck{6�G�w�c��*��'�%�4��]�'�`R:<�Z����GV�������*K��v� �^�E��a�%��P;��ۉ!�F���ڞ	�h��5D�gY6�����\M�3�~2���JIhf��"�'�&��7�M��{���	\U��\��$:���l؋���w�ո��.��&�h�g]�٨�.����'��)����X^��-�na ��nR�!�1�S���P�Í�JrA�\�<�?�2"���1��X�À�%d�%�k��2�D�<�=B
�h�y�(�0��ߛ_�6�J�1�(4�F�;ymy�O���b�&���*4��<ܶӕ=9�K$#Ǒw#��w����|�}t��{�4���NU�4[�=�:�H�S7�E~��_T,pT1=�oC�b���7�]c��VS7�I���vm���W�L A4�P1�c��Yi�Z���*�"��2Ѯ6�� �@��j9zwj�<b�]��v��11ͶY���9��`T��NC=a�x`����
B�\!f���6Z��s�(��Pw��F�}ב3J����L���j��1����l���R�-��$��B�)�|ɼ��5����l7��ھ�s!ʭD��Q�QZ�b?[y�|����(�A��q�@��� �3���	��],���>�َ8����hP����e�+�JLa�C�]�i����5�n�q� F���p���� ;���4:�Mg����{�$��a���Pԯ��jM��;O\�!�*`;���*[gcM�w3p�H�����xl^Ԁ���8�4�H����z�fJ�_Y��t��;��BA��o{�\�UnL���m��!L��m��w�����V���a9�?�-0;pnhN[�&Ga�w��Y�z-�����Mi�#�a����Jz8�I�X��)�p���\���j�H���8f�{Qc���=,?mb� �M�[�f��G�B+��9�:�ʼN�1A�&��E3��"�-��"��X+���X��$��c��YhTY7=�M��*M��"�t�(7��K��p�FyZ=&�1N����>�NʅB�[r����]�W\��"��ぜwb��&Ӷ�C'�W��l).�o�J%W«�#3·2~$��ם����r��/b��L�~Z��>LC��qu�����L]��8���8�Dw��	��c��Vs�.-��Wy��Z�wN��o���N�I�;&���n��z���5<����EH?�Z�U�G�g'8>����3��G���mAs�\*��X�r�l��͙����ݴK��6��W]aV�;���X�oVeǉ��� �cR'��}�b���܂&�o^��_���(�GZ�/��E������cn��G.�oƯ����n�'����Ug���>��)��T�0�'�3z\�7��w%�T�� ��z��,�8�b�e�Բ?�'�l"O�N���zⲐw20$�x �`��
���&����ĻՓ}ϴ1ϧ���(X&C�ܜU�/���-Im�I(8��q#�4 ���������Xv�N*ۋ�������X�ꚓe�㚋,����̉��:
Y>��_�2�Y��!�o'S�x!���/�Z�4���g?� �908č(��X!1�n:��(�q�[�VW���W���Bc@`i��[MA1��`G��_{�u�Θ��7��A�ޗl~S%���$:�f�e��Q���#fw�H'�Εe���� <KT��>z�� �Qʢ03����7��}y9��*�ؠ��߮K��^�����Z���*��ࡳ19(��+�B�~\r�Ұ�^A�n"����tTw�P�[h&��l�I<3f��*H8�=8C�ׯ�������3�Y`��E�d!�'��;8���n�߇��k6��kkj<U�Z�Я`K-��\����Cg���ܝƝ	�$���S��&�B8���"���͜8d��)f�)�F��k��V��4��0D���0�'�3Vc
wǦiϚ�9��H�܍�g�zC�yRD���������i��I��ˢ��[��d�Ӗ�Ѭ"�.���;�8���h��s��V,��L���9H᮴,��|��Z�2���XD��-��+�|�����ʰF���^W�@��ɑ�ZXf�+{�_:�L��q���=�U{R�Q�|��[$��D4"��mw�� �&|=�%�,Z��u³��=��oܢ�.��j�L�Xt��%��ԼGY�~3�5�Ϥ�t��	��K���0������1���b�Ɛ�n�1o�1Z&\& o���$�yۏ�Ax�z)�2��d�F$�:?�s������>���hy{�S'�S�xyt?�&�	���D�s�9�P>|��?{9�ϐ#��o��k_([�12O<���+���H��-�&�l#U��ӿ����[re��w��Qd��	�/b�ꦢ�++��w�ƿ񁩡�y�E�����fW��:Rt�F�a=!B�Q�.Hvˆ��H�m�R�9��& �f����b��	�d_מ;��U.u�%l��p �3y���^=�j�$'���l����no)��C"�:�\�~~��<=S��3�˨����N�X↑�=/_��l�z�|ف��K]��R�re0�	\\z���VFBb�߰�CH��IpΌ�3w�ۿ�[;�}m/�Ԝk� ��sjW��H�z��_l=+'�"A�{I�����&�{<�yb�� ;�c3p���E%�\�b�[���:ɐ�#�_�MU�@��y<Y�chOr������O)�1�*�X%���Pv#5d��A�"�Jݗ����ij��h�����7��<#�/�<|xU-\�m&P�M�2���Uscx a [��A�yj���J��~p�h�=VNq�眔r�m�mA%�CcV<�({
ty�ɶk�F'����s�K�΁�v�1�R{��xO��!͸&��N�ږ�9�n��J�;��Ed�4�߻��?/��lĬQ��-v:eWBw�Mh��}Būcf�8�����-=jB:����@�Р{ 8�J�i���O�����������q�+�������3���B�ng:�V�z9�p����:�Ƒ]6�fD�~9`��Ũ�\�evi������|�ֻT^��7����g��"���F�~m���;W����!�՗��fO�ffXS1gMʷW���o(��ۈA^)oX7n"O�|����
���ʗxޔ�/0h�N��.;�$��@�$�f21O�3�XYd�%��XŪ3�j=��ms:/B4�<-��1i�a@$��������d��H���
�E�pmNށ�,륐�����.�
:j$�*���Zu.��5���
���d��;��85e!�(v#��A��->�:P�F	f���[�\��z�g��.�:�cg���z���TI�v����6�(rSD�#!�`Zd��*��[֊
$�����S\kd���r�t�Zm�Yr	?�����VGl���0;����3��ѿ�EH� ɄC��N�l�ѥx�S��WN���@��K��Ciu�=sW��h����mF�<ȸ�Ƈ���L�R,�Ze@�`5|��2��Q��2Eء �^��	�D=�rs���V�JR���9�:&8+5~�N$
0K��00��]��d�̎t�X�1=]�mX�xn��u;����R	�7�]�XS�B�v~h�)�wJ��C��.�BO
��b"��p�P@<��Y4�����s`,T�!����7!�N }������-�����"��'��ʶvd��Y�9}JJ�M�H��
���ˊn�����v�R�/n��yk��
,.+���f��A���T�����)S(� <�Jhvj�$+��dZ�-�p=W�}�b���0[Xk5!��怟�c�N�ˑ+�P���	� ��Y�'��1��9�èF�$�@� �E�@R��vyV ��Э��2z��A�]a�D��,]������ҁ�����OI�z����[o�g�G�&��Ey�]�����W�V��cn��;�A|"�# >k�㑑���5Shȋ���:��K�3���.�I �;}��"ǳ��YK� �*}V-ʽ�ԍRֆX:�ԉ�ŷ����+������]L�ៅ0$(����92�r C�ϭ`j�ш���/���k�*���������^T�����`�?#��g��:%Y�`$Dr���,^|Ը��,X�}G9�v��-JQ��i٫myrūM� �yi�&um���|"NG���Vl!s��W���� ��HxJ�<f� ^ �_�d�5��������ݨ��N��ZZ
�F�{;�#�{�\�S��u�ok�S��Ȧ�JW�w�
��V���ϬI�Z�+2�Z�2��v?[[/�
1�ኯr���Q��}�e�����XH�ld/�-���¯Ф������:�pK��;c��f��ʱ��r%��b��ܷ�(��g����1��m��I�g�"������<t���{hs�%���L�]u
�=
(E��k��8mn͚㻛��8���?HHQ�X�`�3a�\Bxl�R�����+vD�v`�d��j.n��T�C�8\p&	�ª��6���M��Wt���3����mr� ����c�S*�t����m������i�C�Q���U��ȡ)=q�˯$���q���FY���^Mb�.�䁉���7c�� 闫)\n�'UwQlЈg���/���^����h۾�&�c)A�f_l Hd9�6���ac���Yf����A^É��ZhW�+�lN�N�2��,,���Y��SP��;�����NxФ)Ħj�t�k��~� �=��ᬫ��熽��;�Awy�Ô]m�/_��j��o�n���m�/8P؄�qKJ{���7-�oĝ5P���@����H��ん 	P��mX!m�ҭ�?讔�dp ����Z��qd�#~�&E��ng7�X
��hOlu��_�����~ew�>m��&1�k_�2�ĵo�f�"�n�Y&�ka�*�!�w��(�[\Kw'�Fy���xb&5��v���Q>�%�	.wK$~V߹�?Y�Y�@� �9R�����y}�Y7�׵J/k2<7=Y��}sd�n��T�v\giV�ërf�o�cé��.�	K������gz㶲\����=5��A݃R�=y�v��K�s�x��L�Q�y0����@�^�T6���77�Ϛ������'�7T4`�D���vh�3�œ�
��ϭ��n���HA����V}(��<����ȟ�R�N��}��d֡�A���a���:���U
y�#����� �V"��:X��o���*��w���ۺ�z�.<h�|y2�7�y���4�� ��<0P�֞NI&DXJkP�	��s������,��сْ&�e�ee�f�8A�:�v�3�������v��d?�b8�&��4����+z{�_�^��U@�o���NSd��f+�Wn�t�V��J�d�P)6�KbK���M	l��RvY��o���K���J����8�܅�5�#nb����ՃON�c�3�2�%Y�	��0Y�Wr�H��&�%�y{�6�ש�4���ȶI������VSsu�ouXz��h��7�,)��0� OdN;,G3y�ۦ�״櫒��>0_A�.ê�^Q�4������˃w+N���#s��;����~'0�����@ޣ��J�M`i#FSm� �]D����6���7 ^a	����a��&wg�`��K�G<�4�`�V��)�ۛ|�.��TɁW)<!g�Q��BӪ@{�9jJ�f���(���-W�<��{"�s��]�A������z���f<�z���<^S���%���e1bO����TøNRҭ�{gl�W�Wn�\��M�a(J#*XHhy�f%.��}(E���w]/Jt���%_�ڬ�.���-͢X8T�媬a�h~6�FesA�����jc3@�O����f�]����d��{{ٝp�S���6�ܡD���@���t�����Tz�)��u�&E�1t���/M�c������´��@�뛫��Tu���[��M�:?$"�f�����iA��BuO��M�G\�8/��-֥�-A�����^���!�L��p@�ӏR˼��ޙ�}�h��XC��ڑ"D`,�1��m�eޟ�k�y7)�#���Vhj�L��1'b�\�Dq��gu�\A���&F�w�ܤO��)ŏ�ҁ��:J9Bvf��.��PG#������%)5)Ƣ��[ڡ$�4��rr����%���y񌱜#Y��gᜯ��^ �K�0Ȼ��n��FTbfG��W?QCp<����;7�mJ\��Uܠ�%J������.�܊�� ��B�`����sq�xf�=E�3<\T6�P�Ø*�J�!n���e�h"_WD `��5�����v _;��|���LHd#71�8S8Ä�N�=�s9}5e ��gZa�f���T�Od��/�\�D��M����$�"
Dۡ��>��'h>�4����v�0SI���I6��[3�����-��2���qK�a�+L�Y�X
��4��>�8���
vN
����	�E��#�C �~�b�8������f�3ʹ�(^�9�<�����!ߑU�tH9�5��܎�3lEa�"���}T�q�5W����C��$���3W�i���K'8���og-wM�%�2Uamɢ���4����w�w�l��'��zv V�,w�	�L<�)�(6�<FE�-ce�h� 0�4����lQEa ��o�r�S���۵&2�[������43�l�n��50M
� �@L�Z?�ղx�z����Ht�ֈB1�)xטxn��x��L�����7���b�r��L��<�Q���$#�܊]���.�@Ui ��ލ`�t��)+�{�͂�U2�7���)d��2[y��p4��2��q�ڧ.�1B0�(JR�&=2	��k.���+
�P�#l�g,���3É����ؐ{�6�?f$�+*�4;���+e*�q�C�*���6����]���FL%ܰ�#6bͲ�y�ɔ�M$q3�J�=�͐��UW�
HV7�Z�2�$f��@�:k�ة���t7�q���g�o}RJG+O���Rب����S$�#� ��+$1�r�#PJ!z��+FZ8.da򵞄*��CJZ��bDǔ�f�r�o���X��	u#a�g��d�Ěg���=���K'�ǹ��W�����ݿ�7�a�K���D.H���Ly�g�{N )���X���G�1f���lYd��t��9�Z :�zt������ 4h�uI�י[i��JYV������O*��n�$�~\�� ?���/�!e���'Q赠ו��>q	�X��"�8�GI�0�wϑL>�]�P���)������SHx�t��a@�U�V���?@�Ȫ,�.BPd(Z z4��r�c�ek�T�M�� �>�zv��ߧ9e�Y8J\U,4r���W�]G^1�	�Ie�%*'�y��8��o0��G�1u��D�[ÉwЁϿҙI-��I�#����J�?-1��q�Ea��!��"x#�����I��|*�rk�5h8���f;���^9����Q?�g��}Q���~���CJ�p�:v��� ܖ�v#\X����䝻��l�(�BOx&�~���Q\'儚N'#'� ���u�s��<'����NF�Ä�Ҋ����5���3��Y7q�!�hؗ��¹�������G�rw�:�p��aeX�+�)*I��� Px�B���n�gD0��<`�@�*���`fHd#��7�6��N&������r�tӮ���i��m'D^���}�p��]+�i@�b��]��L9B`���Wc������V3s�a#(�C�e�[F	)
�H\C׆NW����C�k�ՉW��A�b|[�{��هI���5$d�ݢ�F�C0��J)�MV�	���`���* <D��s?b І�w��
�N�p�:�`�~1� �J6sD9��o=6�!�SΨg�
��F�B?�ƶ���(��I:��X8,��3��� ��5�v�1C>�!M����F������LzB3��������C6WT~��4 Q�ś4��J(���'��-�Ce��iv���V���,��( ��9���C�˳�3��\��l�n�=KM�t�����^H�T�W����/Rn�8j�pP%�f����t>&��{�ǑG�ʒMV�O��)��ׁ̈I�<5�}��M�v4��b��D��ʯ{�u��lUc����3�F0���I���|�]@��f��Vq$�0N��u��m�����|+e��O��H��;LD5�5�-8�Ƭ�*�2��OY���3����g��]]�4]G��4�8��MM�1|�7dO��5��W(7�E���4���C��w�oT��5mң��F���p����Uqp�^N��JJ�E�9a�}|*��L�l�m}x�Sބk���e�f����F��	hB�X�f��"'�:v��g���E&�z<�6	i6^�ޕ/��k��,7/�/�кFP�u�dr�� b2f)Nz��|�6�w�,�7���GF�c�����*�Q�-�:�͇Y׼�]D�W�E�[��e^��Nn@Я=
y������\��H�odr��
]��k-�4�[ă�]y�F� ��BYP�v��0av
�`L�(䣌�Bx�}e�[(?��X�)�̳�1�� E�띦��s�[���NUz��]GPvۨܾ��&ц}�����q�u�ɸ�I�m�%�L�^b���j��u����=��{PK�G���	��#��%y�>���c_tH����`�xQ���R���}'*5��>+����N��6c�c][���l2�_�@+�Q�MmBV��yTe�"A��n�HR���Ϧ��_���a�=:2/�C�ζm	u��`U�n�ݧ�>�:�v�d��ޟKBpP���F��T׶�T��N�]���$�f�v��*|�`�>��l,�zW�~���3�V1�2,�F�H��>aZV�~+���ı�5JS��������Ě�����Jo)3.~�?ӈ�S�	�Q|M\�����oǮ��Q����\m�)#>�Y;�6��cc�d?��zA+p��.��)F䓴�x��>�E�k4Q��Z��u���E�U0�h�7����/�6H��g�g(Y4��q�-�Ő*������7��X��˔��*���Y�}�׮w.�C�, ��������Y���B��(հ[!C�������,�r�y��ع����}���Yȳh�@Ըt����qb�e3Ŝ��F�2�`{ֱ��#ˋ-s�R��pO1��y���v����E��A.�8LC�s5��:��&��/r�����y�������L��sy���^_�����P��qu��V,s���U]�?Z�8�,=��m��s"r�z�Jn
D�7&z�"�I$)�g��$��RGY����!��~����4b.θe~|����D�O �;��'��G3�j�͂"�st]\b(�Y|�s3��hEh��"3.h����Ѐ �"#�k��m���H�Dǋ	�<�Y��P>X�.�8�g�<A#ϱ�W����7��5̙] v·0�Ow�
���2�p��=4�}@��0{n,����<?��3�AZ��֩ 7bp q�zM��m
��g����}Mk+Rd,�B���a� yၓ��̓��s��9M�Do�`�zM�@��[�?��wȄZӃs/W,2��ǫJk�HF�!XJ.������ҴC����Й�P��m��]�XfA����.v��W�1��B�	o۸��,�d�UB��n�?gZ���'I�y��
�cB��\\mt�:�f�������ڍ�139�B�D��5�a��xm[Ȱ���ל"6��R(�_-d3_Ȑ��}��k���y�QX��d�6�(Q��@�8%�!$�_֥%�0g۸:G�tuH&�:��t�l�q���n�	��A�	,����U�N���t=�c�m@w����%!�mI�Y����p�
�N]\��������(�f��G$0\�?��T$-Y4���k-���[i�����c�f���B�`x�u�B�tF7�b����S���������چӉ�g�KL=G��Lܕ �Z��n9/TS?�6v�6�jh����F��y�f�8��C��=�� ��K=0���U7�Z/@�#ćm,�!�XAq/Bjq��@>��Vx� �E"vˀ�Yl��R�e��1�66z۶�����#+��OB�\����D0x��A-�eӫ�x���IS�Bk��'�T-w:�Q��8���}�TZ�Qn0	SbsUv��}��e]�9��\;��'����1��y�w&yv�ʼ�0�Go�q���!rj����aa0���[-��������짻�?����o�Bs� MZ�*�v�~�}5н1�g�	+�rzc���pxd�E9�E�������6J�aÿ��6���S8�b�h���C�3�t�.�se)d[VU$�NN>r��?F9��gߌ�d��;��4���bN�f�ݲVջ���Qg��PJ�vTud�S+@1i�'{��'�]�m�1��g��*�7c��0)w!+��a�- 1z����#R�����V��9����r�])>_�8E�#�ђ֯��o2�t��	����v�&��䏞����.�N��_��c�6R���e�ì��6G��<�>@|پ��g40u��o�y�T���"��,�2��7�[r�a�R����^����:P����h�����ܦ�q������A��ӑr��A�+(/5K�Sd~�vM@������Y�j5|�N�S_�;fC�]���C�k�S�r�P��{@���n%c�1���y�JS�e�Y��巠��W.qΑZ� \HN��}9�5V*\S��D'M������>ps�9�P�u�]��Zc�5��J�%I�P��z=��2��j2��tqg�}�[@u�T��-#����o���+,�������Z�1�����W��ӊs�nb����~�nI�7[A�խ� +�0�Þ��?����M I�@�Z��']��7��� n��R+���A7�y�@�=�KG�Y���{�H^W$�:gUj��}[�6]��� +���7��"�<0Ӛ'�W�f{�j����cHp��lØ��؏PR��>|��V���{)�u��S�.{���ѝF�q���%h�#��
��`����]a�R�'g��Yg'�<�NAЇ�2�!S���Uh�����YY�G8n
�j@�=�|�%�:�*VL5�L��QL��;�C�NSR���U��¹#���JƦp���v%͚�ƣώ{I܎[<���ˈ������z�.����3��q�ir��wS'	ʳˌ����Y=d�B��{���?���G*�"��R׵섔N�,�-�J%O����־����c[X������'���H
�)ٮ���Q����2��E7˩'����3V"ds��dn ��z����X"S٢��2x��sxn�i���<K��A��xΣW
���:W����m��F��r=��z����°��N���1�]N$&�!�Z�^�(?�������`���o�p3���AN 1�l��A��k'c:[&��ӯ��!��w����~3�T �'���׹T`H�-�3=ȼ�"���
�`{)}���3��1��jo����VpS?�� H�	س�����-$�����j�U���E@bD�8��Ғ��eg�Y:���nx��^�����
���ѓ��|�ǹSr��ܱ7��U���_���u�-�Sͺ�BX�/$J����QU��>_}�CjC��/�\�H-U�~����o����qݧQ6��
~w�;�*}7�n(H^�E��~���$����,�u�]�\Y�(�� �%���Y,y���A����U�E�X�XԤہ�b�����[[k�+l� Y�M��X y#33GmX���{'�ϰd�j�4m���7�=e�Sq����EF:�Y?J}t!��aht��g��S�n�}3��G���	���TN�С��������"�9��f�>L�l�n߱��� (���+i�����!�"e��uB ��-��`�k����_�Wo>tPw���*��o�3���<6�,�wX�`4h���D�7�iD.�IZ��ڪx{��t�6j�ȰD���d	�9���,t�s� ��J�W̖�7��Y�L�5Z�6ra-EL��+Mw�hb�{�P&Bnb�O�XP�jU<oX�k���o��y�3|֝����M�����x�A)tsk��$���}Y�3 )�xf�y]��E����T߭�|�'\r��.�?0	���-��m%��b*�Ia9�E\s��^���5�|��Ȅ ��^���z)e�q�z�g7�����6@ #(Ih���:��|����q��<:�&�"���V���&ǰ�.�1!���z�i��><Y�((ދ�����h�+�87Z��ꕔa��!��N�Ud��% ����=���ɫ�OZ��)��l�P� ���J�Fh�I�@P��}�2!7�׳\S��4Ĳ�M��x���)X9h��1-	� N'�ޞ���ָ<ԼV�:�!S��#�S���Bv*���ku��_Z�|�\����i	3�zǦ�s��������F��:qt�R������q�S�4AzxP���|��֥�%,��|�R�d�_�V�.,����@�?:a��ㆧ��'�,��\��e���3�b�XfS���C3�|�8��������N^JB�+;�x<�ĥ���KT.wi��((��7%`О?;L���(5��O�B��s~�W Q 0s!�de?���.͸�$���4�,ǎ�h�"�`����P)�E�U!K���M�����_�u�	&�̜P��
�� Y�)�����U�gP�G J��1(>*�����~��v��c���n�0/z��~gl���g���i�����k�kEp�������a|ţ������d0��l���G¨�^&x8����Q���c !8�@�NөAo'&O�ӿ�r��2w�CiA�p��������㔅/�ǥ�H�Z�K�Ȟ�!�?��yt`��#y�y�X3�	���i����q��h�i5����=W�rI�1XPnv[��þ�����>���}�۟����	0�hɨ~T��Q_~���XC	}x1�.�r6�����#�"e$҇ܤ@�ˬ|���FМ��X�G���끫�p~1�D�;��7�IRs�1x�A]�9i#�-��ف5�� iq7�{��`0:����P�����ϳ�����5$ּ�'J/��3��%]g�i�eB�6�{/�T� _W����jhhD6�*:y��`'_����r)ҋ��.�9RzX�y�!�K[N�]�n[f���%�2-�����)!��f��������,ٜ=�������[ib�܄Ӄ׉��T}7�9}T'\�+���&UYPlg��dg=����`�,������b];^�S�ԽDe����5VY��>�
���{u��w�����'8jQ%�<�zY���U�P��*9�N�L������ne�����2��!Ͷ?ۺ��T�j[Ҧ�/4�<o`��x���F#VW��~
8}hVP�)�y���OA����ҿE�K-&�#�E�.���v��GNK���)�?��Nq���Hl����9л�}���� �*���l]ɷ������`"⤴�����\�Pj����W �x�S�W<��	a�T�c�ʈu���҆�HKq�]���ߠ�3���@]�"W�t+WK�����9��=���q$��.�ݻ�	�����$0$;!�=x�/?T%���^U��T�Fxgߪ�P-��m/��T�	�����7��//�2�XҪ��U7�x���QVS��W�#E��/����6(s�;i0��ƴ18ß���d��%���74����EF����gO���EHO���D��	�8)�{��	ǧ�Y�>�ߟ�>�+�!*bj�������vb[����@��Ѱ�Z�n��Ö��kH��N^9[3���d����-_{v�-U<�_j`�&"6��ZP�4v �Z������?���L� v�̈�]p�6��*h���%R|�:pf`4��{}|!���)9m\�<��c��
�*��.g�4��Y�"n�e\��j��# �p� 2	%,�Oک��? 5��Ya�`�9�$9
"fR��LLoox���f�qH��F�k�g�&?jÇ�����XH���F2?�óW�^�@��n{�=B�يw����__�)W�,s_��mh L�5��m���KE2��`�CÎ� m`�Շ:�B���9>��ht�
�/�I{Ir +1�-
0�A��+ג,������q�$��k;��KmM�ē�~�S��!ƤH|���M�����M�`���p\�4����@�G=�g��"<�}�W��;�JfVx!U�pX�	x1�� e�i�ڟn)�F%�h�*�x��ѐ�KE\ZWmo�7��|�	H�a3)o��1� b(��V��g��V�&�j�C]�I�G��y�w2��+��I}�5��*���qd$�B^8�@�7��XB&�E� V��k�!�P՟�<��@��؝F��7-^Ai���9���3���	y�r��-�߅��j��c�Ǻ�t�$��dQ��ە{Z��}�+��C��Vh1��%�0x\16�����L_���u����T,��;��e��ג@��"�ؘ;I�ŝ�`�`3\��8��P��0O#6�s�"����$9Z�#� r�6��t����m�EZ�O���=)FfHZ;��ƶ�wN�*�� �J7�D6��$5=���{�0��(��Gf�����+���z��|P���j�&o��Ks�6�%m�{�'�lJ.����m0b���m|@r^�{�h��ӑߓ
jd��ȸ���NTk�5E��u�!-���!�n�6Kx
Qɠ�8����Cuj����gl�u�l�]<٭5�]�����~k8���Y*Pr(���Dy�9������2��^����j~m�LP��f� Ő��TqŁi{����n���4�*�2�qEm�z��F&�,��}������Հ&3��U�Н��$&��\������c�)��%�ФK��P��B���D��s�jL��U�g�$���P�Vܺ!���E_C[�@��HR�~�lʂ��z*��QN���O�˪�n)��ߗ�|�b1���[(ʵ��h]�l����;	�d��0\d�}�@�m�c�%a��T�����JYn�j���<��b�.u~mw���M�	b��W'����&�_�&��L��g[�Kܿ�m�wܔ�2��?L}hۃ��묰��B��>�%��SJ��H�A��&U8��ޑ���1!k���1恂ܱα� ���&
�nR����չM�_����K2B�����s#^aMc:�x|	�,��s�y�\C,+VE��(�K�~|�3�\U&Ȝ��F�<]!Y-���^.NJY\��\aè�,���]�hy�����>Q\�����Gx�>AO]a��ѫ������p*�~���G�8�sj"j����h\��wM�;�w��ra�n�$T�0���_`�z������J�� Ysf�V`ꔖ��0�[�@�;�W&��8� �|І(�Q�t�a�G�{l���Yn/G܎��-���l]�b��t�.�97w����. �]�n3�{?�v}3�8�|�����د�3�w���q��ϊu�|�̤:ncBʄ|$_��P�[�
���H�Q."8�t��
 K��i��ճ���U7��e᪁���+�ݣ7��<4�0lq����~y?�^5������g�a=�I�z\v]'����K��Z(*qs���D�F���p���!�􍛧���qeH��3�����m#ȩ�r��s"�v����'�p\w���t5wJyG�n�:Ȫe�-���)*�E����T}��jiC/^�$�9e���q4W�������r���`�5���<T�
�K����eT�l?��(�m=ޮJϮ]�E ��9g���݂�S�p5[r$�g2�
�BQ1�.̢?d���  �-�❿r�0�vW�A9�ˑv�V<�9u�%)�9��j<��6��P5���(�_�|㐿�W)g��+#
�a�/uz֧=[�ɛ�BU�|I0˽�C��jA�V��ˇ�U�a���?tD	rn2�	= ������zHc���5�e�O0|V"��� ����SÂ;�M���)�`@�~�{�O�=�W$��Z�Y�&�6���,3�����'͆��tA��&J�"�>m[� �kM uE7j1%�g����<6�*�˓KT/
��{� �Gm�d�#��K[]P��P��!\�f�1���@�xH��c,���WX�ѿoHW�k�8�q㶅}��	�*ɺE�Aǵl��/���GF�??�x��T��X�2m�	?�-�]���0/8ƔK"o��d�?�^��ٺ��sk>�jmI�&^e�A�U?7MM���\S�G��L'��F�+r�q�5�g�[>��6nx��m��2���TT��z��Q�P$�5��;�ޢ�}��#՘1��%�����Ѕ�Es����%Y�-�5>v�2�xG칖~<����h�鮕.����:N+��=��/&Q�N�ߕ{��x��9Z��J�?�-��=�^�S�}���hb���m>�0������@�	�����jR �j�Zs�z)=��5�L��`K괮(w�,�Gz���a&�b@�p��D���l0�-��l�����1�iS$9��i.�7�p�/�oY�#��Ѕ2R�(:�ZC�x�XHr�n�O̤4$jD���
�;u��-q�Y��K�E����梚�!�((1 3Lj������� đK���ȝ�^5�ب̳�х�a�:,�i���~'�e2C��vD���$e���i$��k;�{>��&�=zgƾ���]X��s�F`�ţQ*/����F%�{��	�?�?��g-
���6��!��'
������'�o��}�ޅ-��Tܚ��"�}�Z�e`���y����,�_-�v�h6�x #�$���e����%�hH�p̶�UY���ak勏V��e���D���Uo�n�
`� <�08��d�޶��=�8��(�ז���B.#z�0I�IZ�,O;���b�LŒb�*r `(ˤ�*���	���~%��^eW���[g��g�������dQU� �rr���iOȠ=��B
�gan�dyN��+�M+����(J�B�!�����ʘD�Y�����N/�Y��*mR��<�2Q��Ӭ��~���s�q��K�s3�Y��@/&M��?�>����i3�'�fin��ݓ�>ɛ��=H�<
�٩q�D'w�>�Q��G�y006CMR�_�V
�m^��L11B�s�l���-9,�H��x: ���6���t����f5Ǖܪ���$3���s7A�@��$�2V��F�gʪ�SЬ�i D�٘���ݬ��*���}��6��-.?�"}�4�^*���d^�khG�$:nT�����9�tE*9�Z���J��)�B�a_bw�C��@
\,,�]����q�P{�h6,tك�#��2a��������+ޮsJ�5 �1���b"{�]� ��*��Nz��5vu�Z�?�"ڜ�������?<�t[i
?�S$��s�@����}���Ɉ�1�Ob�#�ƭ�9�6�ֲxc������������	�c���,�2��xi��E��@3]Jua��VH��,�>����y���k�+����qF���fX#3yc^��	�4�u�P�6���,Y�,g>�R�Ǌ}CKW��rMw����Z:�\<�� oB��A�k�Q�#��λ�D���09)?};�����u��gd���Q,�؍���0ɛA��d�+�4���V>�DA�7��*�6V{�v��a%�t�A7��ʓ8Z'�༄�����z"1���!:�S�P�E�H��Zaψ;���O��~ʶ�9B�@���F�+A�Ւ�z��X��P~5ο��ӥ��)+|9�KҮ,�1�P]
� 'b�;7(kc��tbr8��^Ko:�ȥ�崙�
w��Lӄ���Ӻ`��d��wfup�:�F���:�bJ�lr[�B�J����1���M�|N{�NV8�HV����Vg5pƨfہ����?q~8r詰6��_�0����B��Y��h�����zlP���(�fRl}"�̃.1V�@���^}g�OB�\��R����O����7;�9r������ۦ`�4�l�}�5=�]p��4�e�x�2*!�#���f���ot��C�Y�2GH�l^��� �%�.�=m_�����KFQ8X�+K��RX5�&��r��VeAT��U81�d甮^	�����> g~�|x�o��B;��!jb-���ϟ��U����ɢOL3�A�������.�bt�a���W��~��%��oE�G��p�aG���--W�4��F8AEM�����)��r���Ƒ�(��@�{��_�$&�u����(u�3�2����e=Fb?� �J���u ���T�	O'N��5xnV�܊�֜&\Ǧt��� ��_@M�x�:��Fc�Q��r�0�8k,~�O�%;���k�7������源�� {�"��6ñhI�k���P���`voP��Rs�!��c(h�G���
/��F�^�Kb���?�:�o��W��H>ֱ*���
�]��d˔���v2%�n#�'[��b���~E�#�=�E�n'u��!��+�26�Y��%���od�%�**׭g鮜�ٳ�wQd���H�ì(Y�֋	�ܦ_�2����f�/�+��e�ც��M����R��8(�D����k$��������x�m���r[�K&NH��2y��q�X\c��%�J]�E;
��PpL�c��}�~����m�iʡ�TE�o�+L�X8�f��p�`��_���K/��ڒΎ/1���+�7T�4j�d0��:/����h�USs��vq��3a)A�����t��!�&��0H�|b�k[��Mn@�ጲ?�ȴ�c/ҽ����Gӳ_�o��ޣb��GGA�����ύ�l�^��J|oAb�E���.P�ˤ3�VՍ���Ul�ddwZ���t�ӌ �*M�� A��+F���G��Y�P�MZ^����A��(Kʂ���鋖���}ʣ�䬸)���m�f����/k�z��R(EF�L��T��#�4��+��wH�=#����T�C�R?ISc�������F=�l�4���{:��v�uk������H��J���.������`W��ͬ��a'f�I{�ơ%�ꍒ�>X5K�-�P����kqq{������F����-�c�et���q&yc,n�ͳ`f�f(l�ᧇ .p��5��x!�K��;�X�:#����8�1��;��)j؊�tV/M�CyV���orb��W��&��C�7{Gm5���J�x�{�txb��߼�R-��(�* �l���~����Q�{�I��2]�]��"F�)wD4�B�*!-)���]o������u�/���N��2������?�h�uut~8���t.���E���R߹+}�R�eJ᝺�&kY�&O��)��Q|)���A���'ۭ=b3TXЊ!2����g�=Հ6X�K��.��ў���8w�;E�*.�sh�̴���<��=ԧ1t������8�㾮��i��S�O3Õ�4$+��?��q��x3����Cؠ2�g^`�z�f�^doE��OȎT'#��������=�BiV��K�Ƨb K�R��f秣�IHy�&�б�']f|��[F�[�ii�Y]�BܚZ�R�R]ds?���5m�b�.�c���bּoN��MHP9�܌x"	9�o~����ɱ��䐿@NH��"�XC
�/62-�AJ蝿��J1�ή����L�-�7D���7����p�#������︫ʵ$�����������g���7%����=��C[r��jju���u���I"pRW��6�0NF(��=�f>���O|��27�	c���K����a<���x��J��]m(r�^V� Z� M$1�p��?�1is�ǧX�j[~x�U䧘���z�0m'�UO�\f������CyL��Y]�
�̐�9�G?��D7�n�;�Y�Q�]�Y/+x�8]h�Q��i�����l�������
�f��i]y9&q-�Ƙx(`��V���RW��Cw��;Z�������V�J��t�8򁮹7���I��h�t�1-�9_�C-]�Y�g ��^���-��)+<o:6�j���0�򓘲Ѫ�n<M|��A�۲E%m��gpO����fx๊7"��%�:ٰq�";��f���`�;���Cb�v\���<jL�O�=���GO�	�2&��GcrԵ;w���1�l�T6�u
)���:?\��7Co��"�J7����s�r�0)]�̮I�#PG��ˊC�k��dkUc%��^<Z_�WN�XMV�{l�%�^�*���G�9�k��
F@�v�E��H��"�d/\<����\��-�űM�!J�"n��,B�rS<.lC5 �5����(4~��6����N�i�������6��?��7��(uejuIM\�F�+��G?%6��zϐ;��`Όm�N(i+���NZɫA��y[�����L�1t�V` ��9v7T�4qit�#����Y!n�P��.�˯�>SlZ�ٽӎ��'9����;�0�E¨^Ϲ�7˼��rX�;;�3��$42$��ͧ~=Ic�3��`�7Z�iu���v9�j��K��3��'�����}�Nz}�b�)򷄳����{��f��q�z����}�	��3�H��1�o;�L��7��s�EL�
Zfk�a9�w{�h�������h��M	0��0T�`�2�B���j�z<�G� W�9�+*����W����x�������jS,#5ϲ���JW"gA("��{�B�M��c���vV�#�G+�v����"�B���tyK����y�I��m�Q8����-���3!ygg�#�֑VN �Y�.����/��c���& Ggˋ'$��E\�XPE��\��rz�Q\Fn��a���4m0C�DD<߄ ���}���o�y�.�,Wz��"ފ�C��n?������)��5�G��+�1�ۢ&pg�?F�$�����C��7���/p�H��^qh�w����2sf�Z�ׄ�{��"� ��́.��[�9��`�����05��aD�O�:髻�_.	��U�|&������V�e����º�%��8ީ[>a��J��{ґ�l��N�oW$*�8z:�/�c��&�I��H��5dҐd06�u���z�{a�k����/M���c�E�L8�����բ�D�Q0�AHP�1v��D aI�7j�z�1@1��#���C��]��k}!<�(g�j	i���j�M+'��F0���Z����)�D�A뾙r�Q�d��j{M��6��H`�T�V���j���ɇ)��n��¿�$���/)`V;�L�=HZ�/	� ?(Ҡ�)#PK��s��?Yg��`Rt�KI�|�6:���v���0�.�͈�Δ��8\'�7�<��Q )��$	����,#L>� ��(�c�1w�#�O�%!��0͕T~WVo�$�]����V��u#�ܨV~��nP>�ge�\�֣]�������hU���]3��"���RQ@��Я��D�U`'в�mr��4�|?�;�e����B��ƹ�Zg35`����Ƴ�R������"9'#p�2g�$��������S��:�����q��0(:R�lNP����~�ؕ8�d�����PL&�<r�����IZ9��82y$26��&��V���A\	 n{v�^�1+�u���E_�Z+��U�& ��7�90��{��!��	��H"�)�\�����K��B,x�(������[����czD��m���^��F�1Ҽ*33E�4�=��/������}�Ul���X%�^m�bZҏ�0;k����}U���p9��{uqo��� ��Dj����]�4ǋ�F��{W���l��#�VMЄE<U����� �dݞP��$�t�j5��bi>��h�<J�������19^6B��#�U��lv�qpW�q�'I��|6�Du3x�������t�j8c�Tq���6"h'�I6 t!E��\Sf��Z�!������5
X~����ZA�Y���<�A1J�=���zP����^/E�X,��k�_P�#��������i��˗�����ד������ȬD8�aj�f��a9_�?hy�ǲ&�k�E�f� ��x��/�
TN?����;��JUe�g� ����,�9�e�$Q�)1
�.���S�RԀyċ�����i^7���ŒXV��B���ᣛ��CT�1��&��[A(�˛��؎�M�2ɗI�mʋ[�t\|ˢR�S39�$Цr�x�2���b�Z�Fy��
c�栅$���atS���6Cw�R�9U����@`�	�lȳ�Q䭓����:�Q���$3#}��=}�D��Bxn`8���%�+�&,��f�w�-�q�q�T���,4�ƨa�����ލSO�)
gDd�L �Lg�U��V�E^!cA�r,��9��4��uC�8��@u�:!dA�z��{��u����X$
Z�Ʉ!x��M�{�x�?��i����àM��O��H���$ؽM0}�+o�C��<;W3���f�ċ�g��6c��󈬼	�d��\ɓT̿���c�C�r��O-3NF�o�:Җ�C^�6{Şǎ3ai�'%Oّ�Z,�ܞs[C)��B��?镝�ƪ`���D�̘�h��G5��xp�D_�X�L��j���&����=~(���֜Aq����o��J0���)���h���2�=��U7s��Nn�[`;����
t��'�8.��5
��ӺhX�r[����1�Z��[|�1�����_(8z�k"j��泰˄�I��4GA�\��������kI����,�Λ$�Ep!W�jKr�2?��K�=!������5q��w(Хr�m��4�*<�0���1kUt�D�������M��=}�Kb���)�YJ/j�#����h��v/Wmyx�Ҿ��̇@a3��������e�I�3Q~ĵ<Qf��q��`;�\D�iHzE�b����w��Э5(�W։'�l0�I ��1�-�SZHΫ�i@jV�w9�h|�Ҹg���EL��T���=j������m�f���2�柼�B�� ��3:	�B�](F^#�I7R��O���a�Ag�-��u��}G���D�M�� �x��B��N��jĀ�:8vtq�������L���3%+$WV�%�%�'d=������I�n�]L���8��	��FG�J�V���7�IkIgA7恟�I�в�{���Y5<�h)#�ۅ�h8������Z�n<���/p�W}!w�U�x�=��x�M��-�K��'����f�c>^��t�d'9�@�+K��<�+��F)�
p�Hm�b�^��cp~I��<���cx�f@�24J�I�㌪%=��h'����H�F�x4� '�+!q쯼nSo�W�PST#�4�<5�����-��(>,�K���Л����Y6��3Y�E������G�s����)�9epTH	}o`�Yo�m�'�iu�Ŭ}��I���c�^t��z�]Z{1�&����6f�ڐCܶ˷��@c��P��WЩ�1@��E�T�W`�z�^�Y�t��:M�|g�r�\���B��1lB�8VLW��͝Ȳ�$ O�8�h`︢7�������� zO�Μ˘D��LѪmӣ��4t!��##O)�b4e�>���`��^�ݱ5z�b����Xvl���Q8���+U6�|�)�R��/�P0/u�x��8jM�|c�����͢9C(ď,��X��IS(l�%A���Hw���6x_vF�D���i��k�@�afG,�L�DI�t� �?/���o�X�Ű�n�dW�4���b��r)<u�3��G�Jʈ�O�f�R&�Ԑ�^ ���"I޲��/C箽;۷h�Sz����M��6g7�F����4u�������^����t0�p���\%}}#��ݼ��Wv�8�n�dG�S�"�\� @MA��lu#��gI% S  ���sl�=��*r5þf��.�C)��W*��ae'�z}HL�(��ܕb�1���I'f���mY�䮟��{�ߝ@"E���'R`�HˈR@R1�GM6t�v�Ɗ��leS� �e���S��7�0R &��6��X���׼��Y�i��7md�rz#QS״��_@��KH��QYN����=��Z{��A�k4Ľ��ey?�Y������f���}����q��ϫ�Z�� �6K6�����/!b ���ui�`Q6�:��<���:5U_HT�a��Ԑ��cEcUg7F�_9�ٛ[�I��>z8475���g\���1�)xؾhw�v����@A��т��ɡ\~���H׾�>
�ۛ{e���wW:����p�J_d�Z�,Q�Z��̇
aȪs�U��i���J�$�}&O����g�s{ZI�Zwz���.z< �c���Q�ʅ�8�R��=>d0S:ט��3eH����K�H��e���Э� �����������ؙ϶g�󉽨I�N�M�7�~�y�
� �:���u>�
d;7td�w�_�9�؄,o�M