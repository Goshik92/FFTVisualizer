��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHnǨ-�8wV�}���� N�L2{�p��L��� � L��0];:�G�����Ü<�3��jTЋ��2�ܓ��@i��T���V��Vnj�%���k
6�����C��u@��og��F�XNd*�n���!{���+4a��mc���%Η��t�Ԃ;h�2�_!���]+.��S�����M��_�{<��Dw-���+�8)y�/�	땄�B)��*�fE~ޭ8�񍵹|��VSiH�V���" �F�L�cJ�~����ꢢ76K/'Z��u~4ȵ\�D>4uO�k�&��.�<1pT$j-a��і=�%�"���5h�e���t�!�}�y[�f_�-R~юb���!mZ4���'��@��q��m�QĿ��%�>��<�"ۨ���O3��,^^4q��U�LR�a�@<��^��3�X �w�W���)Ń͠6Y"^*�/�}߳���Q��N��ht+We|ɏō�� ^g�y�i�TXԕ� ��S�T�7������^�E����rj�VeC٣�"�O|5@��΢ײ�v�t�@�H���0J��X1Yuq_��.熳�]i�а�g�u�������`��ykJ%+��$����3����Yr�L��v��ʰ�]��R�㍵�i�Ɍ��8�)���q��>B4'��g��HQ�����K�J�2_�Q��:�ueK����w�Z��q�;Z�A-ah�k�{���`�$s��x���r�G�5�/�j���ǝǮ�2��x�������G��ʽ]��̖���`ix0
�~��I��� o	<X��ާ��U�Ÿ`�`ޤ4�#~��kΰ�V�(Ԉ��p�@J�ӄV�~>e���G�E�v*��e/S�i�$D��,�c��y$�9�xz`#=r��-̦#C�F|>fڻ\qt�PJ� �Bũ�{�ՠ�O��+��������k��JBM��ƕI�����a]+" go�!>��)�,ܤhв��J�gl<�E8ċ���3��:�O��G���%����}j���&�g-K^6ŝt��͂���7p�a��De���W�b������\�7d�ך �9�d�c�k��`oX��K_J��L��q�hA^�6�9}��X��C�r�FȔ�G�B�Vr9�3����Q���	�A����'9$ *;�2l)�ӣ Ȧ���d�xk5I4���%��ÅE�S�� :��<�Y�����.��;�]�[��,>7Oų��8,���d`�n����Xi�t ����S1�%���3��� ��� &�Ũ�_�yh'y��hv������C�
9h��r��l2П�NJb�0�ыލ<�^�[۷�b��|[%Ӡy��R�+1�FD9k�ߕ�q�1L$�GJa^7 ��򧵲��$�Xݴ��X���16p~�y�ںE�:��Q�l�wo~�0� 	�V@q��}�S��y�U�ۜ�L��
\e���E>Qg�Ub���E�|���|�o2�m?��H��i�O��� � �<H�g��P� P�������%?��
9�;����$=Ųo�⿲�fҺ�]�~�������9ڦ��Nd�	q���ظ����8��[��qKWLA�7�?��BK3��'r~����I!Eo������pÃ�avL<�a^ѓ��vD��ls����<�����[�ol�+tO�M!�6C�B��*l�'�S��0�a�z'�3ڰ8�>#b���r�zQa3M���j�h̽�D���8%����Ǌ�<n����6���߅P����0��)ǐ�y�d��;�j�'�s�'Tpw�s"L'X��/��^,^*ث��1㧯
"}\L�R鬲~ذe�J:��]�Z���?a[�hc�km�+�Ο��}}:G'S	EKo,�X�tb�M���/����u_�e�����=�YV,c �$mBs�3�&��Y�.���F6S��R1�n�s=S��r��-���.Aᣦ�Nd7�='�)��5�Je�B�j[Z?���VҺi(R3Q�x3���\�~�!�젖��O����
��L��!\�ob�!b�a�D��L娍HI�Mb��q�\6�����c��خ;��%K�Z�%��⾦%��+ea�1G8	Yh�301��f����;���m��Ms˦��Y��v<�fn�u���L�v�Z�k��_�W��&�8��$A���6$�cH"�}"�Q�)Z.������L�pUiy����7�77����R��Lα���q/���Ul�U�x���%�Uʅ���o��Y�[�;GO#Q��{�$�Q=��!���K}P67+�L%�B�j4mY70��9*`Md��e�(!�?��㏄�X.�I�[w�2E����Yd�vu)�	�J�0�ɪK"�|�I�CZ�!%e�>P��i�	���l�0cT�誗կ��[fnBZ��9MfvJ<�'�aj�^d��[�`s\&��#�{3��YZY�}��G��e�Xhb��n����?�Oc�gV�a�;Y�������
�L��j��4��3�EzrG,A�h㢩E�:6�����H��+!?�@�ds���ܸcT�88t%���o��^�
�8��_���(?e3+�g���}0���é!�P��
F�B�/[�!��d��cO|l%-$V89a'7�H��b���Nr���Џ�Fɶޝζ���?����w�N��J�J�G�W�.F����'�g����r
�ޤT�J�v�f���q+kB��@��c@+��)�b-�=������ʹ�o鴜H5��>�K�b��|�u���&scb52�^�ϧ�d�5x|�~�=��(@�Sk�����?�H3��[N�b[�.M��r��������;�C�'�ڢ��zˇ�2�ԔL���z^���\7C�������<rY��U�=��8�#�u^��OE6T���'*- =y�7��m&����������drh|2'5��E��������2_ �ȋ���D��F�V�������ܨ6�l���EFi]��D8F��q>����%>w) �<Q�ɘ8��Hr�."ÐG��UM�2l>���,]�ט�Gl��A�d>G�eE�|�9s[�d�8�f��s��S�KNk]~Mw� �+��o���*����i�E�o-�Y2_����I(�1 �y!����VD��3	W����t��T�Q@Y�Bj�ն���HF4cdW+�I(c^�z��*t��ci��H��hL$X;�)�@���h��Lf�zq����F�~<\.�fZ���Y�0^��@�ָ�p����Gk�l��W>��NJ\r�2�#1Ǥ�dp���7)���HN���j�y5�{�Vc,f��`X�����R��Ŝ���ݷ`��.C�KB��uM7`H3� �A�k�?N�:�Qs*��?[��߈�PwP�C�Q�Rٷ1j�2b��|%&^%�L�c�]�r���j{�6m	_KO!���e�m$��Wn�9KB?����44��߄0��N�ԫ��Y,W�R��Pgj�d��?�p5&�J��S'T#��R��(Lb# �_��������Pѿ=F�9�/@�Dw�Ҕ�i��}#}���\z�uat��.���DХb*�ObH�
)�=��JŨg�z>�q%S�k��o$��d�0$�_�4��vlp�:�";L�>�Fb��0beH�1�\fH{�Z����k�rf�\��L��Z�	|�*J���r�,�7�E��d�U?`�=<0!�k(��
k{BX��	��Ǧ���U�f�61>ɚX㗉m{�{z��m�3L���<D��r#��6��.��m�(�7��ߣ��T�R������q��Dw�K����c.�CZ6ʦv��R��p��G�ѤQ
�`5� �b��k����&��FL�Y`f(]�*-J��TQ��V�!U$�W���]�Ħ�\�J��������>dC*�?X�6����<~E�E%@&"F����l�*��s3�hI�r@���l8�.W��[���@`ԞG�L��F4�qa A2���M�[#09����,?����2Mx"�$�����}�+H����,�h��L���~@k���'(Az�0X	  m�7�������{��56�P�}�:�v�����eU���Ĺ{n�&aYnk�_�Ct~&l����k}���������������^{��,[v3�rbYn�2\\x�ߑ����E�M̘�>��t}����Y�U�T�m�ı������\�Z¡���j,t������vh=��"�JȊ;��<ʏ��u�>(���A���,���LۀF�R;���s2�Y|݇s���%\3?mh��tM��w�R.�O��"m�d�Ϥ�����ڤ4����e�	_H��n���n_�D%`��q���d+�W7�&+ Sެ��8m,�K�FS�rN���,��«%��6��A����}�߭u���^!B}?���;�Cb'��D���<��5/wݫ�*��o>�@�;l/m�r��c�akH!@�◁��%p�B�a>qQ~��/J�1�o��k��`�Yb��K�5J��ڴ�1�x�`�7L�}ȟ���铢�M�g@K�'�~D�B�ӥd��n�2�D�S��[��7jU�ֽF�*(��"V��R|����gTt7T��GH?J~���(\�l�F'F(u&;y�t��k�_�}��,>�����R��,\�V
S h��<�G�~I�h���8�ZZPg��5~/x��H~��%��aL"l��nuOG�ժ��&G����'��6܍�[j ug/��m����W$j?뜙�	Ē����M=�@FNcޛd�)⏱���f��y䌃�>hm
yoL�~��d��`�D�P �Ђ����|_S����,�
CU&�XN�@NWf��vu(D��CQ2pD�I�ޙ:��)͂���6HK2��c�V5����P񚵅��b!`�R��T�Ϯ��R�$W�l�c�<�bڗ��V4P����k�͡$��h:��~�������·�-\�T{�{{	+l�#���ߤ��U�A$��V�; ��-}�A���	\1��'}׳Δ� �6C3�H�)�Q��N���D�_.�m_���O`�K�%���)	 ��[����?E�6��'h(���n�?�`���
s�b�A_4��KD�D�`p��
�sW���������U��+���*�A�t��#ck�6�8�-�9�MW�X���R�^B?�:1��~'�j:��Ctq3>{�kl��y��A+�O���V����Ox��TWd����,���P5�4��&{G�d;������/���o�����ɢ�����|�G:)�{k.�pG�9l�Wd�����5\f��D&v�[���������$,��)�h^�J䙷�,�����ڸ	�`�
�9�?����ޫnP:�����펽���I�39�b��Ŷ�\T�u[2���J41Vȕҽ��V�������%�W'�Z`��A�r�����ʠl�7��s�g;�U���MRl�`��t���E~�ݿm�K�9�P��y�ت$o����8��C�Щ�q��xFl��r�Z�v�t�E�7{�ڟd�~�"r�y�a�7D
k���u��\��T9�������9�<��h���۳{��%z�|A�V��\UdM��&kz*0�_oX�4�ʯh��P5�ǂ���D�=%֎<8�̈@��]"F܈�f�A�r:z���tǠ<�J
RF�k�b"�GNM��"�ë�������J�Q���H�L
����^<�X�M�pa�H��ҝ��G�I~�@���>��<��ﱭڐ�"'65�*� WwF��+�#Ldh[�����ﱳ]J:l����(+Q��� ���r�U�S���Hn�Mj�R���ߪ5�|+\4 ·Anr�K��	����4r_�ڞ�Qb5��ql ԍse;��aN@*������2@Q�EԜŽ�d�(liV�i���hl(w�FA��W�v��1��$���ҿf����\�T�d�7��I��I�x�le�E�
��_v0��(b����\Qi���"�a{j������߉]s]p��4!���<	#q���H8���>�����tׇ0�N������ ,�-��{ ?XE)�F5���А/Q�!9�+W�n����(k���ȋ�y��L�A(w3�=��3����i�YL{Ś�`ƹЖ�W�١���Z�P_��Tt��_J��C����H`�B(�����;I����Ԇ%㶲����q�@�K���$�sp)�I|@��Ó���/�<C��U����� ��"��M��J�К�\n9Ql����p��P��9g�H6Xh�|�o޸:m4י O�����Δ�M�ۅ��Z�At�1����P�(���@���-�z/��I���9�2.d&a�M${�"��	�]���~r'�0ڲ� ��4ok�Y�c��Z�J{L5� ~��/M���Y�{��{��*�E���"ld���ۇd�hB���6"@S�}O�-!+ʃ����!Ѯ�Ҿ�U��P�ok��Y����d�t����C�\�G	�r{ӻ�P�:oz�
jyb���%�aX�֑k�К	�zRx�����)3�����o!�pßk�P_�rE�N��j���0�.��6�8�,��2���9*Y�_��16�!��^/1'P{V���ᝦ�*�\�ww��#f�N����J����/�`Z6�|#MGE#���(��%rt�~���q�Kz��C�r��LPq��ځ�獆BN$�=h��􎉳BC�N�_No#	nuQ�r��X/����ni�~�ޅ4klc_�pc�_�06XyK+6��b�:耑�1Z�Ɨ?�L?�L
�Q�-����@�l�O���{S���fz��q)y;�R�<Q�!�d:�I����xo���!(��ǁ��0���O�ɬ� ċ�lg�������
�`icOªڔ�5��ɫ�cח@ӹ]0a��zP�i*�eC@�je�\�x�Շ&�^����q5a���MC�u�K�fɛE_ V.uM����-lMf{��S!Ƈ8��+���Hਕ��/Kfz�M?j�7�L�����'�P'�=/*W�[�jS���S�T�[2naSf�ɫWc�FD~����+��d��0��t�Ѷ=v\������'����$����"�m&F�ʭ�v=]�c�wJ,���؂$j������y��Ӊ�J���(�l<
@�V���{o��eT}	����!>/�_�d���A��
��j�h̹�_�R��7��UK�Kgb
�'�Ed�I����d����=�1�"�
���b�h��U��H_.P^��wX/ͧ�q����UA"]Y2���&�S 3�l{�@�6�8Nc�S6����5��A���c�|Yy�.�i��S ��D[���7MagWh9�E���!���,'�-d�]��G��_W��	��!�	��K��GBr
%�&�U�iY)�4��E������I��Y�����D=ʆ_�d?�մ`�� }�Z�JR�����>"�kK
Y�.?�܌�Ợ7+��q���G	��S�I* ��D�l��p�4j(�'�[���U���T���fa��8�b[>�f,�E	N�$��jj��-��*��A-B	�y3�W���[�b���K6��Xχ\ƻ�iw��'��#~�vU��~,�Z������Q�誯���] f3�&F��y��0��C�.�ub�>nD#�����%�Y0���	m�>R� ����P�L$Io`8���4�4�
^�E�G&9�n�47ȭ�ip���e#���-��8%�"$�w%�]g��J<�����|�
�eUk(�dI�	�xSY�y&����%$��,Z�v�"���q{��&�d��ژ����I�� "³|aQQ3>T����9�`�N��ڐ����&�м���;�8��p|��Z�>`{���8�5YFd��'={�&=1�ۋ�1��{�>͞�u*�r���q�D��Ҩ&��o��ޟ�/�JjD�+vWY��*׺sgy
N��n��]���冠��;��L9b��@6��5�y��w���W`[��
��	`���z}�ۓ��ض{��}yZ��ߔ�E��
����ũ�'�i|�V��ғs<�_ ��h"'�Ce��y�x�m�%7w���E<����C�'9�/�b7 *��ɿ�cw�o�M�]\�~$�$A������7v{�%����D��=C�>d�`' �&Vv=0Y�}��M ��D�g��K3��.3AT��~�Xd��P�����SG&�;�'��qhf���YRs�/��&�4r��4b�B>Iۗ���u���yB�G��ѩ���巬V�;�;.��g�:�@�(�|-�\>��E�r/����z�Ah���vG0��\R�����݂�p8ß�TdT�"YWqFf B7��?��	��	��ÐD2L��Dp�N�3�u�Q��ژ�d\�N!�����"e�^� @���;&�P�sz>��إ�A��.Owl���eV+z���)�ZF�ԡ�����k�S k���*	�L��J/pǫ�"��g]T���le�3�_�^��hq��J�cp�zF�M&�y�r���3폺��gX��o5.�pV�Ps�Sr�>����Wi#�R���f�[
<7+:`��C���)�8�A]�!K"�1�0��L�a�
�ý����jU�$�a)� �PJ������GVe#S�m��D�xFp���coN�G0��t�5��S�ݢ3��C����i�)�֓������{�i2"A�I2��(����sc8�U**v�����nA'U��ޡ�vl��<�|ȗ5h0X?E=3�jm��+n8c�:��L���Դ��V�� ۋ7�edH���$�� �G�&ƃP��u;�7�������N퓔��9���ewWh��������W���0��?��m\_����k%[�v�\3iSk�ԶG6+��S�������%?B�C=�gO��F��U,�XR����u�0�^+��tɞ��u$�����mvog�ғZ[%ײZ�7ξ.��NUz"�Tvח[!��Q���7w�^?�_���v��R����#g����O��7^MI�׈�ӧޖ���߃�U��ȴ�tԾ��_J��O�������'�(.*�c����!�l��g!	�xP{!��f�^�����!�g�
����֢"�"F���,X�E���Ê��Ǽ+��=mmfţ��)^��������/�֧K6/���1`;G\RLG�	�ti��7hw���3��S*�R��������:�8^�N��d��ɿ,�蜛��+������
NoiK9�<�>|���D�hjVV�W�bX�������Z��a'l����`�{��%E1��}���{��2&����9�~�tU��K�0�C��� @�1u��x�ZAP����Ύc'YW��;6��Y°�[��"5ٓ:a��.�r�՛˟�C�u.���f$k4�T�YN���x���6l�4FQ���%8K���p�[�S�*Q��1׸GR0"�iݕ�q�q��}����ζ?�V~5;��hmn������<�>.VA��d�sb�X����E/���m��֏�U�m	��[2v�9$�
ֈ����c6/�xS��$  ��2z���0b�0v��[nv��L,�M�B�>�
.3���dJM 6�^���N���O��c�i!NX��S��&����}e���qu�pC��=��#�QX��֟!���ٹ�\�	�����wS�[=�!B���]3ߌ&eQZ��TMGVƂf�ґM|	�jH6�%&Dtb�����)h %[��@��1�,gg�}M������ P��D*
|�\:����#7��J#݄�jG� sB�*�
E��<�m�l�<�
��_�,��K����J��tQ�N�JG\~��M��ET��\0J����7AAsԎ<�	h
��vDNj���Mx����}V>�P��ҲU��2<��`��Hn�����ۡ;~Le�ѫd~��f��s�r-���^���'�> '�C�c�i����W�6q�%$��[����T����@`����)&,��Y�W� ��Hm��e�z�8�ȔK���]؀���!o��=Q=]�4��_�}��-Hk�i7�5 ^^A�E����Y?�����i�KΥ�eOLa�*5�2(�h ]��~������h���hng��xd��6G��nu��"͖���:�o8ҙ�Z�g�~�j�e�_� �����y�S����c�&��(7ȃ<RŒ��B9vi����0ƿh�h�.�T[)ߪJM6��(r_E��y��T1�]�}�,{��}�����=�*q!HBH�A�4��6��`N�Τ���0t�9���9�)$-���';�Q�mDp�Ff[�5�N#���UqJSs���k��/dx��Uns_}�t́co$m�`9g:�EҗB�Ј�7H��Bڷ�6;�[;�A��`g�9�tw�G��Z���M��XG[�����~�o`'���n��̻�-�s�,l��8RmV�Q��؎���hGO�铷�����Y���CʁJ��;!�����k>���w;�3������~�;ԝ���H)+����$?anf��7S��q�`v�ԩ����*{6W������g�e��s/�{����7UY�
��a�L� �;����X�.� P����VD5��g�Ԋu���~3Z���W�8&Z�%V����������+�L��:����[��&�jqW��Y��ނ7�+�;�߻~}:�� �	��o�E�+\쥙>ԫt���3wR����ÈӘ���x�2E��pJ�0�#d�F�\F-��t5�����;��-�Ԫ�D�4m2\	f��K��ΫK�ת�D��R��E�C]�. �XŔ��p�U��L�HSK{X����p�dD�#���y�<�'��6���Ox��V�7Os�8�D�E�d:Θ�������7��U<_M�ׇKe(H�
��]�y+�q�~��ܪg,/%�Å���M����oZv�dI>�XX�\L6��J�j�M�bn,�_,�� *�u�."��f6�5�;��QK� �_ ����PƢ���o�%])��!D6�v�g��A&����3���� �b"ғ^%��hӲPR��;(�Uc4�R�ؾ3���ᱻ�8�T�Qgi{����(({?��'��V��7/9֌�����6.+�qD$(��t;ٱ�����m�<f0�V��a�Q���}Ȗ�b,���0wi�2�KS��s����p;���"�I���7�����2=��v ��M�&��pS�����	�r4���s��`���I*D��	���C�ry��c���Q�!E�z��԰��~E��m���sj�A�0Q�(=�(v����YtBo�y ~-�G��x��q���>�"sdɞ��Ԭnϗ_�EzP&��4�uOdZ�U{���&�sJ�W��}�RtW�_,xt�����@��Oǽ��a����1�7W͠�76M��3�"%��m6��Y��sqH���Z`і�8X��o� ���ȳ"�y�pw�g�."t�Z�����kF��d�D�t��~L�痚Q��"F��ί5���9��h�tt՜Ĵ@��zQV��H�c�Q�\JBg'cj�RS*�K�=	���К�����F,Z��OL��9��E����m}���3mh����PK[lSU~uЂ�fN�aI�7Mwߺ8�ތ_��A��#sf��C�����{;�mC a(V����J�1�Kq���B����-�l��lx����O�FQ��>3�wVV5\�S�F����*5Ɣ��l4y������ ��Þ5��i��e�GC�1�K�~)�s�P�޹�z.�+瀭���J+u����D�2�w&ݲ3��I�8!#�@���E��Y�̐���1t�	�2�\�Qv�מ�+]�ZY�]�Al�����c��*�4������5q��?I�/�)��L~|�0G��".E
�-/-���c��gXr����;���]I<����P=fS���w�Fj�?8i�g
�����ϵu�����-�
���	�Sv�,�rg4�<�����	&y|�-������V���`��+(��m���z-L��{O�`I���Q��u��&3 Ɒ�5�S�\�F�WCV��`Se6M-U���f�[���
�� 7��u�p�F���5��X ,�.��[�s�H������bE�eޒ�m�*A���Gt|a����9k��D�G�~}�?�v�1މ2�.���-7�W��Kt�j�r<�@�YI�c����	�cE��z!�6v����|�%c_�ۃ�xV��c�B�R������=?9"��횥��-k"T��a�N��Z_f^!��C�[��Kն���������?׀ i��A��f��_�K�;���*�Чq�w�D�����d��3���yҥ��y0_�w^��-LZw;6��j7'o�jeڋ�s��;������{4;>8)5��}!�əolo��j�~�@k�@���~�G���Dh#�o�MqJ��\v����S��ǰ3�qZŗ�^��E�O<��-FMc���Z�[OF<���v09���-6�e{�2hT��l�_�Ej�&*`��g/�&�W<;|1���ŗ�hn��/$|[�!b��aR�p$�f\hgHq�F�n7k�tPv$n��+1�ƃ-�av{K[�^���ox��5��h(�(���i���"����rs6�q�o:O�,�Q�2�:u�%K��Н�	�l~Xܶ�x�����wI��#���m��E�d�G�_����:��:�����t�߭͸������V~�;j�w�.2���,(�t~ǭC?��OH�
}�S�l�EP�\I����M��q-\�zC���1�i�[Ƚ7_[\xwM�[��+��hb��HD�!T�T��̶�����*����؍��C�:����y3V��n�sT�H�+\��~`�6:���T���j��O'���}���%�f�E&�l��?^���<����G+�m�ڀvz|�k}�p�6�n�(���+R��ԉvt"G��ķ��V�-��������q'�����v�'���{�9M!x�?:�$5��6��O`|����3��j�#D��vR'e����b��0�|2ļ�L���E��U�t
B�P�W`�dw����ֆ�<S���&{�^�	W��w%ч�G�?� ,��fհ
	n�Wi�yV�E��1l�Q�5ȏ�s=K��5}h�J�����f�s���]�:��YPo�)�ȵ���:�u�:�" ЖiLB��\�'b�����59v��@|�6 ��p��9m"L*���;B��:w�%tFEڠ���.=��R8���DbYT�w��F�3ĶO��=�'�%=��
fms0Wg�K�9��Y��y��
��lX�j���j�e)�ŚBj9����m�{\��=�m��/�=����8^0Wl�wP��2�g��Z������"���ΆR^V����+��tc�>�5�iV2˫7�G";���!��[��k6��D3N#��5���a�˂؇�Ljl�gt��'�}�vᆩ��P�=j�k�J6���6ޞ��-�O�m7���N��F��?��V��Dܸ��i��?ƾ{�1�`Ƃ'՗k^6�&e
��K��}lW�� ���������o���8s��Qq��� MB�h����[���d0/����4��`+�>9�����ϧ�;���Njcd}�ɲ�Ԟ�4��Ն�+��כ��'�G8���=7'�T'�q�b�h��@vr��~%��m��)��G+Zg��9��5�|�W�"�=}�(�>/��sgqrڵ�Im�Ἐ�������$��� ��)� ��'s7��Y���6���`���&瘳q^��,��˳K:���\�o�׉o�*�o��dd�pW���o
�w��9���}�Vz��>��3���%�6<�s`��ۃ�j��}JzF�#�Q��xo*�I�u��̖T_X�=��M���m��rێ`�B���~��D?��mj��c��h���b#Y���y��҂n,�x�#	�KW���T:�����׵�� ˇ@�!^I��l�hJHlG����	�l������Iͤ�G=#����M^�ۈ�]%�� ;t�@Y�g�bb��nB�]|����Ap���f���J�/��L�߫{2
��~ �'�w�U�/Ø�/�QV�2���.���{H���&f��U��3���D`0W��⟓���#k` q�Xg�[�od0�Tr�l+Xi���Q��n��rg�a�F �*:�H���)�2̮�a|a%�/&2#h�`���l�NĘs�����3ݴ�-I�^�"&�a�<4���/&UǑA�@���a�[N���=���he�P2�o��}��3�Nm������s#��es�)��y���kC����0tR��w_A������FQذ�NN�\C��v�\�2hx��wϺdS�q��}�~�mv#=�?^�':^%�wՔ���������>}��4�vf�hМ��{���z�fp,���T�1=���O���(r�iG�AO�w:��u[຿��� �ۻ�����X�0��F�g�	�6��A���&����L�:�g�*㡀��w��-_���Q�y���ۑ�Wr�WnR�~�?b�[k�����@�G%_v;��q�^"��g� �_�s�"{;��S|oB�����S6C||�L5��G�|p��Kyk�[�ݯWo�7��c���T@Kx�Ez�f�27�i��5���p!e�N��:2�Jkگ�Cׁ���G�D}����΁M7
�l&���EвtΧ~nA� Y������oU��l�w�巣؝���#� G�J�"��q3�h�̱���(�@��f@.W������i�P�o}H\�Ϋ�yw�xE\�x���T��i3�ub���(�E����_F$�lԡ���z�X�Q��=����ņ"Ӟ�;��k\	����� V�DpF,>���*��J�����dgŞ��H�&:�N�/(������Ki̕���X����,�*��_k�Ě��<L����Sy����.�GWTPLH$��L�5��	Gy/��1m�m[����Yg�?Z���>�j*g;�i�~�%��{��k/��Wޡ3˽K�Z���&@�2��m[�Ep�æ�`Qd�/P?���c�� �G-�F����>
ǒ�� ��-����Iv����͸S�I���ؤZT?�e�6^�v6Ѭ�	�CQ��Z�J��A%X��u[�I.~�o*`K�:t�&g��ׁM��*���������x��'����>Ȱ�"KP�*�j�:��r��ˮi%������,��3a�/�c�9��Ȳ�ȭ �8G��6�� ��I�γ��m\	ݨ�[.�1<J��g>�u�5�~鋀��Ӆ{�I�������)��~3�H�CUH�N1��Ђ�?_��3�����Ub�?���7j4"�I�/��ϔ��_�dG��SB�<���I�m����a��v�M+�%��M�>&�7ZV�*��lMF4�;�� �3�0&�N���`G��rz/�v�����FK푏c��3�@|�q�D}�TWn�r�B[V�6N|T	0���<M�i���RUg��gA��`7��`���`U�����(�`��_%Z@<�΄�g��K��:�Qq���l?���B1���Y] *2 �+�l`�Ll����0Hy�QU�-��}�X-iS�pӋ�(pĂM����g
i��%��Wn��N�$�'6�]�+zǘY�� ��7��/�(��I���Hs<��:ܹ7��q�4����oRwg���7�@c�n����g��WZ9�����
��{\���'A�7��$EE�n� �v�H�e��n��L�}t->,o%0����^f��5�l=v���A���@n�Y��V�quxR����O�����ޡً�<:��{ԑZ)|��4�d�F��a��м��z����}dO�{K�<�pQ���|\��
F��E��qH���cò ���*����t5|�J��E��[t:o0��w
7ğ�t_9j�����߁�{�Y��멨lM���e-�] U����1|�D��"�-s����(���	e���R�o�o0/a7?)�91�{�*��k6����9H�^&��NuC���H���8�I.��g��<�	���&͗XhS$ԯjA�9������i����\X{d�t����'b<�;>#����<��Yõ����+���6��D�M:X��ϱ�`��gs�zr�� B�]�?p�8�B����m2T.Xq�����z��D��C�o�= ��2<�2�G#T�;v����>(��|m���w@�����$��B��!.�%���]QG�.�(?}
P��=�{��q���uN�,м�ԉM|P䄺���}����p�px��_%��+��/�F�-]Ķ\ɒ�VxF���[[F��a���<�}>`<�M 
 	�.x�+e�� f���l�N	Z��_`m7І�ϒ�%} {����7K<�'.e5IUX����|�����H��z���	�6�:����I@�D�6��å�����t�Y��U�ܜܘ"�]	�4�4��v��850��sp|��w�z�V?^��pl���M �3O���u�x���Ae	D�2��^�
��/CM)�D���t/��X6���S�K(ن/Mc�Dk�ҢFd�#X�0K����4����]�����IU��\����wA������V;�������RD脻�U�N�+銊,Ll�����	5d�,��5�Lױ��� 5>]�}a�-(��=P��/�,�~8Jo�\g镊"��mR����W�X��}��-/��]��..����`u8D>�w�rP���s{��G[��K<=�=[��7Y�b�T��R����Yx��n�=��x�[Em��e���%�'(6�ؽ�lpO�S���G�2bG�h/��v�"��yŝ[6��O@ֹP;�d`�Y��AZGߘ�B�U�����@`-�T&��!���G���8���?ॠ$�=�q�4�4H�y}i�cN���P����G �&˗�YM*Jd���W�`�ܯ6�z��)7�K�����0Ζ��f�W{z}�
~,���1I�4��R��:���Cw���"C����SKk��CS�mt��rb���LWL�X���D���L�rE���~FO�v�W�G�F@=��7ٟ&61j	n��#�t@�COX�1��P|Wlo�J�\�j���%T����>�1���"���B��xL)=z��1����S�'ֈwy��I���n�T7�����9b�^e�с���g�t3N��ܨUc�G]i�P{|4~Z+=�5��<t�)���;5�	r����z�#��%����#����>��}{^6�`��PJ7-�y�������S��������ț0D�gS�{Bba����^�z�w�eM2�y]�sl��/��˘�vF���?1��A�	{�}��p=�?�Ȩ���x����"���۾a���x|BIC��_�5�őg��u��1��\Uվ�8�Z��/�ao�g;���L��iK��$�;PMx7�.����w�������X�� �&I������f�)th�ϦR�E1f[o�v\�ą&��l}x�����)�1��-�	\,vk(~��y^��}M�֏_=��x���&՚��4Q���:KX!���1I�ٙ�R� Mt��3�J��T��0��C�� ~�{�3s�U�'{1�̍%���� ͝��ᖲ������N9 �D��Z�*��la�寇�������x�a�@'��˽ ��u��1�M�(R��*kV�_�gh\-7Wz�=vz0�Y�@���t̘`�E�2f:CD��w���٠!���T����ϚW��^���k��(���옷�ݥ���CA��Pe�I��i�� �#&w��W��E�Bp�f8�aM!u@{%�=J��9�4��<ӏ�=���a�ٗw��^��v�I�8�n?Μ�/�2�-� ��C��	���]�Ñr.b�
��M�q�,�+O\��|(�nH�{����=��Z����L3�N7i�j��&$��y���.�\�w7��w�`js�������c8�'V2��	λ~W�E���d��\��D(��"+��Xs�q������#,Š��'Ld�"�4��h�H���
2�<��A^6x���^W-�F쾖�~����&����(CD��3{'�(����jj�3�}Mh�1~�Ȅ�Şnp\}U��lŘ�ɼ�7=`�h����P �
��+W���MZ<����s��cd�E�*�
E`�Ye�$���5�D/4:nP����4oY�I�<���*�CJ�(����,���{�Q��s_�U��XIl������	�xj�
������8�:�+z`KL���2&n�:�:����3m��$s�z�?�ׄ[D����]__-i#�j{םpiCBZ4	/����jy�^0\�?ܷ��՘�}���X�F+4�miJ����B����4��F�����6wO�f\ߣ�����X�A����@��l5����< W��+�0\���������1����T��;�y�w�zU݄q�w�R�Z�-sEٍ-�>W��l$�B#OjR��:��G�Lď����B2@�{��Y��"S&Q�4y��|7��s��u�8���2>E�L�͆]��3 ����_�,T���1���d���7��/![�;�J��7`���Q#A���J��[��9��m{�V�oCJ�+���3@�T�s��'W<�T��n|l���"��.�]�ZA�bP�P4��*��T�$uA'�W3t�|�>��,�b��e�K!Mņ0U�h�5��3q25�ȦR�q�&v�o\zu�d�v��s y�n@�zb�?0�v�zP�ݪw��!2�G�x���0!��]a�;��0>3���]�;o�bB�j}ځ�e<��
�O�'�7��V�Ξ�����9G����9H��L���m�?ӓ�'	���bg���A�m�E�I2�DO��>T�K��-��5R�j	8aAG�G��_�|�����C���}��x�6☧4	�B�e!՞�,8@����+ed�!<<Kİ�$�
��&�2
�A��z�����%q�x�]S��@�:����x�&��Lޠ����>�fq��Oqz��-���/�^U�Z�Cuܡ8�쮲\R�KU��	Cr��O���Pj�e��V�N��,���<*e:�������X� ��Яe��*�ʔ��8�_S�=ʠ� �!����,���u����jpoq�b� g_�&<X�H�R�,�������qc68"�t��:��xѻ���vGzyЀ�>������]�i����ATA�D(7Wx��J��e���\�ִ�3���.�r�!Xy��<��pY]Mm����dmX�q��w~VC���sk�Z���O-���~��{;�T:��6w��0V��*`�3��=�;�|
��&&q�ܤ
dCҳ+���J(�����B�jp����HuNm@*�=��3���Ғ،�}�O}�v]'��x�@��a /��A��.��(~F�h4#
�A���2{:�<�0C7�(�OP���Պ$��I��l�%+����=�މlي�ʩ�P��Z��h�1y!���H��D�����Q�.+���
s�l,;���s�-�Ӱ���m��1�����:�[2#7�$���ȗ���D�W ��o�p?�L��uE��E�`��YPt����3�o��W�� n�C	�����*�����`�[5 ~%|�k)�h��:/~�cgNR̀:j2M
���;>dP��� wv1�>8�	��Z����yW�
��:���l�  ���f'��	J���`}5����T^I!ecE�������'�\����}Rd��{��9�({���
Ybr}�
�� ����M�wmu�ŗł&�EU[�_�"S�THsO���7��K0W���Eq95�J�bU"��J��h��W)���8U	�������}e8�Q�DD�)J�v")� �"�N��e�([�xu��� ��X�&�{c�nw.0%H(� ͘]|��P�5^��嗈L�M\�FӾ�� �}��$�m��%48�5�&��O�Ö�`�����\�Ϲ�(���N��OQ��c�qLJ�{�е�hS<a���s}Y�(C)���x��7���®��O�.w�Y��z��mcַɚ3�g��FmR!l9V����������Nh��ki%�1)t�S%���W$E��AaY���e�5@@��A��AU�D-�_��Na4�T+��f�=�ؙ�%ދ+y��?t�>�ǰ�5;�)��E�7���w>�F��\�)5E[=�|-7���<��L��^rtKw�SR��E��yi�B"�p���wI�%��eģ9GꚀNy�6D�♮|�}��o9;�!C~z�)�z�Y/����|������ǒe��� ��v�dA��[��e��O�Ma����ie(�nCFHh�KbTiY��B���	��9e��5Lo2��%9�w�=����ԗ���7<*o:� ҡ�lF�E��&����u3X1»V�R-z09.|'F� ������wg�5P�bz1m����xͶ�_q$C/s�#2�S[�nA�5~森��j��,��m��Z�)DT
���Ԓ���~��j9Ź�J�^X��x�fZ��C�����awr�R��ִ���/9�Y��s��w������1�
�9���p��Z���Kr��%����U���>C^*@���W]����9�J/P��z%��1=u���e��j�����{��H^߳�Ί�k��E�W1�	7�2SyirJkzd~���a�hRy�G=�R�A�_�e����2B���	cU`�C\Q�F����3N��N��E��S]�d�2͕�ط/zO��n�Oo�����zi"���ƛ�p�"�С�!K�����h_G��D?>$C�b��=�ќu���{�*�Q��Q7:��E�@�O��RSC�7�,F�^W���Bq������`[\P�Y�Y�rH\�0[@�/�c{���n�u��=n�5����i��P�(�9*qn]fQ���<���ʕm>���8�XlL�(�LIqc��`n�8���!�!^?4Y�;�k�h5X'��ye�����^�Q骋���J���yMȓ�pؐCS��br�zm�
��KG��l���ʢ_���e�O�M,4��G~�25⽵"���ɑ�x[�.�o� ���P~ �l��n�Ƒ�id`�/� "}�l�i�RĐ<M#?0O�P��dec+�Ω�Wb-#�;G%-���ը�����%�VS���n`�ou`ͦW��I��ͼ2�j�o��+�=�än����D���h��g���'\�7�p���|��XXѪ�Z�#��U�y�@O��@-���Y��Q�qm�HF�%�^�记[pA:r�л�2��f������c���n�/(`h��CT�
���qxlZ_P�Jl>&��;�ރ�"	2�?/�s�,.���?@Vd��8�n�=m<f��>n.�V�����G�������\�z�{Q�9�n�g��79s�2QZh�S�6rdQ�H��Z�;r�ݗ�v�E��U�w��?��l�!7�k��Q8��bS��FJ���RX:Vm�D+x8���܁-�!q.�/��ͪ�u�I��Gh~����by�ٓ$ݢ�z��su��e��Q�Y+p���-�`D'N�c4�/+�p�U����:N}+Km�]~�%s�宒�
iRf-j�����T��Q�(���aP�u�9��"��E68�����/�ĚbY̽*��\�v�nW��pǏ�%�ڲ�@�>*��S����>�F�em�T���/�����Ƅt��H6m	�|O��O�g���.����&��[���]���GO9@$�g���!V��xHi�%���jypU������|��Ɛa��s*t�����j�Y�[n>�^U����2I����fD/�xm2�ϸ��n���Km����m����d����z�% �����߶[���֚�]�Y��b��]�K�>�b�&3�����;F�,z�q�D�{�b�BL�1�#E>��n����A �
����q���K��vPC2��NCΦ��PI9]or%p�">�p��R� ��*�ӿ`+%�8��1�t��(=�E��𘈇b�Ǉ���H�+�q0��PƠ�"��~H+�������[�ob	Đ$.���R#�σ��OTH,��<��%$}a&�j��ʘ��2���V�qD=�'Kx+��F���c�Z_Fa�`eV
$*h0s�56y��&�{݈o�?$� (,�6C���*U�ﲅ�a��8�҇���#�%��+F1� V��r�?s��:�eg�8u(�����J�X���0|#�r(�������[Lb1|WBwb�Yh��Cu��8`������o�/:̐�c0�Ӭ��c�3���(��T �NR�-�E���<�vp�1����B�1l����Q���4n�9�Ub�A��ey�vJ�Tވ�:'kf������<l ��KO7mr�{����x�#/�M9Nꎘ7�_���=�v����c��������b��(��'��+9Na�U�;j�E��%��J:{g#���(_�9�W�J�q���l�^+�ѡ��^
S9��Zv�C��P�>¥�ɋ4> (7��iġtG*��r�U��_�}*�-'o���Zvoic��f��+>_;j���L�ܔE��o��|+6��P�(`1'Ļx�m�t%�̙�?]vf��3��^IBx�l�_�9��B�Xz`/�+̅�w'��U��kD��s.�`e�Ջ��Q�,�SUS�8��jN ���U�޿t�����K&����j�6���>�9_����JN�Cl��9�Q��7,���=@���������N%�9m�#F���T?��&�LT�m��u����&|D٫��A�eDr �d�����j���JF��c���*'�B�����+�dۯ�lYa�_6�r��byh\�OY��s������x��~QL;��8����m����Mim��l�j��l�2�ܐ'�C��&�1�lv��%�O�Zj}��w57$��j	�V�<vix��[8� ��F� �&��g��8�Y�d��Q	�yqTѦ��XRɻ��� B �-�B\1;Z_=1�Y�Tm���i�/�`}]S�S��@�ߵ~I��-/��p�)�_(����s�'gL��I"���u��ʊ�'w�+��`�Zԣ~ɸ�ٞX�P��- $7HE���~���{J���Y��+])SΘ���"���xA*r���;��y��\���_o�Q��)��C�|��_��*��������˝�R!��Ta��u�lS�azy�&��=�*�9���ⳳ�v�O���а�pc�_�N��m+�:>;
$N�>��A��K�-���U�)���X��3��ՙ\��R�UӘW]��d a)"6qd�i���[�ֵ��"�Q��K���Jon/�@`'	�Y&	L{����� 1��נ3�"a�O5[���0��6�e�]z�M=�΢V���GITr�o��U��K�/*eE��j(�/I�8�B�-,V"+;����6m��
��r��N��ʚ,p�%�_�i?߽�;�8���=��N�bT�����c9�/��\�vJ-@}^�ق �l�� r;�tdq���"�����w���_u��M�
�n�	x��%�� ���ʎ ��If,�����r�j�k&���>!Gl[�����w=]�y.�az�6����0ν`��f�*oa�_d��q����1Z�X�����S�U ��5��D��C`�a:���U��'?e����蘯��+���8�Ϭ[Y�����Q��B�Ёr�k����}�d�.�V���\e�ڶNȓ'��6i{�}Ľ�Y�-W q/���Yx�O�z�"^8K$�C�W�2���>H}J������r[Q��4���J�D�6q�I{86�?��yK[� �Fa�Įd�z�t�{)��<i���Z ���i\�<~\�u/Q>QM4�����MM���_�~�ڋ���,���f�["Oa#bZY�F�ɸ'�V|�moj�]N;7ߨa�:�`�@N�Hh�g�B!��������1�Λ�ӷ'+B��X��7�$Cz�����2�~��UL���d��Z��zf;:�ui_�wm������N9���Osx� 6B�֪������"E��n�Y�3qdR"[���V�əeܯw/%�L�x��D'�՚J��=y��A��p~^�u�¢�h�ּ�#�Z�,�6t�=ꉴ
߬��)���тO�, �e�W���V���m4�D��cN����č��@Ǿxd0�C�Â:�� �y��)go{;S�F�Z-FLO�#�I��|�ts������@�v}�vȴ�~D-N����>,���)t�t��o_��8�e{1�3>����H$��*;N���Ѫ9���j�V��k��A�@�'δ Nc=O�%�rp�r�׷�fo�����f�L�`�)��I���i"OGt�X1{԰���op%�^������U�e� |*���0�ޒ k��(&�5�&~�OM�8������_Z�>\��	l�RYD�e�׳JZؑ�s�Ȕ�"�ȆN��Z���C�\s^,Ho�l"^�&�1x�����􂊥�1,^o�'�[�Aa�Hxu��dJ�?{G�� ��4=d�n��o� ���/�h�W��L������Y����NW�j��� ��p���ɟ+��4?�Y��c:�o2��Z�I����ӵ�(ħ�g{	Cq�PuK"�*޴d3')�^�,4�h-p�Ċ��x�fGgrS!���Y �#d�'1��T�,����h���Yt�r�p�	��瘲1s�\�� �o�8�<Ȯ��BB��{�`V��n^�_����i^��}�/�l��xq#�x�ʢȈ�H�Tp����H}��68LX�Q�ޖq֠wعA�u:�|��US9���X�
t�_��(��t���i("�9w���<*���8x��q����^�'������_�A�_��m�%�u�R����t2H�poQ�����e��}x�")������(/�`<㍬�����9�j���e7�������y� 依����b_n����r�~؊(�Gmaj5Q�q}EPe�/�#ƍl@WrU�]c����jow��g�S����8+�����i#�!��0ػ�8zI����_\8�6T��$m�m���_}Lv8�NZf�,(;ּ`�0���$�?�/n#��H��Ɗ%��`�C����+	�*{y�.�����K��:���5��k�&Q8�o;i����0�Y���_�PpL��"
��| �N�ª3mF�Ӄݻ�$܊���;v�0(����V��r�$�%��.�ʆ�԰�&��Ȓ`���{J����~���#��-}d���LN|2�S�:Q�qE�P�?g�J��s��%�3g���1J��-�INgH_����s�mɮ�G�x�<�GD0������Jx~�G�L�c\��nq���[���̩(��)Y~�G���*��s�g~�Q��^��Reޭ48&�F���5�1�5[��T�]�;:��UqGe�TeT�WOJ�Sb�I/���ٿ;/3���>�|�����5��PU`p+�}�}�/�h��xp=藙�E?ۯ��L·͈'�MG��05U*�R�lqFj��9E�  �A��[�?�bU��Ե6�	�h���v�});�?�L-��Ƥ��0�X����״��Q�Y�)%�s?y�8�7I�(�P�wq�W6���l��\�g�~2��'�ǣﬞ0�����7�����CQ���'��^6��-A	�"��y�"���y��r��(w� ��-�W��#Dn����z�1l�[	�}	[*V�̌�����D#��UH��38�3S ��	m���.��|ؓ`i`�&�~�Z1���A(w��hYv��^�3��]@�/��e>5� �r��xH�^Re��$�tML�F���ݚ|����N���h-H�	��c c�e�wR�$�W��M7����*%�[�Һ�̎����Vj�2��5ߚS��-�2���z�ꑪwQ���l�֯ں���M2p��j����c�k�Ym�T�!>|��}�E�P�G�L�Vg*�D�L�:<�B���������n��-�������NF�@+R5��ɍ��÷��"8��~�e�:{��Z�6��}/���7�㞢�%"ۥ\T�1��Y1�K�(�����V?�8|��h��BF� �e9���*�E
"8�>�0����a*�8��"[��"^@���� �����ק������D�
h�5�~���2Lأnq��zM�H��z�+^����H$�V9��^U�vT@BT�LGy�ࢅ���5Q����)gM}��/����(�e�R����w��r>G�|�b6��L`�2�^�9�T��!�Q���7��Ɇ�'������M��#tv���J�4ߠ���!a����܌d#و$A�D�p���9+[ 5s}�;hj�/F��&ռ]:`7;ƻ^q~,�v	�j��|�*T�Q䡝C=i���xh�p��4�-�%����!�Y�kzݕ�g�
�&5v�ӭ�zĵ�� +����(s�O5��1"���v��2c�k�v��XE���2��%"{M4{�˹m�?�p�Q�ރ��;��Ug���"Q*���'�+נ�6:�5���U�H�f{��@͙�~���qd)^�%Ů��i5p���d��>�fx��亡Y�5lC��]�@u�S/|�6r��YR�Ffx⥇�/S��z�́邱)c3R
�.
�l�̀K���SO[�z�p9,E�Z�d�5�@�h�u���`����V�<�y̣ϣ���<���h݂fI�3׳x��w>�Z�6��7�-���k 7�u�!:Ve�{��Ved��
�j���[�kL���:��^;��(	s0sc���8��&�gO��?@=�T��<T@7�{�2I'Da<�V���#�G�3�"Y$�#EqÅGS����:����z�貉Vxk���ٯ�OpC�`���ZF�5��AB����n��*A��Ɯ]�^Q�]�����}�����@�?͕���97�ũe�"�L̩Iǽ��������r���A���z�~�ؿ��$�0��Ѿa�-"�?�q���5��x����nR|��2�#��؈�䖌-��/�V��3K�J=(���(T�֬%�Z����d!a�W���&���j�q��TI���d�r��y(S0Ʒ��������O4��Q 3��U�a��KZFW�FR���m� ���;���iqlo��������N6��]�C��>ùx�]Nt�.W�V�{�O7�Od�5L߄��~G�$� �U2�'w��K��q{!(�LШJ�g0B��Q��~�6e�X�s���*$js�T�dU۷\����U2
���2֜ΰ�B�^>�47p!�#ܖ���=��ƪ��A�-h?���{~C�����/kg�����~w����-Z��+zs��i��@��{q�������j<�$��h���[Hk����d�Eo�^m �&��,�W�3�>��,f�?�?b���f��q����2�p�2]�l�!���Ӝ0Y�}"��2�LY�9����W����,�L�� 
��=QE����66&$����~}�4����zy��
��-{T�k��d�h)��,����NT!��^��"���K2���J���C�����9���Bf��3A�>Z�~�%U�_�Y�r���
w�Ta���]D��Գ�3����?Ĺ%��C��O��v���2�J��&8��ݲ��@w�k�Q2����R�~�Xy��I�Ws�ܺ҄��ϑ��	�bU5���.���&��æ ��&χ�K&d5D��s����*�G{�*QN�&��Q��XR�X�oĀ��~t<~l9��ۛ��^�ߞ}����=<�:<�"��]�G����]y���P�%.rNa�����}�-"pL��к��㓒/\Y3}[׭�]�k{��S� ���'��LDd�@�'v*B�U�]��.��=�M��vf)�����:�=;����E|����=��y�Vb�#�����K�.X�`�T�!��P�պ]�D�	���t��R�	t%��$�L���S�Pe�4�nIz�gĶ^Ϋ��4J�|iH����|,�TT��2��`�f~t;��!| ����o�W�?�����rg����7P#Z[G���ڋ���5)��ݼ�� �����+�����H�"�S�ѲЃ5��?^^�PHn�F]��[�Qe֮�I���׃zU��ydy�jv.���vB�Њ���rI�d�|
r�$�X���j�8��B]�ʎ��Fx������1�Q�Zq?�PېU�N��j��2��� ��,�"oM�s��B�*�D$((蹗��E������#�I��(�����x3�j�gêߕ�u{�(��W�8f_%c��!� w1���"q�cT������40�Iۮ���W;z��"Hl-ɣc�rA�⚓1f�Mm�s�J�#$�!�U������R���y���n/]���Ŝ��%���C��>>�ܱܨ��`Q}g
ۉ�l!+nƻQʤO�_3ۅ��Xˠ�<������#�P�A��q�x�f��IcB�HVz#�L��ۉ�kmq��Q��W�ٝ�'�
ٲ��1D8 �lI�/(_��f[2W�i�S���m	�=l����V�]�yB�qۖ������򧧱���7��<�"��p�4I1D*��E?9��}*�"��FhgpǛx�%���a��&�8���U�6�2M���deW�� :~�u-�G��W�����l�f;E�5�<K����}�ۏ`�f������L�����α~,��.�WW	�CĆ;�RxM��1��~GN�,�N.Z�g�U*����m,X:Y���ɥ�]2s�܋X|�m���>��e3'��K��h�\�.vuDyfBeY�ƪ�>��^^HAA��lf�E$9B�� ��P���=�k�8�f�	M��ظ���f{F�R�#v���u1_�5_W�=�8u�գrڂ�������^Vp�,K��;���ڱ�L���W���"c��,W�I8Յ����=��F&�;l��I�ZJ!�f�,u�:[:��{��>D�htEdJ�����]�:���A��H7z��V�G���*L9m��}.��?���7, L����=���ټ<DwwƈB+������*b�DN6��w��r�m_X������A^�	�ɸ|��r^R�_�;�֋�U|}���h(�SՉ���[t2-u�\�uݛ��ϝL�����˰>?}�{C�c0G��4���*6�9�K�q3�%��;�#��vҨ���<-�ɕ�&��qI�?8x1 f@!
�?>F�_�oɟ�ԡ��1�����۔!+GzM�:Gu�v���i�u(�c�eih�>{��b�W�
4��e+��2���!�] ���rHa~ˬ�E��WG=֑s�`��Ҕ�S���r��z$1�˓���7!�(\:��F^�˟*å�9Q���� J�|vo!����*�s�ey��B�N�Vl'��C��n�U�A^,!~D�Y�43��� �� �8>w�����Kp!"udJ���eli�T*�=��8K�#nO)W����p"�T��o�����,�^'x���0���a�y��ݖ'����4	��:e}����f@ElبZ#2�ԯ�������a�>��(]�M�~�L㻄��pD�\h��n�KnR)m:6_'cڰ��$t�����NS�F�Ȼ�9�8.[�06'�$훜��X���-^\�M���_��{�iB���ߙ�g�d�:5vB��lc��jy�M����@����hW��,�؀�W��4W��Ag�\�y�#�����	�ٻ��b�7�NA��w��C�!����M�|9H8�k���M�wy������s^�lhڜ&݀5��@���Ym�Dd;��ڋ1�}��IWg�����������/"�_��x��Z%=RIΝD�N���{��iJ��ɧBa�x�o��l�(L���[�4W�=�X����l-,;=�-�C�r	H�87���MK��Ό�o���D�������!7����>��1��s�i��F�'����W9�K�Lb��j���Yi,H���Q]f�H�Z�³̴�2�Ќ��E���J������O�Krő��I]�-�^�b��f�y��%�xوmp�F�l|�S4��4��&<��_~G3��)]�I�(Cq��	��{[�ˮoy^4��k�7���R��Td�P�vM7�A�5���C�+�g*i���y��
�[��.��$kb���p�W-@9�3��y��)��xj4Bu��^S۟���8��E�;�V��G�Z�W'j��l�n`�Y،X�<Ar>^o�L�B�Q�QD-亱����Tz��lT�~�K���Kr.o���U$��:��I�Y����&9���:`��r��`�?u�}LuB�_ǔ�Ϯ�c;G=�si����{8��n�Ȱ�Wkú�Ukh�L�^+p�n�l�5�>���A�Y�Hh�א�#�v���r�w�����)�V7;.������A� W!�SC~�j6f�H���������LF���1:�1���<����D�,1FS�*�Gj����bg�a��D�FKk�����q}q��cA]kpIj�E�����M�m@��Q�ZU�x�,�5!�	U/I n�[�6������9��ƙ���0%�v	�%h\x��P����
V3h��I�!��^�6%fd#���~�!�k-i�,(��S?I�%��3�mo�7�(��g���.b���M1O��O,�ț�c�Dz�Ov�d��;��(s�̂�p�,�����?]A�7,��56��w�*)#
������\8���;�.�G�e�B�E=Q�L&KЮ�5��h�*P�CD����#G)ϜB�GJ���nB�����IД۟���vO
���?��_jYh�%���)5�ka�l[����j��m����|�/
��"�36� d��+��U�S�x��(}TV�/-i�?XX���K�!<�	��s��c��ɫ��fI��q�3��y)~A)�m͆��u(���gf��5�a⿼�,�ZWSJ�a�1EZ�˙�B� ����3T�a�_{��h��I%B�����L	�����9�L}N�]��Ѣ(�ǀ�J�;��� ���� }=LT��׭V�7>e
�J�tK�޹AZ�cI��x��=>�5�5lOX�����y0<�X��r��0�u�^�v���� �QgeC����gCh�WS^
N覀� �xDþr�й8�ӑ�>�%� zIӂ�]���`��]T�f�ަ��V�,��	hi\�1��mf�Ɛ�2l>�˭|Fݨ��/��ӽӛ8k^LG��==����B1y,�1���锺���7}}���#Ɓe-X �1ZFkbL�R�W'�J�*��5p���
r�.Hg"��d�q}Yj�
��B,��_��e+�v(A曙���]����,�s1T��r�Ս��_L��ǉ��*��r�
�Ȗ�	��c`������2̣�$�Z��;!W���������}��І����t����Y�6pߍ�a����锊�<jk7!���cXǲ���;�yR� -��3�	2/� ���w�6ɪj$������A����S[7�w��Wk���&q/�	��)|���4*%�'"�����.�$��5W�b檍�Z*y���3@upٝ�P�)
����~���%~ITs��o�\��Q�Z��z��������?�@6I��ۨA�l�N����Ӝ�˵�6dNe��H�l^^C]����\O��w�}O�%����^�����8��1��P�4'_��F���H�����%�ȚQ�����_)%�o��K�H@�*��W|��Q�F��R"�׌_j\`�٫�<�*@\˝#7<��i�W���_���?X��]$y��AJ<����Quד��P��|�9�[#5� Ҟ�]���޲T۶l@
V�v�scR��(bS��P�moOϟ�����k��@pa���.�m�����`�]tg��CU�J/�ْ�)�9��C����81,P r���#�i�=�Eov�1p][�"mÂr�3��F��yH�٨�?Y���j�D�`���{�z�}��r)��]Va�ܟ���+zx�?R�7tX�c�6�ho$�My+�+�����Q�-@��-Z�mF��`kM�~K� k�`:n�[>9�}����=H�D�����
��I>f�8�R�E���E�}��q�a��e��)ļOc)N͐'�1<sl�m�.�G��Ϟ��=+*\/9��y�.&~����*�:^�Mlmu�Ȩ��Vk-�Ч=�c��RG��tT�V�þD~��rVYo�d�|K�
B]؆G懭�����_I��������R�+�	Ś��eiP��	%9�7]%�!pX�V$'�j
���i�o}NdPzB�Bb2�G��=�QP�qB`H _=�dK�XIb�q��?@���~NjY��UkMQ=/���;�~1�N���M׵�Nx��/"�ǭ���1�IJl��E�K�M�k��L�Ǧ�}_��?����Ȗ����\gt��z�_:�Ik���ܢՌX;�5#W飴��5d�6��\c����'C?f3��s
l��@�D��:2�����mŤG��sW�dd	���d���wU�-����?
U�),_�=�;K���o�f��q�!&��m���L��u9"�_��'�>t�(\ʷ���n���QαC�!D��0z��ct3%�CB6��eV���������߆�s��[
�9�1��A�}%OƐ����y�;���AJk/��j��{]{Y� -��{ڋ� ��y���nq�o%Spr0���3�M	�]�ҍDϜH��N�[���ZJ�~���b<�Àsh]�w�I���՞��u�8��k�=�~���ݳ����	z��_h���0���;��l~�,g��c�������K��煋��O҅V�ܼ}�B��$ʶ�����y�q�~E�,mdt_nECg�yRtT���e�o��cOhH��%������WE��:a6/9~�9�;t� 5�8�_Vs��V������M�#���DdC2H�ɠh�8�G]�� ��z{�w��jA������o*�:������)�_����hL�&�G��egfO�j;f��4//dd�:T��p.[;����G�Lv��=�m�Ϲ���"u��:��c�?.V٫xO�J?9!�6� 9J��e	�5��W�膑0�<Y��%S�2tG�G��N,S�r�;9j~���q������nm��K	D��T�pg���`�0Y.��_�� �s�#������a�v�^2���-}t��jv�b��K�ʺ��k2�6Ho1):�;����-�?�pE��J��_��^�.�9�4/�_bI���s�_bD��>��r|��U�Z�s��������M��-���� j���ء�b9�҇��;.!�׳�iʵ��zF��ؾ"�I���r!��D��=;0?��j0*X<S�B?��>Wܧ�ϳ���ǀ ��h�{p���������1lC JQ�APR��\��\w����V2|?���3t�Z�1*���}��o��6�b@� ��y�o��g�	؟-إ�T�A� �ڒ���S2
�'є"��c���D�������Q�w��s.�|���
wڜ�f�3���7 k�h����^�=g���-��α?�҃�� ���Q�K�D���"𶜋4v�ZM�`���<�������i�Ì~�Dta�<Um�Rs��5���&�w�̕�Ѭ}�4��(�������h���#�.�>O�ִ���1���|�%Ta(�#�!����� �<�6�����┄r4��.���~�}X6�D���0U�fB�ſ+�΄nh��#�~�1?3�.�^ҁ{2����Ѭ���G�JA*�����"���%Z[b� �:������])��I��L����zํ���ir�u�kH���	���?��{%���hK�X���%"L�X\1��>��kL7��K�,^6�P�� �f���9C�+���?�xA󁗂�_�Eb�Sq�o-{-!�u�6� �d�Xl�4���sG�$ה��P�!@i� 0uO��Wz��M�S�	����]�: �ϝ�z6�Bu=�{�Qn�J�گ���/^�*�(���cjq����xy`��k�`;�'���x�vc՞+� e�������.]�$yZ9��q�T1�@�arK�9��R=ն����8F��cy
���Ѡ~�_Z	q/��r��k�sP0�q���/��Bwg�^�@�ۄ��N]i���N��p0�1V�g��I�mr�"~��/kBG�֯zS���݋�]��?P�
ۨi�K��M6\m�TA"��c{�� +�F5q7sY�fSv�
'�mT�k����]f����?���K@�'͔�\7��6i)�-��a�k�E�{�oA��Q<RZΫ2�Q�~���+��r:l�|b���d�Z���ƞ%�%��H?',[Cdɾ0��Lū�;�z󯚾'glɲ�}���C���i�;����(g�{��UN'�����a��(��7�ب=Q����Ag�����tk�/`� ȼ�	U傺���T���Vn��kx�Ϗ�'s���3y����{��_��u�w(mC�,AZ�"�����Z��X7E ���|�u�[���[ ���T 6 V-�|����Ǫ1�3y&I��K	Ӭj��|��a�<��pee��@AOva^Ш�߉X�>G�N$�K��9�0���U�߂C ��YHZ~��HTH�����W;���Φz����kaau����ʹ��B��u~��$D��0f�H�'H��J�j��N�g����_����v�0��ҋ�b]���	�ҏdJv�" N���
TK,:��nw�	W��Wo�`UA�;� ��D��ˁ(��R37ނ��?��xw�&H��0�t8�o�4�����criŃ��E�D� W1#�-�lt~B��jpn��Kb�o����Mi���	]�x�~B6>�I:�5�㇭���1���tI�C��'Ӌ'�s�O�tu��SE�ꪜc��PY��Au �Y*e_	�Q-ND����w{G��q�7�A�[]Ɩҹ&���IWm׃2�z�W���XSw�Oh����[��7Ӫ��r�����6���<?���i+߿�V��i���ei%��8�O$�^�!s����� }�a�r�ྌ�g���oXڒC��%)/���P��R�����]�.���	��y�x#1�\{p�>�/y��)M´��,�Z����mX�2)�1�m��Q�\.,�rا
)�1w7�Q�z��F��B���?�<&\)^�eO�/��L������k��l_��׼�U��Ǝ���傑���q����5Q�p����)�](��Nԍ��B��Қ���_�1�!of�&��n2,�FD��~��<�x[F����z�}�j�D+|07�zz�TB HY_�h��
I�!"����m*�4o%��B�$i���o�r>�-TUuy��L�F��Q��>XO
�'p�l�M��vsY� �zso5�hb�+�����9(G��{��)Ҷ\�I��O\E���C�:x�t�#��|_ߧ���}�`~&ݜxՎB��*4Ƙ��8����y�o �������HO��V�QD�$@�H��x�Z<�b��e����8�H1� ����D�E*��{�����~c#�����r>�hX�2�������_B�{��n��T��TM�Үc���x��h+X�s��Ɣ\Yo��[ՠ�H)���K� v��C�n��D���M\@k���S�O�&�-Qq-��!m}'<���c�P!�ГpʽZ%�i/S���n���L���n7�;�۫�l�d��>vm�
2����"gOp���zp����u��"�X0<z?��@�W�
A�@�Ԇ���J��m�z�b����������qr�R���}d��|��|����6CX����Ί����<Ov��^!��L��	z [��o1�Z�L�hC|�P�D<il�<f����}����ęw�k++}^?�'P`�x�m�����eBw�k���zjR�a�X�;���!M0��o���݅O8x�1��T��=�I��DU���&(�ek��42��Ο�M��[�c�^����9՚��"�{/l�"a�{����$�Z ��]:B)�E��T0�ݙ�
�+O��p'55H=��>�q����6�D�@n<?�{��u]��l��@�ۗ�X����k%��,R�Z¿n�����&Ӻxb�^4<����2���+襤�q���Zk}?JO5#��5�t���C|I��J�dp�J����oA{��:R�/}\��_2�)W�i`O��bB�Hq�+)�ʓ����������p�,�љL.`��PZHo�5�����#ݨO�	#� ����Y\r�Mf�p��\�OQ:���IaK�BRm1��vL"�98Q���c�� ӟq��^��e<�q
��g���H���*���*:'U��Aa��|\���q�oiCU�O�]\��m�z�X�Y�	W�ePb�B��~�?Z��ĐF�Ɖyr�87{8w;!@?_���j��.��B$ĮI���Ug�>���:�U��՚	�<�	1�5qH.'������Zxh,�A�,��.��C��F~�n��N�#��}����rN�W�Ò0���sr����x �f��?z�ιہc��uj�lW�N���%`;iz�� ��:dX�0y�A��x��O�^�;J���D��|�5�8����i�~w5J��J���'�ԃEم;��'<�
��M��Y������t�6[�eusQ6�WLM�J�f��(ۓq����il�����76e#�<�TlFC!�S��I�:kp��� ��<%��h�P�7�I�qUAsPFc�����Μ�)AT6�ue�!�K�\0��?i�u4��.]���q.a�<�s¦�]x�ꤙ^D�h���5_i'|5�ԩ�(����W��l �x��Ñ���@�1)��Z6����L��h�@�M���g������׏YtN���������&��xJ�M}Jb���A��B;d�T���x�Nf��9��x�Ɲ�v�L�u���K,�T93/ٱj�:2.Q��^8#H���b��������[�di�~�ӟ��nЖ�2w3�3�R��'.��E�t�]Q����oQd`�;�.ح^�.R��\�	�6�����{�7KS�V=�����2$1ߟ?�2���@�5[���X~��]Ǥܴ�Ӯ#�/��F\�d�o�+S��/l����E8�'z=�CFf���9�[�ٿ�z�B��]$�`����\���B���(B��6F� bC�*4�������>���*��Ew��
��@�A5rfmE�njx_y�b�+����k8�e�Lz��J͒���y �Κʦpg�s^Ĉ{���+{,4�x��i~��,X��=�"�v���P�B��Aba����������j��
����^J-�}N�v|��(��|/,.�^�Kf�X)���J\�Ft��h��뫵6a��5��;rS�T�X��	@��".�zg�_t@�n�~s{�1v�vz��[��⳶8��Qq=����Q���ҙ�u� #X#��EQ�$
}o����R`$��GHpH)��`�J��'i��J8�I��pZ��˖�@�G��?�p��p[��*�
��e���W��W��n���{NN�OH�$r���1���$F�K�>:U��q~����N��Z$/��A��wmtB0,�T�k��1T��zk=�{��� H�Z�=�6[�{�t�J���)�--�U*�ǤĦ�x�QRR�êum5��п�����@���ߵ{�R�Bv�HPj���W,���(������vlˏ��>��GڟQ� \�*]����G��r�0n�LF!�ݵ<��������&:��o���`K7���XJh˝d�k�0��:�ޜ&J?�ziY���ж�-l����[n���p�iQv�Ycv�pظ�;�)�$ ���5w��#��=K�&�4��M�P���O�^�����>���%��-�{��ί.^�_����m~[�}����v�m�L}w�e� X����nZ8ں ����vL؇�_;1D�ڒ,6��=��G�����lE�D��z����Vm>3<�(���E�J�b������Ι������5]F�nT��s�w嫏�UL:�H��{�'�Q)�����5�k��xnix`�x$wF�O�������o�:UE�f�2Rn?a���r�Nx.��-璦^TW���$���SC��(5.���|�v���꿵TJ+�<��x����M���Ũk�]`US%��r2'� Ym��--��vq�hy2J�pݥ��;��NE��q����sg��b���9��+_��~j�2�H�˹�	p;������Bb�cYb��b��*��;7B��IC�B.H?k�d�M =�g����U�{ټw�����P� "Ț���
�$ͺ+10e�<�6��$+�.���m��y%��^D���]쮤g��E��N<@h���XGMl��l���2G��{�0B;k$���?�p�"�,wYX�`;~�`��Z'������=�)����Sѱ%��ö�a��ɶ]r��Rd��ԯ���Uk^ۑfU�]����J�R֐�;�]�ifgzY[ �_8k����Hb緱՘������p|జ�����]���A�'�L�6��D�b;��T���s�7)u�:��?[+x1�ʖJ뽺�r����Ԉ���<kR�F����}�uz-;��vϋ85��~;���kߚ�{��c�K�`����e&�&�*�vC�����5���v	`I���9�y2�L_���*`����F�?ބ�����{DC��"��拺�&?Cv7vk-���c�����N=��\�b�R=0��1(v�.����� �&a��e��|��>~�qV�2�gӈ�bQr�2�l ���j�9�~W>�ɟ8घ�$���F:�>'����2E�+�����4��Ez������7ߎ��j�!�d���J��6^��+��|��F�W&�S#B�t��Y�� ]��U�(8��d���gH߰�?��!#��L��]i�:��)��k�^�ד�A�� )��S#���H�g3���h��k�`cX�,��:K�w Ӂ��`�ع�����u�F���,����\7".��E����C�띨��ը�u��=������毚냵]��81����� o�y��+`���S�f_�nQ���B��f�v��AL��(;�{Kb��+j�m�!�m.	�C�b]��:���.�Q�{ ���2�A����d�If��<�MLV�����p����pf`���D��γ�_�qVJ���L���@ p[���fG�"g$����	1���ޚp��~����j����w^}����� ���X(�������:(34f�k��B��F�+I�����T���ug��V�JU؛��Ca��ȓ��S���������ӱ�g�^�q�I�YM���k���G�6 �i�3�&CH�����x�	[U'�'7��k�4U�l�p��'����= ��	 ��k�l%&]N�ҿ�o<Z�^{�2v���j���ZE7�*v�>u�*�c�l�N�*��?�H�R�����a=����@��^�q0J�@�����N{����}����g��!�jz�e���V�rZVݍ#?ᱏ
�c )�%/��A��h���7�Z�x<#~P"}P��yx�D��|y�����-�A/\��rl��F`�cOS#���S��7�J�m��ͽ�#����ڃ�;l�گ���v�S�t	���t���:5P����zZ�ݘ�dB�霔`r���ڼ�	���]�ѝY�L.�H�P⫬����ݟ�d�3ְ	/}1y.Wë�F����V�֢���X��o:z�,Tu��� mD'�2�d��W�Ac%��@f��	@o�"�i�y����eZFM̒�P�+�)6��t�;Rǫڵ�&՝%�$�Ey����%yj��Ϫ�ɟm���9��������]q4��3\g�`Htc�W���߬^u �ma�dTpu�	�3�Ccu�k���)����:�
���#_�3�t�߷��W����3*Nd��w�������I����w������������A5�
J���( ���8�r�hy�\걝�Mƃ2�d�m�S���������I��e֭�AoWo��x�\%�u��L���wf^�4%7�x�#nW�6xH��.�Y+%\ŖǪ��烶r/���$�A-�� 5��7��$ ���Ή�p�����*�,�bD\H����'`��Xq��Yifx��_�j�����tǚ�:��(at}x_�z����TLtf?R��M�ѫs��7�AZ~P6F�m>��6C ���5�CiyG�v���*��=\er�q\fT��@��~��ڿ�{�0��°�)��c/Z.����^��w�.�gr�-}a�pl1��i��5eb�kx�����-��̹���s�|��,�o��RK��m�K�<Wrh��!����]N'�'�w�>*N�V`<�ґfj���$<L!��: qO��j0�5���n�ʏ�������+����<�7-�W�#����i�Z�S�2^9r�i�f��PFš�Y�l{�� �X��E�}DRI�'D�&"�Z�n�	�d�f'8��'޺��N��xV$�j�Jm�
����B<u/ζ�"���=��"<y�*�#a��_Ϫ1�9���~�������0	N��[/k�O�!��_�b��ƱK{JI��>e�]SL�q����!}�f>�^x�2�Hp��Vw`��7(V������!P������t��_���W�=�}��t�����~�����f�⒓&�jT.�7ؘ�X�UsM5-��K'~�|b���z�--����^��|f�?N<�)����Ϸ.U��8��F�ZGl�y��m�V�.E�ju)���48n�?=���F�0�Sq)=�� ���FS����C��+N��t�@���C��f�J��ێ*��n��������*x&�ߔ�*r���:r�ή��lB�]w-~�Dp��_@ ����Z2�kMh(|���}X�n�r��9+_~O�L�Z+�� ��n�����Q�5x��D}麭w���n�5�j�r c �I}nJ�D�qX�-c?�s�����¤݁�e���H�V[��RK�N�Q�.��vNе�3f�c����WWވ�6m{֧Vԉ���/����D�7i��!z��Sm6�|��/`t8ZN�6�������a���/D�y���g�"W��S��I?c��ZÒ�tc֜Ʀ�]���h�4#�gS	�.`K?3ۓ��/��Y�I���5~?��oX�N"?��$���r�)���MB�J��v��͠b>Wƀ�>\��q�Ġ�1G"��M�]�ղ�*�\֛�'�ćp�����Û�x�����,���*4K�$�s�dH����e�͍ټ����&�������K&�Y	|EyQ|��O�G��u�`����rw�� ����z���͒@tYW/ǉ���DcA��)�r���X���ll��pΖG��(yTZ�8LU�f�Ex��v ����V\}L^�"0�h
</�./6���Ya`��N:-L�=[u��z"
��!�O]#�۵:�\>����?!:98R$�����{�~�y&�)V�6c}�6{�Z���垗�s\S�'��S��B�`�1�D� %ɯ{M��(
k�U�S[6��1�tɪ�Bi6�&Q4�Sc3b��,�&s��dv�.o2�cp��N�L9�܆�)\H�Jv� Fvj��Pn������i�^B��bi����B$ļ��
�A��2��S�)F��_]`:���9���<�E8�ò#%v���Oэ���Ԗ\�̻�yj�_a�]�5L�[ԥ����'P��s���\�~��֞7�N@�_"I$ JfU�`�m�I=�4�<�t��{�gm�����XoeԷx>�
2j
�U],�U�TF<]P�T��[@u��C:>B2>�����Aw��ʣ'���ݬO�vá���P��"ߗA���2��axPj��5��������-!������Aw�iռߌ�K������L��^	���J���z���?9�x�0V�
�*�[�-�'������1inX/l�f���O�
.�C>�L�ݱ^(�^�*:���(��uu&c.�q��I�N�\�d��KК­kf[����ҟ� b�$^3)�e$~�yt�6G�d�%T"Ԓ7�L9�x��tӽ��Y��V���^�MB3�0�i����*,�����A��E�Vwcql΍�䒸<C���V��7�]�B"1��0]����`c��Lg%��.�5��Td����∥�Us+0��Q݆�
�#P`{�w6��7�3Qޒ:�̻�n�Gvb�1f�Xbr���q�	\S��_:(ʎ`Ƃ�Ņ��~lO=c�e'IAȍ��.pp�`��v��8����E_��D�pl�'0�쥻�&}��d�>��YM���D	����b�5���o�33yZ0�m���E��;���u5����W�q���e��Ղ%.���W�{W�aE��b��\k�١u�c5�_�O�F����0L_���
�a��8S~ck���l_�[߶dw�Ra������Ǔ3$ 38�Y�.�KlG���Z�r���-�K��0��ő�wj��|8��H��K�w�J_�TZ����_��o`Q�^��3q�/e7��H�����l���Zy�����:��8ē�|�m��72�h`�������R�����8���Z$��-֢Y=�;*�;a��P)�t�V	I�����J:v�>\�һ4����I�f�o�a1�ʻk�pL˫�D)a���ː��w�\H�l��1� o�#�:��r�?Kd_�P �r�@{/渋J��)j�\�X!8�yVpFRۗJ�=(s@c�s3$@�Ԍ�O[�Hٴ��������T�vT�{6��Ph�9.���j�9����Zj�)~�BK��<�T*�;�A�wB���L��e���{9k�*��5�+԰,�#�Mq����'�}^t�Cʮ�3�L-�����{B���*�!���"�:�*�!�\< ��D�d*fa�[:���`���/�Z
$��e��MI>��zd{�[�~��E��-"��D:�Oυ������!��_r���5Vz��YN��N1�f�R s͹�f�oG�v�o��F�'9*�{`v
l�a-]�S��R�S�|?O�i�״����)�:lU�*�wr#�k2�ږOD�o9���� ���o���F���n],���N8��3��k��N����?�@�fZ��ms �C��T׃�<��ލ���wVK���N%c�P�Ym�R$��/�doJ��l:�WzY���Y;i_��[�(���p��,՞���{�94��|$��3����~�A5
)	ӷ؝\{��5�<f���˞��<X�Q$e�ũ�0�+�{�W<#��e���w�쥆f��x;��k�k�+>	�MVf��K�H�}8�9�����w�W�2�rG�@B�7�b��:�*�B��ge><����D��̓
�p���R���l�K���}1����8�i+V۹-l
��ƦP��O�o,��_{YF�D�:Gjr��j�Cp���L$(N��MJ1�ϓi���I����y�ɒ���y$�u_�؎Ac���8}�i�mlLo��s���1)�q^ҽ@���2&72�\xEx��$��7� t��Fd����&͊�<
蜝y�-;��G0�28�=�.�h!���o��Z.6h��{Q_�a���I4�K�Baa9ܵ�A]3�t.u�®-����ƿ���s�ye�IFW����]��i��J"�~G����b^�?&kIl�P�Γ�V�K�*�b�[��)��3�8 �a(�B�d�yʛ�4ea�d�EP��e����?�$I&�	P%@�����{����u�F��O?�`�8���a+\nA��C�~�
$JO*����b�H����>�7�G��q����?�r3<z���w�&t*�=X!L�p�ѫM�mO��O�Q�d�P��IB��3��!����]N�4�u�}�h�4��;*�'��߸+! 4hإ�GF�]��Cg�QT�E�Ҝ�i�P�l�'y�X<�+��\b�P����~4=��1����5_qºu��+7/�ܻ
A�|�J�阓i�C�o��{��g�
A��焽��<)�3o���=*c�n�N�ӡ�z�y�����wq~��T|~��6��n?����_Wf^��ω�z	ќ4���i�z��B�yS�FQh���p,��d���?g�����:,^T��_�{Z�׵�t���:���br��!�����Nao3�t������
f�>��/_7����OZ��|���$���5oIς��B��M�=���3�q��K���Qe�0(���ʭJ�)�T���l�����M��.n[h�TI�v��M���0���nqC���x��y�D:�}���>_�Y�8]@�t�gN�9��v�'1t?�}�JtYL��Nඕ�2�w1N��?�Lu<�oe�0򵥎��}�i]�
	/�W$;��OX}� g�d�sAr\Ɖ�B�=�#2��Jf��d�l��M�qǜ�_\�>8�2xo�]j!O��~������1��(8ы�� h#�������X��U?�R��N�Yq��?�e)np
�T�Tad`i���2���r^�K.eUk�?�ʻ�)Wr�Dx�C�<�ƀ_�O�}�!*�g:OJN�Y!����$���M��~�e�S'��_���LC��*��:"�d�Ԑ����d�>_ ���/c(<i�ӊP��p�, �}�'�6J�]�,��5&�� ����yoO2����|�*68��H��J%t�Q7u�#Mt?@�����nO]��I��i�$4?�ʎ1��=��>�.؆�����)��[�Ӗ����^A�
��p��7���ݣ)�
p��$�k���L�^�'��!���ֈ5 �ZuE+ҟ���b%."����Dzv�T[�"�A:���t*N۴�_$��*B��n�b�, �m�n:7+��&SJ!J��7B�Ҩ�C�AH;��;s�6f�?(�M+���#�Q�`�<Z,-�Txz�*���8�+)ݱ�>�%ɠQE:�Y!��4~ �4v�˻���HbIz���(@ȶA�(k-�ڟ�)�׽�J@:lգk�����K^!%���4n9��z�ˌ8q䕾�
d�0ov��I��}�'4�К��r�������.��̍1�q�I�pT|	��d`G��%�ZB�M���2���Mj2Uz��X����j��"2�e���9��hIAk��w���l̜�������4v�Ӊ�&��i�iHWm%���p�>���ù�W��s==׎�N�qd �����wa�Fc)�N;ar��s��h�!�ϯ�!��<�fۚ���?f��'r��O�e�l��~L:'D�"��W���̠�f��N��a݇�a�ƙ�U}����l�al��'�dD�Cn�%��&y�B�D]�'��ȃ��;oN��*���F�< �m�@	uh]~��h8&�T.���8C�����AB��$���|Sd��:�A��*��}[��n�}���Ob��G�2m%{<�C�Q��b|HV�`����{�L-m8ə�}��-�w4�}�S=1��CHM�.�:���|�n#���W=��ۻ;��|�0N�힐r���tI@�kv_��7�[Z����F��9|����%U��Y};>���Ǆ�͓�W�MI?R�W\*�K�{b�:5qe,]�>LR�eL���&�Q�� E�(3/
F�{�۵�G)U�A������J*Cp���6��
7��Y�%��=J	���^?����*~���v*�L���y#����)���e=#�T���O�����*��w���­$y3v
Gz+��ә��ܲ-}�;��jm��fW���l�ϕm!�y��N��W��h�ˈ���T,O�q��������:�k
z�u�H+p�:^�fS� 3�aw�o(mS�/锼����٘��񿔄X�dcs�7���e�/j��h@�kb�m<Ăpw�X�Ζ�Ӟ|�.c����y��<�Q�oza^Ϛ��%:DT<
ME9�Y�M�ͨ�U)���Ш�_����9<���D}�x��+��Qx�Ǖռ���Ձ_���c��pi�@4<��$ײ�+�r�t��#�(�E$D[T�y�*��=�l#�����T��z�-������(���J��Q�'�,�m��9Ad���=_��1�p�����?�${�Q�+�v�3��� T��Z-����\r�
>���N��I��`n��}fP>��/Pp�M��`Q��A*R���BE�+؆�����S�2?0�X`�"����u��.˾9W���eg�F�X���|7Cv7]�������D�v�m�|��ڦ���&Q�&�c��~�R�SHXG�>��3~��JҒ��&�Z<O�����0c��B�����i�y��+��]�&H�m��C���i���-���#���/Џ��Ln�A�u͎�/^1ҩX� FZ�55��t��$���{������ �w�$a��f��~�#{���E� �ELR糵��R��Z���R�6R�����>�pZ�@"�x�ǣ�����g���5�`}a��}��J^�WiE�.`>����B�%����D�4O�:>8@_j�G��[a���|�&�vX9��{���u��z;���<)x��9�?��o�A�l��.�G�]��]fx�9�eə�{汣ӧ���J������^��ѩ���ջf¸�Nzc��M�ә̎Zs��}�̝y��ؠ|`s��;y�y��K�n�a�R �^�aG�H�y���YH��+���7�������\3`Z&��S���B��/��[ҊV��SN�+��bSkd ���*2�w&G���HxZ���A�Y9Vȣ,���4=$2D����+bC*���.��VZ%����;�=�vCz�5Ԓ5>F$>��K�˕��|n��`�A����7Q�3k�r$ʂ���o��	���c�v�N[�m���q@�F�悢��g�J����,v�e|*�x������u�kz妫�8�1TɅB���-�N������.�(9���|n��ě&����#�)6�
 �M��4�Й��O�6=O?�١R-r�ؿ�5|X�~S��=��X��C(FC���e�ǛJ�ڳP�5w�"�PQ]�&����L/���uM�x$�zQ1����uҊ����~<֟��4�S�C�X�����qL|����x@jcㄊ ����a����?T�*Ak�^����W�Ȑ[I ���nC)%ƵP�ѻa����Г�im6���R� Č���
�Pw���f�U��s���y{���1c'�Ľ�����T�=�u!���۲���Va/�3��9B"!�iFW�p�C��e��t�.z��򾖍�Ƃ'�F�j�����B�3BJmA2P?����T�x�U�=��j��|�|=dһV��kƂl��'Q��Ji���*X���Y+���F`�]	�Cc&�R[U�톥yP2J�;�ܯ���ML��~�%�(铳���1����� ��׿yA�Ko�I��P��}bqmX��Z��K=��Y�ni�����"{poH�e&�d��Iҁ��Ȩ�)�r2^�oM-u!	*�ʹ �������=�-���$�G����8�E�<�m�ɠ��Cˈ��y�U��"z�9/�[��&�I >X�M�,���(�_=wWZJ���5j�6�X2�[�a-�s0�:�U��儠�����6�]n�9+�VJ���+�1�����Z�
a�ݨ4rB��݉M��|eWL_�����3�P}Y�ʄ�ԥ�(w�C��N�l�nҊ�n���'*W���h�ͼS)�[X��T��"��i+�;3��FWZ�	(��̍����G�g���nPT�Y���b��_��j*�P'ӗ�-t�s,�Ö�5���>�bu���Nh٧�/�pR���-IW�}�V�fZ�(����ݽ�eԏ)��T�`�,�|�F�-�v�j�#�Q�;�L�pd���/~���nC~̭���т[�2�����0���3u�c�f��Z�hlm�� fh�����`h��٬��"�_X�[�����%�.�xIWiGZR�I��y���	�S�ejHPֺ�T���~%j۩�oU������
�d�ͷR���V&��C���hѾ�� ����%��7�h��@�Vn2i����̀C>�NQX��4���]��JGC�B�:ukg0�� ��(�4Ƅ���{��6k�Fl�u<39��;=��x�����Vؘ�-;'"�o��M��$;�%�`��n��=L�濽�ok�v��7C�{���9T������EHA-�PQjV���@�ĝ�����E�ü�{8}Q������D@�>�E�����k��Tt]yA������؅�#c1��W�:Q��4��%~�,U� 6����M�K�9ܢ~�1�Jxf�/R�_$�����{�e�͸���pQf��C&!��ˤ�ʕ۱��ߑ�#�b9��VdvD䕥��Wd��!��(�Q������[�܅7l_��L��7qu�i��px�Q�}��;����GP��aM֨���G$Ð��XE�`�&�^��$�+wj�c�)y�u�3WV�b\���9���F8��I��N�BA�F�9.�LK�w�i��<�$���(bC��"�oŉ��[��Po����`�WҺ���Ў,�Ǥ���=�آ�i��*&��j�}z���w5�h=�F8�z��}���Y���S��Pl��&c3��!����
��A?L���+|h��n��n��Ѧu�m��U%P�Gr��d�A�>�wmm,Nv�����jN|�����'����/V��;��d�J��@z[s�?����	)ɕ%e��������x�׿ٸ�Τ�켾��F�F�䡲����t��_���nO]��P0�S�
z���?��-LN@�;N��=3�q7�'<�v��4'����U�o ���T�'�t7�b�� �:@��x�9�u��
�"�M�7
�5���L,��V/�l�r-X��uD�W�ն�ݴA*c��]^
r���\-
e,xNz�%,\�k��5d�ּL+<�;s�+$p�l�$�ݳ޵&9q�h�k�kcd��KP"�u��"���3H�`��n󖲒�������ߪ;�)V�ٴ�ﺆ�>m-��O�,�n%�[���H�iͱ���K�4�\L��?�8h��l�p������>���ʐ���8'��}<!'�ff1�%YI�PG+��S�ɟc�<��[l�St��χ��4 dlO��e�����y�1V��^�,�T�oc�?�ᣰ̈́���/��9��m���bbS��-���ϤΆ�U�;��4Z^ۆ*�6f�~똅t(��S�N9��'r�z>�t��K�/��~��ў���q��[�~�?�q�;�Ӽ��������&���C<?��0G0*��/��֑S��(b��-�y:rH�>��bU;8�cH�a�#�}ʭ��_4l�t֜�e�j9x�dV`0v��l�LW����o�r���t�$XnW�tC%b�A}a[|��KgB1>�"���`�P4s�Co�I8u��\���|4�*�뮵�u�Kk��΃~��Ł����4�~�7c'���,���&_a���ct��_1% ���鐆%T����
�`��#2��4�/Ŝ1M�Ҡ�>ʜ�O�v��e�V,��6O��C�`1u��Q&$Q��e�Z�J㓘�j����7��o���ϴ�����HM�K���%pH����-�S1B��%���?�^���\q<L��>�5�?\C��P�>��I�-�b�Ώ��ܑ�e}/���ur)�1GB_x��;.���$EՅ;U!��ͭgF`4� �5��mܐ'b�U��r0�9Eh\X����*]����`��(=��
'�u=�������_y��	#�&"��8{�����C��ڕ�gNR�<27��*�`)�Y�	�$����$]���xM��/p
�4a�c����}���Z��>AEb'�8����%	�TP[����x|\���$
��?�㳄�G��*D*J'C�g'[R+ y6>���r	�[��v4����8��)b�C��X�R��{�����[ ��x�L���9�����k�b���H'��-�Qz��Rs�GPf� ͝����J�Ҏ#7�r\��D�B���wjY���~R4�
��'�X=�A�5	�3���Ա����j B�~|Fe�v<���&�~��9-�&{}mŠ���s>]ҚRGD�5c����"�n�paZ��}d8�3E���2e� ��;�(n�ر�;�o�B�P�7�=�Zc���;�A-;�KvrD���Xf���ؽ����!`6�Q[Jg`�D�ˇ���#���c�-jG�4z�i�eMdG�����o$�dF�-��rA�M�8���1f��dy�'��Z��pZ�6��:� ������'w��� �l���e�9Ý	3 m:���4o1��'ې���U�#�*W���2�����&�qD�������a���0�.8[q�ͼn���/O��b�����O1�Z(iR19�)��jr8�Hs	���{_�"��<�Rwٌ�虳�m�����K��`m�ܿ|��g�p&�[����G�m��8ȯ �k��	�X�t��zMx?��^�&�~ ������^��v��$�{�s��-�Z�ٸ�Ԩc�o���������,����0���v1"�y�r���h�o�צ��I� E<��h#�k���'�����ymȹ��Fp�X|c��AaQϼ���%�c9�&g_�2Ȟ�> s�G�Oc	����(�L�;1��lP����'J�,�OI���*��*���H��/cd�ә-痄�B�I�q���G�<�8Z,�y֞!VM�2*����7�c=�:N#p��9_���e�CHF���S�n�k�u*C��zTҥ���Փھ�E\��~"�g̃2N�@:��WU.�7��<��zf`���X�t?�IAo�P!/��o�Q��mk���W���2�5�~�����W��<�(��f���C�@�lǳ��v�Gj�䯋��x�)�Xڽ%_�9*Z��8���	tHQ{U������=�I���T�5،�C�B>Y�a�L~�U�@���Po[Qp���*i�F�v׀�/�A�nT��=�4k��7)�aL`t(��"_C�4�zK�f����s�r��O>G?ir��z���?A�����ΣZ����z����z���i>r&47|,nWgBhu��:�AL%�5rKft��V@lل�Tu�L�����L�~��Ҧ��`'�r��QU���=�$��>�⧗�2_	�ߵ���a���NA�?���_|]Li^��X��B��q^I>�-X��/XaM��"sf=>~b
�) ��NUW�Ha��PYEx�M0G&���F��bԐ~��Ś Z�Ғ�ʆ/?*�\��4�|���3����i[�ct29��D���K��vܪ����h@���Gs�]��pw�xI��ř{m�~x:T�>�U[�/7cL�>3��?�F��Y�Zǟ�I����ob��+�E+(�#�9���_�����a�v���� o��(V�<��4dz���pa����]�nC��-o��<1FO1F�6Bjom��h�v%��Y�����2���I@! /�� 8@��R���	�r$ʶþ�7bC[ =����(�\�20�,�[*'��Z;L!�oXǩ�-&��y������9�	�/���(�� ���:��_W��Ug��s~�/�Z�a)y�ai��w���t��j�a:�r��H�#xy���b_6\���~�FwYh��I�kRa]XY��C�y�a
�����xbj%���=�i;v�*ߝv0���&�U��m�Y�Ώ�O7�̇�Θ�<�*?>�PDZ�	��$+���M�M�C=%��e�r04i��~��Y)��5���(E �&�ob{�����a��z�(�&^I'Bh| D^~������%p%��E$��XN���Oa���O2�JVA'u�J�#�n�Em��s�֬�~U�q�v��3�k{��V��bo��S���5�o%�j�&5�Ar�������c�nM��K���k��y�>��yz_��Q!mq��}���>ൡ8��>ʪ"&Q���D�p�w�9e������ط$����&h-'�9�k]f�]�
C�<FT�$��?-��ݍ���f��2���X,��/g8y҇�C	�=%P�(9(@)DQ�>�r:����@�� ځX$� V~)��X4b�"9�,�_C��n62�L�Po2|��P���4��j._=��׬@Z�u�,lk%!�S�o�ZƣX�n�o0���f�!�K�j�9"?o�ǨD�≁V���OqN
���'p�5
��8�̲t��WΡ�x�n�s�)�=ďQ��S��Cqܖ�ٴw���\rV��&�mO��**uS����� o��I�*A�@�q��}a�@u�E�P��(H�`"��v����0�E�x|�1�pBz��@�wH�M;�%�^�+�0�Ґ6��d�(Ap��^��ˑ[�s2���آ����s���]1�ek�n�NӅ�0͌��`-����c3��1!��8�;�Q�VdÞ�.�+ 
����*�mQ�)wY�\�A�$��1���_˾��,�&oP�%^��c��7[X��'!c�'�4� ʖ���`�Ǵ��ȋ�4K�H������F���P��Ս^��Qsx珏����ٛ�+�i�[B�Ȑ���SI���Y��τD��U�[�W�b\�f��w��}�Y��14ٷ�B>:�1��	��F�2T���R@�.@\#����+t3��ʢp�4j{Ê8�P�%�4G^ó�nRe�훔'���rث��W3փ�����;j�0$��SmuCyu����U��_"$:օ6���>T�:�$q��r�{8�gJ���l�9^�S�)}��̠	��aJMU�zt���N���]�ɽk)�)��pQ���.�a/�(��x��'��d�Or�� �7^J�s:0���k0pS����Ej3[r�_|�;�R�ų
~���B��9�]Bk�l^{-���O{P�ִ�P���}Gm<Sλ��)�ݬ?/.��$ļ�O�6��K���x�ۦm���L�{(pt:��]	Gm�ϧB!�*(!u�!��@u_4,�ÚM��t�>,sK�Zg�y;�f~���I��cV��q�?�y,���E�n��p�P����{�C��
�5��E!Q@��G�!E�D�CGf�\��P.�6U킂�T>@ٲ]F��gRw@Lz|���v��n��}}�� �q�B0�@�P���Ýe �(�mFw���L7��j ���������36�W�:��YQK'l�nJ9�w;�y�T�ŀټ8��lO~��V��S���j�M�b� ���{�a����w�*��CM~n���e&�[i�ߗ�K�>&�9�d�u�-�jZ�"�!�{s����ye�%A�5\��F���Hy�_@L9���w�,�[&UvI��6� Z�C��
|��S� `�����+Y�
N��^ �D;�<�s���~�{���1�XT��c�-�Ke��h#����^t�e��z�J�WB�+�		)`�ŝ�FG$��ǩ��o/�(���x��`|<��ѡ�!�ϩ��H�LҨ�ָ�ׄ^S��j/E\�jzF�t��!�M#����c���T� �/M�0��֞���5��Y=|�ؓ��^Z����,�����c*,�ҟ]�8����P$�����"x2�n�eA͏&�����J	�D��>���Ah{FxH �T8�V9�4 �J���[JS�
����v���w\ɥm�y�3�*�q��2��^ӄ��,�d�P^���S��lK�T��W�p▋?⟥ݰ@�D
�ٔ�F}/���w!�����ϒ��ٙm���ڢ�V��~�"�o߷�����kWz=|��Eg�v����^^�A0v��G�AƂ��\}�!�7w�%�<~6k������߃����w ��?JE��-޹+ߛ����s<a��p�e�x{V&/��v;�%�#�bV�3�����%�Z�f���ͦ6;���,j�I���Y�����B�����ճ��#ߓmA\}]��z:���H���&���\v�<������&#��F>�D�Cq��&$�_x(r��5YNrlQ0|]�;�~��O��3�����J5#;�Ag�q���#��IG�v8��M���e0k8�G�T��e�l����X����y����G���Vm��̕��3HW��e=r>�AL-�`�(d5�Q��!��7��`W�(c�П7�V<˓C�άO��C�/�껾���ٝ�ӫJz��ճ5���\�8��oT3���&Yq����R&� �noh)0��y{�TZ�1#�D���tK%����+.}	8��W�	g���2�-	l7<(q�fVk�-�����*'�@���zd���[�6�h�*�9�u�b j`�B'��#��ϯ����](zr����,a� J���&���!wV��<��UH����6Tx�"��bLٸ���)C}����C���e<������]�����b������R���\o�)�8��y`�ҿ6��d�u
Z]i���N%[��֧���X��x�4�NMD��},�����!dU�E�Dp^��pxw�u_)G�����O��.%)�&x0.��k����p�<�_����X�<+$Fs�^y	�o����b����˷�7�or�DĹ(94�ǥa~$�<�$N�ω[�3���$I�HB@Ѧ�����t���/i�g)A��#�u]�J���δ���`�M��4b�jw+����D��Z��b�
�C����\��RWBri\Q��H��ӡ鸶<���������sROi��2��vw<'��u\��>47�*���y�h*S�6��3<x�Y�|6�|B�������S�����W�co�ut��I�')=9���t���Xn��pxjX�F3Re0I�(!�1�K�(���6�$��dh�wz�Q�@��w�3���(���x���_n�W��,�s����Q���P"|�9�JC�=�R � ������z�hZ5��Np�Kv�!Ǌ����+5)RP�\���]cQ��
;`��C�D:���0es������$��6k��4���\�p�"J4S	$9�*�d�{��D�r>��T�_�
~h���H8��V�QO����n�� ������D�M�,7��������4���F��޵�hY+���U�t-$�;du�I�y]c���G�V�G��|�M� O���b*���q���qS��es���읽M�����l�	Z�	V�^ћ�CԥN��Nb$[A��(@���\/˚*�*�\�Hd��9e�\�ي�N�~�'��L��2q]̣~�ߠ,����̵���Ⱥa=�x��K�㲚�h���f9�-���%#r�N�x�p�����c�k|E׉�hV��Ol>��T�f\�!	���uˆ.��,v���wn��lˠ��}��;n������NAO��5X;���7F��{Y;��"ixE���ae~�6�}�id�k����4�ڳ��s�b���Q��b0�qƭ�BPH�ӿ��|ж��̰����(�F\j��}��ʫ��9�7�4����F"w����oF3k��+y}��=���	�-a�m7�
��}|jH@*��4�C��y�h�R
~нq�H�}��U��]H"��P�D�G2c)���ѐa��E���{�gs�Fk8I����|�j2C?А#�Ji�°c�;�Em�����=O7���O�2�̯��X&zP
�5�?�E��>�}i�k4>�Lu&�d��P�E0���d��R|�>*�]鑙��B#2���+���3�~D�l��Ny��TȐ/�V�s�ڼ�3;��&c���8"%j9��8a���O^Y�|��j�T=4տ���fj���h!_�vFb�cN�S?&�F:��c������]��:�dZ��3I*6��	xog�0@�ɳ5��L���G8�W�����bS又����4p(�����mM%4�\�,������W�F���u�P(��f-g�cQ�P��M'��Y�͌��'�6N������C@����?���K��= �H�?�sqsR���K��ع�Ё�r�I��j}�b2<�	�������A:�P䯰�Fl	0�3JT�D���~����� ��'�"�,J!��]�r	ro�Rq���n:�Q*AH_�%��{�����).���%�jM=���D�V~7�����ӯ{�����*s�zԆ�}����eu#'�hF��Ⲗ��h��mUu,feen?ܭ���][���Z������*�����t��K���D�zU�Shʭ5��ړ����d?*�*��:�{&�x����1����x4�	�D{��[o0�I�-0��W��pb�W4,�kb�����es��OԖ���}��SF�а02^w����G��Bt��'_���n�T<弐��"9`Lr���ri�����B���'͡��Wp�#�X�p�2
��:E����}=�J-�Ks���KyU�$��
� ������/�-�:���F�Ϩ"@O�z G��rQ�w���1;K�us�9[�S�W-d
Oɘ�����7��{�X�$Ύ�G�1��o&<_�>�a�� ���,OS�S_�ۉ#g�LX��^O�+����%t�R��#iH�'��=O�/������$J�N���=����A�g���zk.���g��9!dBu:���:L\�>�)�Y�.�
��ӛR���F� �5M.4���0�39�YX�W�ֺzK#7��+!�SԂ��!�?�ߒ7��5?�\I��1*��ˋ������s[�m~� �QܿH��Z�	��&z� �h!O;�(�gPm&�U��;"P3?k���1�Dַ��ER�Xj<�gD��Ԡ��h#%�� ����:�"I��O^��"-9+�%�2���� �i6�+K��O;]<e�a��?�]QxFA�Q��޻B!.�s�ϕBʨޯ.�Qq�,łg�D'籈طidS�����,�MM[9J�>.����\ۥ��N�1o��+����n}	�>�s�����z�����-R�5U�!��\�Ѹ�xb�UҤϮ�zF�-ت�+���k�t��l�]�DE���T9@e�@F�Mx��
W額�M�fs��#�]
҃���O����,[�Y�&�����u�d�.5t�����ٜ^��1��/@@+���"�Lӣ����<�(Qo�5�ȣD3�F�����i�z�½9��e	d�1��0'Jhy����m���p���#�u8��WV�3�Ҩ=�L�������F��Y�����D���ha����
X��2@'�?��q�:J��z�j��V(ƌ��!YO���ip�:r�T���ģ@�%<���ֱ��)GDvCo��Z��.��eEN�t����ï���Fr�F\K��w6��	k;�g�HC��ʬ|�#���sx;�.
�� K��;-J�+j
D�.�)�a��ͼ�K}�jh���`P�5h���J�Ӆ�J���צ3��ip�p�l,�����UpOd���"��N�z�B������{�����;�� ���@�����ic+�Y�'���atZ�l�X�T��xr�u�����9��v����%�F����}���1���6�˓3l�Qz�䝗7��?K.[�IQ���I/7�� ����Ж���ߣ<e+��h�\�z�.B'f'���؝W�6�n�ۧ�n7���O;rK��_T+��Պ�l;#b��55E ��	û�<:`��	#KDZu���$a�ZZ���g�q}E��ǩ���X�9ia�bK�D�Sئ���t�y���'���i��p����z0��9JE'�f�ΙG�д�e��+4�}q2�D�פ�i#�����!7�j{���^�b�t.$ʏt�w_/���ngb�M�i�ϒ��ʰ6�y����a����~DZ���ʻ��3.Cn�e���::p�s�jy����]�]����&{���"��^UЈHh"��[��l��qT�%�z'��n.ʗI����wL��`��fGo<�Vn�����_�om\�<
/��tj"��[�A.�0��6J���Aͷ�4��3Sߋ?��)2Z�����5��:�X��LX��hJ�q�F_Es�񿿔�yɇ�R�p�hd���*�~�pB�X�e��a+d�T�:I(>��Yo�|��;ǁ��DlK_�� HGZb�?�G�y�fxͿJIY9,�Ѻ+."�2X��E9.���aD� �� �g�l���t%�ˆM���m��n������g��!g�u�E�r�҇�9�e�V���:����K�����AY=�cr�ͫ��ƶe']�˒���S��JT���1�Bx�3��	�O)P? �ڣ��1:t��� �x���%�D���}��I!��h�&��Ր����f9�Quu^^���#�����O�%������=(ͫ�����1�!NlV�YS��7c��`�'�o=,������jō����C�1����Ea��>x5	G��)���N��.=��$�̘��Hf��턋*� ��1���<�k�(�������)�y=�ˮ�K��X~l���á�?���m��4̊�ob�I���Ŭ��5H I�QEN����c�����8Pi����d�yǙ�)�uh���cR�S�Y�Ƶ��1cQ��Zn��Qv"t��;����)��8[��OQ�|B:.��u�����-�e��[O�sw�Aȇ��'����:�gB�4h�%ٕ^c�~r�ؚLjP�)B��- ��.�]<џ  �^(�'��C`\	4����n���x(�3af��-i�Q��0o�e�ȱ���@dE24X����!MI谝��֪wPo��lR�N��y��N~��2A仚KbANʮ�+4!ͻ����$��^
A#�꒷1 �#]�^2k�r�Y(�m�0��T�t��q�9�O�}�Fy
0�J��R��� N̫�x'{������o����7�b	�l��j��3r!׵���-�����3��A{,L?�n��{�wbL=��r���`-�u}}n�:��XYN�%��կ^x\��:n�^��Ɨ��t�kc���>9݈�G���վ-��nG�-����w1��������z��ORy'J&�!�t�Aީ{���kЬ�ӓ��ע���D]ȳ�JO�J�������o��X�u�Eb� ���7�!q2�M�D�0��i$om�d��\kLb�����O��K�gԺ��4)2(�LX>�6�C=�l�|�����B�!��U7���جʌ9��G�"��Gk��E�jg?+}�Xn�T��ĉτ큵���������չ����i��
aAF̓q��v��s"o���'pAE+s��ڜ�8�����i	Q��y�7�lvV��^�c57������u����0���P��3ĕ��S�����!�-��oKPD,�g�!��_˸n����ຍ����F�܎�A���8)-0J|����%*z�|�*���_������4?/�C9��]��k��P�))X��y�,p^V��7��	s�PDt��܆�GP�B�B�����!�-2�4�ھ��:���6�x��Jt?x�.u�2�u����c{h�؅Д�4�Q�3�B��C�D�\�c�s�]ď�4%�䢓`M�5Ƙ
��a�j�8��ǚ�c4l�E����k��B�=sO�u��S�GFb�*�����=~u�9#
���j�2�YT�,�����-����$�Ͻ�Z�	�)�a��}���e���=���y+{&d�SY�7�%�~N��� X�A�bW�6��A��A�̠͘��9��t>�g`�̏�x���9A�G���Ú�M�$����P���i���'g`�oQ.M��m���B���]wRJG��R��z��"~uo�QN~q����`��K���t8
`�-�"3�喃�BB���>�9\v�,�XK�2��6��r�ԢCʙ~�$��x�/1�o=�:��I̢%�>�HIR����-iK���o�����b��9�����68���A���b�6ߨ�쉪��ߡ�iũ��X ��>�_6���R$�Jl)�>��YL(�*l�~.�;8Q�ulr[�%7c�%H��R&9��$���&�ڥ��j�y�w�mU83!� U��t�i-�m��DV���?:
v\Xӿp�@�����s� D�.4�Gx�����z��<3!W{" /_�M��<�b��X��yS��	��F}g�!!�h�kP�͹�	]+�O�����Dj�h���u������硊7�b���ƃ�'5Y�	PaH92M\#���%���0Ե��"A�����:���������:��Z�u��>����me���xˌ@ԲQ��m��7#ҿ�A�C�D��.��6	S��ZKu~;y����������t{�Nde�� ��p������~s�wt��w�b}eD}9(�у%���0(N�M�s�f�?��؜���^ �R7F��ܩ(~�� �ٓ5%�[''s�ߊ׵މ�/�*�|��7���n�6|�R��+}�pC��m�u��K�b~&�QTY��YȈ�!��1����H����eA09����+��p|�H���'�*PC����?��Wɸ���Խo��=�j��k�j�c,�#1��l�~�B;Si���+�nE�T1M��P
���9j�8f<�k_�Ћ�+�BKK�j��_�˟���\�;��M����+F�b�,Ҝ�3�E{)�ƚ�3�9�FYUNW���g���>��5-֔�e��(y�!�ӧ��L:����D��;T�6䌒��\��
�F`�VȈ�f�����4`��u$�R�/����rA�ـ����A��\aT��4�N�/Aﾋ��XWE���������!�]m�-������޲(�z���y���$=�� sw��;J�|��r�5	����t�K�0���vs_�|��I�:>���<�߱�����;�I#�W��i�}�8P%V蚒V)|O�t�`,i�hR�'���T����a�=�R���yP���8�;���MU�yG��� �O�D}���GXǂ7�B�e˗���?¬��-���D�C`<�jp��S͉�@YZxϨj���o���WV�7_�A�����_��a$�m��˲8sX0R}�I���yZA>��R
T�0k�D��5�'&YE���`�˨�Os�3a�a��_):D���!���:k������9o[[F��RfZ�=����M��D܆6�'݃)OIFʳ���=A��)�Λ��O�«\�R�P�l��t�4�Ї�O�
�q�\�m_D�%j��ȏK��g����L�2���W�+"_\��鋽��ĳ�v��)��'	NzN�E	�[�*��������IG�eA��R�u�N���-9gc�DG�V�6�J�Tc�h�6�,DdvY"��N��0)�?�o��B�� �I�����S���Op#�����6�cs��}�;e�u�W�ūQt+�Ez��l���7�g�0)bm����L�sq%G%7�wx0�X�J}H4�m�q	�~�B�Ӥ��+9K�w\f ���J[����-�*OP�4m�s(T�]G��.���S��H�p�iT�hA����j��oe��e�묁2������)�+<෩���J=������{��@o�,�05��1��-蜿���?[�CEEǝ��9!֊8[ d�gG���Ce/*ײ�cJ#��ur	��Q��#4G;��B'".��gٵ�/V�����ۭ'��GvHe��#�����=wW���|��;�u�";�=xy�y�B���Ұ��Ҷ�Wxi���b�_���?)�Qe	0b�C�&�L)CG�+>��4�����(��'�:U�;��<Zݨ{� 0���v�	&���M6��������狐�c�w���cߎ8��]^��ܤ����O]Y��zޙ0��+j��n�=�5�j�#L� ��'1}U�*��{� �y�A	�^��F�_Z-Ūd��S%�>�G�՝��@�	����-	����T�v���eY;��a4}֞�ס8DC�O*y�)�]8
tKA���N��^a:Q�d��R>��K<�'\��I��o��/���ٚ��oS|�J�qv��#
��&c���ͼ�-�<��J��6���
��s�!�i���ȴ��p�\�2	�9my��h.�-�~]�|���ϞX���v�O^��w�X��/Z� ��?��WN�S��f���4EK��I�����bŌ��
}�ѺYMY�x* ��\i�\-�М��H��ǇP��v:pb�.aTn�ƶ���t⸝+��$u��֮0�B�Y<*�����ɠ�2�%Un;���j&���<���Ő�@7:
T�Շ$��n��Ytc��<l�8���,w����X-MWH  ����d�U]p�7�NU��D"�PʸC�(�*�L�^�Ho�M.����)�!���4��n�5����K���W���
�i��Q7	�n��������|&uOZ�*�@��?���ԽF��;�_���Oq�҂#�	E�fE3�#y���
�x$mwpY�8�����eX�|/~���5�^bfJ��']�d�_�큟R��Y�^ݛ��ꁈ�6�TXMV*��n%5z�h0W��Cv�U�H����uds�7K(�N�\]gW
�I�b��l@L�bϰQ�C�< y�$۔(��чnf��w��5�,B�#B"uD������v'���X�t�����)&�6#��ß��F������{��6�����8�Z�7���Z�����ݥf�%��Q�٨�d��ؕ���	ҋ3۰ҪѮ��3�w���p#�x�SҚ��(2#p��h���<����G�v�[N�p!4��cƃ����e�y���r>�.�0/m�t�
e=I,��8�㨘H��'�vC�G��i��ݪL�s�In�X���^�4"�%�h���sL��pC;VZ����NQ���B���y1�˶�|2���ŵ�F1$FWQ����A8?�x��8�j<����l���2��/Yr�3�-��+�="P	pjK�7A�)Mw)��9ؠ3E��
��������L�ȡ�欤ם�&np~N��& �ƎȣL%l��:�D5�{����6n]��~<-k�Rc+H�_WS�)��[�b`<z�mhA,rME�A�,CmiisL,U�l���\�e~ͥ�����s�a�n ܪ�v}���2��C��{x�W��(*�@aZ�֩Q��O'�9��tW�7&R\c�2���s�J���"��i�2�#O]n~P2.-��A��^��ĕ��p޲��9l'e�v����fI�����M����v
HM�Gȷǀ�ɸ>�|��q��b159%����6�t�p��-^޿U�3G2���om�zd�:}�K����>�X�� ���o 4�}}���c�<���s�zh�n��dwF`��"�?ϝ�Ykxp���뿢�qXB�	�7&�0uw��	>M�w<!��
�89��-��@�P{֙�v̤��\�7���[	�j�V�>+
;�.�u��rӄ)�r�*xR��a}�?�[0���P��ʟ�4#�*��������<�~҄W���� ��j/D����D�B}� b�?Y�)C'�M��x����C�� ��f�E*sR�X���N$<(ک������A���H�v�S�_^�绩�U|ܣ�����m|
�U�*ΡV����{�d2�D�A�2��عV����9	��u�TM)���ȂYp[����XC����Rw23`�q��:s4�c�"X�$Q��&�'�7�)�:W��&���=��Rd�r���6u i'�L����\�6LV�����V���*�4~�p�	~��	�v��k��U�>*\�xO�zu�+FB��b*�y�"ݕ�W��C<�Q�o ��L\L�V���6J2���!B��"��
5��V�/�6������3��{�W����V }T�� J����K�گ��~t,��jR1c*|�]s_,o!:iJ�k�6�֨,k�����m��Ѫ�N����0�S�M�¤1u(IM�fSa���������n{9�k=9b_���^��ىC%p8D3pVz�rùa�<
aÐ�w�˽;�2��NR)���dF�v	~�B��;�g���� Śe��'&��.<U�%�K6�q��/���������}���"G���9��E��)�{Go�f�"Ҥ�ϒa����p�w߻�c���C����~AńC`��M�-IM��x���U��+��2wc���
����V���-�*��s<�F'��a�"�I�N���~0S#��������2��iX:	"�S���,a(��&��#���	�~w�h��~��/ya�xw�`��&�W3�$��Ϡ�_ڛ��M� �m���ܩ`�!:r&3!߲���~^��e�N^�e\ ��N�k���uB6�fhq�пl(hP�Z��8K�;=U<�+и�Y���Y�6�����R��|1�b.�F5S��S6��Wp@�@+p�V��o�g٦N��RO�?�M3����l�W�����D���A�B)T��q� �r�2�
ۮ)"�`�yF�Z�ស�_���7_�ڄ�U��i�: ��'�\7Mu�ԩH� $*��+7q�y2�s�^�B3�U��}Jˢ��f):%,�Rw�S�G������Ա�H�Kc�a/��)�5 � �'�n�w�*�B.�>�E�T�7�e���0��ƣ�����<�SPk��U��,
�+�;�~3ЅTD����fcn`��نٔ�Ǭå̉��na/t��6q����~sٺ�OlT�j��������W�\�{��疀㔼p�y�}5D��5�s����VN�rLCd��ߙ�a�)�,��.��i�>�~�1�̩z�q���g�G6eyю�,;�W�P��e,\6an�e�s:��i y��Җ=�0_Ǳ}�e�P�3���y`��7���j�6�,����E���u�
*�e��!���H��%�
��G�Nh���k�u1��Er*�b�׏����ֽ�
�byl8�̈$�o�Y1�~�\F/�R�`X���wL!Һ!Y�x5$�5Dg�e�6���? r�@�.�_΅�kp[�5-�H7��`B!f�/�w(���:��޾�]u��E>�(����
!+%M��վK�zV���`���ZT�ƻ����{'����~y��@�#o9r�9�@=K>R�I籄�W]
e]��kT_��v�չ�%g�u�e#6����o�}Y�Fe޳@\�ɹ�u�W�2Wy�&v\P���1�?����$^���ݭ�6hU�*�Ƽ'X���Bo#�u�&�堤Z���4en��>��I����� [���^�1�\���A�ڠ�U Xz!�cÃ0����ӱ'�ʢZ��}}lt6��:��fּ{�f�#w9t1���w/��P[n	
��l4/S]2����X:�D[�%�L��]��7�f������;���j��9<ʹa���m �u`��v��sj��o�o��A4�|1���aI"�h�苜�`�F��-��ΑD�}���	�:=$�s3\�U���jPs�2B�i�Iݔ�D ���`�q/�JN~����.�7��Elq�]���J�
O͐;��������hI�!�G�]T=�g �D��ʲwa���P�r�R�A��)�%�YEc���Đ�{�x��}�ȓ�ݙЖ�U�b���nW	�Eu�;��d�Tp(�e��?4n��F=�̑s���;Mx볾.�:����CcA���h���/W�]��?�n(R�b?�c����CR��D:B�g�*�	��=���c��=I��S����9G0�)0}ۑ���1�`��檧*}��]+h�g�8b ��x�W��
)B�:g�P �fHw�=Y�h��ި�ʭzd��s;"�O+Xm/�Zb�����O~�5��!#ߌ<�C/��[@�ջA��vK/����[���d����X�`?��.��P3�#�������U=�̂Q�yޫB'Y5�[E$�9B�0����$<Zu����^��X��$Ж��et���	@mVIF�x8ٯ
���I5���8환@kE���,�r���v�.Lp��3ќ{�㟰۪(r�O�nAlN��(�]� ��|#��~ׁ}��k�Z��@�d�L+A\3��0͈�L�'�U��a���\��+�s~bG�~��ͻ̇�4Í�\#}_YZ�l�h�~P�`�iMV7���F��  g�3�l��A��������Ε$�$Х�|�@���׉u=��*�S؅r�p����Cl��|�����a���XO�����g��g`��<����w�gN��n;r�J9�a��p��׶ܺ�I�qަ�ӹD7���Gv%��*%I�p�M�vJ�h�]��3_�袡��o�18�C&��_�]`Ϧ$����h�t{v�-7����3�3>S�����j:�ո�\� Tг��vG�Ҵ0�`�i��+��P��F\=&�m��<���=�*~�7X�����%=�6�)+�m���8�-·��`�AEY��tR�s���΄�f������룢kWr�Bh.Ϻusko�c����Z��o���@Ħ�kYQu}�!{�h��v2�-���5!̃zf|cC�λ�3^_0��)|�5 `G��#�Su���Z��>e<���}S�ɝ�rT3���X*���W�P~��n�<���3��������-�
�ދ��BwOi��ٰ7��A�81^���Wi��U��Gt�|tn�G =�p�`&+ޥ/�'�Ej�n�:
��F�7$�R�'���ne�q�{�����$����q����J�ݫ�լ� �g�<H�-Q�u����mBJm�Y��)?�Ы^�9�v&��)��Ȭ��S�
����)�{'��'�'TE��#� �'�i�/���o4>��i�
�HR9�%{��&�85.���6yx��yR����@w���N38R;=<?kh�N
b�&Le=`{��Y�.�̑u,va�F��pi���sª+�s�4k6��.=T�\z��h�o[>�����E2�Ja:$;��޼��w�f2�㔘H��������|'�Gguw]{����o/(b�2s�����L̸X�yE�r�%�V�bbv�:,��z,�j�q��)���ù�A��3���r~�)�@�)��8ɵi���6G:
�:yO�T"�o�Q�`*�Ȣf���Y�gZ�Ue}T}�t`]O��Saa�=�#b�L>3�¯*jex�,��L��=w���u7�15I��m�WH���I�,Rہx$�K��[�V�:�Ekot��
��k�����y��b�����_�)��w#s���H�L�T�w����L�����!�뻼������_�"�"O:���޼���m{U8����ö �<~soo��j@���:�惤Ԏ ݾO$
���?�"R�{E�P+a��f�6e��Y����2�H</:��ܬ�ݯ����*dx��.��-�D6�E��z���V�j�-c�M�zgP�͓m~���u�E��	�<�#��[Y%�"�c���wu����1�7�wb�.k�h��U�z���#�k��#�M)��V�	���{f�L[H��8�=<,�0����5��[�d����v��T�y�_�P�P�嘍���n� �}��i,�м��n��m@�����\�J0Km�0�Ц�)��<�e�y$$�A`*���;�6����<�+7�t(���{s��*����`���8Pi-��O��=I����n�P�/�f,���Es^�߫�x>_�Y���k	���eju\R�u?�Yϣ苖:P���s��dW��_[&H��`��\�/a���/��  -�+d%���������ʭ�i>���:$�a��c�}!d����kU@&b4�z�N��C�h9�Ir��?��vN�OVI"���|c�
���vgF�����W��1���!�8�=���!�L��s�� T��a���l��%G�]�2����4>r�B`m�3e�n���"Ӹ�B�i8I�4g�;q$P�m���Q�/�`F}�i��O��{��[����l0�G\�e��J��4��xC&4&O���f����R�����a�Xj䫨�53��� {N��\��s�u�J�,�4]��}3��Pa=��I˚��#)Z3��\�.�坋h<T�^��'d��N��O�n
���,����ŵh6��t*Ί�<��dxr��,�%CD5l����R��G�n��#�|��[۷��x<4cT�$K���=M�Tr�F%��o���22�m�D��'X��c�\�E���NӘ{s�5V��1ш�O_����	ؽ̜&9�:��X�6]�d�Ʌ���2vc��S��$Eڱ߇�V�H��I>.��z�U���zY1���J�2�Ⱥ7�gďU�0|$�X�%V:�~����]D�n������� �S/֐�x��� ��jn3��� R�����]&�J�_/܉ߚa�n123��HO�����t�R�������~���˾,q
p5�u]kL'��;�7>����5�/rmGRqQ�_f�a}�K~37�\$�ƩN��K�~���}W�Ue>	��"��K��L��'�#�k�33�e����|ER9�gP�������/������!P����*&u�g��O�����K�(
�F�48��9q/�y�7�Xc���=��|�u�\X2���E$�m�/��L6�4��������k2^�������|�3�v*B"7_��������^��X��ؑb�y����Ռ�-oE-�2)i��)������ωč�H.�1�i�!�V���m��'"�s���NV�"�;]�A!��Fx�J}z�XYcu����i�{�7���i]�X�2�ʈg�֘Ӵ��a��N*�D��� `Q��Bgs��4zc)�`��g�6�눕J�T4e2B
�ι������Y'��'Uk����q�G2'�d��ǨsHi`e�d��Rx�?;�"����B�!���>ć#�k 7�Hi�}Sq��VZ�Q���ڸ�t��o������]�PH�:^�b���k`
Jc�w��I�'���Q=����l�:�ѯ5²��:J�� �R����*�%Z�
�M�1�}u�YS��".ƙ� J�3o�S/���VU��I$���r!)���s��)�JS	I��\����͠�gl��.1�C"vm���TY|9�/3tV�y�G3d�,Jb�!J%�ە�h�8[lN而[�4�]�ͽS��Uߐ��iK���@�����{lլ@�D�.:X3��	�9�=L�_�#�d*�K�}�ȼ8l-
̲v:Y��p5�݌�x>���4H��eHGB�S^��hů�L�f�q�p'��8ԑ?WN|7��h���F�U��)�"y�a�(?�=}%�O� y��i3�;v��[H�� ��Y`)�ᡓ�kS@n��6��⬘�[���;��M��8�rɁ��$$H�u*�=?�A)8��j�j���`<ox�H{�z#֋�u%���#xI����S���b������]�m�:k�6
�	%gHbxi�qǎE� kK�����;�Ե�!zBc�y9LkdT2�ǆ;���	dB��s_�m�҆�2���Y�Q�8��<��S�g�����9�D6�V~���D�4���*ˁa������O��o��?O�7{;�p�'��Ќ�Ʃ�ܑyg�½"EI���Eip�-����%���ڵ��Ɠ���En�T��8
��eP��9oz�ޖ��F׼�V��%C��AV1f2?i �J=�`h�8.7˰���tD�`)�"���ɴ܃�7�k����˳g�A�ei+W����
o�m���Ԛ%N #8?XE^$Z1�$x�O�/����z<�fBt���}d��2��$�!zQ����6#�o)�7s/��_�u/$�b��x����Q���
8�7� 23�#]�^[��4Jھ��|~�݇�}M��i�FĲv�61b$���-���)���f���]�#^�e�^m�vWp�\C׵'nw��(4�����6�9zv�������;�5��]��%sOW��*<�՛Y��މ��f�U�P_�\�cF!Ļ�����[tQC�fW��Xh��3��I����.릤l+;
Ql���?#z����(���WnO�k�V��<fNDb7�RjZx�;��.:��$��~��!��Ld'/#����*�Ҿ=�+��վ��H�J�=ܛ�镅�K&��S���K>�sw5��ɞ�/z�t��@�t2G�'Q����U� �U�{%x��N��N���b�
�=��Lb����,��P���rM��ӹ2�KO�Dl���D,%��Lxd8ݓ�:�2h���>N����Ւ�Y�{��O'� uLp�0u���.(l�!m���*	��{�"�(T-_�*�ʜi;�|/�Cb��K�(l� <}A���i�pym�T�Z� ��5���L)�D�(�ӝhi��q\q���I9������S���揔�`���Y�w�Y���N�-���޴q,��yp���X�u�� 7���>X���X�A�L%�C��:�a�!8�'����*L���
+�u������;���kf��5��Y��v(� �kt��c���Ο�y����Ӧ��څ�_3+�������K��A�}S�HT��K*��m.\Y,�V����S r�H_���<�����·9�Fӎw�93��·_9!��JP���8RF�	�YN���X�{�������(A�Ԉ�_u��=)�%7���Ѓ�JQ 5�C��J�H=L>G:5�B?T��jb� HxUX��?0��-\�QvV�["��C��2T�� �|�*{����_hU@�'d��Z�6L�i������,�yK~�?uF���D����Lb2Tc�����"��x�o<�;Ca��6�����A8���Rި$����_~�T�,��st0���-ryǺp�5ٹ�bW��">7d���	��}ug`�VA�E��b��3إA�1�c����f*����kL~�Mm�ar,��j�f�����m[��0���ר(U���m|��_ճ�mrW�Yf�:��(Bq:�.E4�9	1K��&;5>�d@��q�ԊΦ��Z��Gw�$#GӍ�3��@�G�.���,�"�;���(z@��s���sQ��;��}~&;�wd+]�g�����g��T�)��ެY�o�TH�4�b�P��E@�������fǯbl�=o�Sژw�% �,�B��8H	ȓ�=9]�&R�t�?�S,�e��� 7׃#A������h#m������2�~��ۧ�%e��^�y'�ŤX�<����-A����3].g�F�0mZ�+q��6`$�,���&��ސ��Z�����Z|x^��ft�6��ϴ	��h�I�PC��ɸ-�CA`phJ���.bA��O�J�S��7��:F��s�����b"���o傍�2B�sȭ�q�]R �İ�YNv�S3���5���*��F#�$�&�=�s]��Q������J���=�\�Ry�Ynk��勠ݩd^yD�p��@��A���W_9���g2�\�j~����VCF�丈d��~y��,}�ؙ�L�E�W�M�Mr�	���H�@J�9�s��L�3��g+���1�>(���P#�0�k�5�a�<�`�ަƱ���T�@{2�i-��փ�*(�a
���Ƽo4թeؖ��bk�Ч�$-�����G����P�������G -pƓ�o�(p������a�<�R���o�y��&��P�Ҡda%[կb�F=�C�q�(���6�d�.�q�W
D�G���G���֥��5a�61���hH2��B�s�1��;�Tb�׳����V�z5�zy�[Xѐ�g�<�]Z�P��"k��BG���j�4a��*gdD���h��M3z�P�x����#q�vi�~<��:�4 �{�.%=�,I�"���)�`>��[�e�J���<��R*��C+� j���_�t7����ʤ�����(_p*�R�\�.��S�uN���1�i<�M��#�����>��d��z���G���,�a�;�n�Jk�=���R(���C�IA��*yMtP�"8�T۳���c�%l��B~��m@�W7BtUɻ�۟���/���<��x��l�u�3G�
�z0n�{��g@��9-�ᨪ��G���,���X�Rs�3��K�!�7SŢ)ז`�tvթ���qA�y�K0��ٜ�!�Z�:�L��46��)�~(�n�k��'��9D�yNF֡���ܠ��J��]wI.���˓��p�c�����2�:�0,l�R������f^^r���5���?>�Ǚ��I\���?��� $�P?�r��W^�S�U�?�T-F%�H&{c������,|N4a.|mR7�MQѣ���1z�l=��ǿXkо��W*��MwXg�&�҃���{W���k�!E�|8?����w3*+�/sDA
����@�x��A�����BY9�K���i���Ҥ"֜�z���g�/�-FJ��8/��QU�������o�y���"�����Iv��0�\/�P���>#��t�\i��[Hf��C@zcY�LgDcQ^��RMFN\��Y?�Ҿ^^��2�cw~��+�Y%�ӎ����h]����)���� ͅ0*ns�Z�����b�J�HK����bp���o���o�2�(E��-��+�9���N��l;Z�aZ�'3���e�ހ�J��Oe!���������������BVJ���:jҁ�
q^��Ŝ�T�=���q�h4�B�
�6E|�~�k�0�K���:��=����m�=�3�/J�3�吼�*�K���c��.�FN;G||3cmX�'�eU�����8�u����{F�^���E�Q�l7,?��ኚs��Qٻ^v/��W��!�VBH�4�7�d�����B���sjc{�W��v/$���	b��#�`�%�g	�!�Or�hIY����}��Mǅa��6wW0K��xz+��.�'D������U���!���*K��o���V/����ܼ!x�Gg�7�6��a:Ake��eX=B�</z}��?�X^���Z2���s�˳�W�]��|�Pj���b"+��.�
$%��U�J��~6�b�R��Joh>^��l��G�-BvC�ӑ��I�ȭ�*⮑��A"� �3ʹ ~���|�4]{�9��Zu�R{q8�^'Ĵ�,��O��1<4��>����X��K݀t�UM�l[�Q%��C(+f1�
��5���"�2��.���f�R������+��V�o�R�����|�
��\?���
���I5${x�?S��!u��doͶg\�}Ԑa�U�[�S��x��q�B�q�Rٿ�P���(������[�:#t/�	�(��s���V�{޸Y�aR(`�E}ux8þ����$��6�5�Z�.,Ha����-�E�s�k7~�':	n&B��7�SF�d�O>�<f{���+�BE�I�`9���C�r�\�ДWo\��:���ȓ�nɳ��&"���e�2H�e|x3\���-}�%gQl� Ś�"%qNYI0C��R��9-���޾��㭗;D�<\�|ҫ"^6e�� b8^a����ew�I`o�?N.'�ݤ��+��@�t�$PK�����j��%�)�P"vp��~�$��C菪y�Qῴ����M�Yl]R�fX�#�Nq'��=��?�7QHM�ӽ�?�i��دO4`�PZ�ң@o�ZA��pҭB���Րk��9\n��JT-'�����;��t�+�J'nrd��-#��	�'���u�l�����q��*un�9Vc���Ĝ��>�|�r^�`C@%%��Zf9�}b�E_�4k-��7���Z�U��r������Y?[�(���ڻ��M\9��gi�k��Ҝ�� �͋!�;$�'�o�H �2͑WSر
	T]t�Q���qXk}í4�����[<*��_��N��1���|F�Z)�zGV�� O�����ƙ���Yf�j���n�Uڋ=���U���@2��<��b��xv�R�jAq��?�/�c~�~$�	���[�P5��ioH�]*��)�4���#�&n��+�h��hFHqB%�,�=��p�!���#�s�r�f��=r4Hxa���d|�վ1ku�ɔY�@�Ƨ�@�@](7��.�U���ҭKMd�ԇVG�]��(���"/g�..b���zD7��2_��M?�cO��7E�r������`���� £�j�oͮͼ��d�	RI�����;�q]��7�ܓ�>ќ#�A��Rul��^Q3 &�xtap��6d�W�M>t�ս0	��K��i9+�>.�"]TBAK��Mj4G�K����]?c��f��gƻ�0 �,7��)�5�2���t��_[qD+2Az�'l��5=yGȄ��nj&��=�U���0E�Īt����M������!1�&��ME��yQ�� ����W7'>�*�k!!$�;� 78/�\���خ�9#����7�Q\dkУ_c�[��b^�s��岪�H"�v�M5-��+ܣ$b=
(��g�h#��mˇ��]GM�	8�1]� ���2�Tc�Y�%�_��9@��)���&6��B���L�:uw�ڐ�������ޢ;�w}��-d5����3vJoUa�Y�4���grù��9-��(��U;�j@���_U?K{�zՁո�ڠ��0<�Z�@��2��JI]�L�!oQ2?Ѳ]�B���do�+(�y�l�����4�[])4q�F�N2�[��+�&}��TQҠ�.y%�}��,�JܬX���J,��5+Lx&�;,{��p��cY�|�LIE/�,�$϶�Iݛt�<�F�g�J}/�����W�dp�",U?RwXaaf�?�9I�.� <�2�5b��a��_��D���u�1��[,n¾��3�iH��b"�A�bX����6Eͅ^�u�N�S�_ �.��|�C�|��_�_�VݓQ8��� ��][\/VT��'�Pk�.u�*E!θ]�ڥ�x��^����ΐ3a��yV�:V��x�&f,�-Vzz�>o�S�]P��4�kHI�2�	�ru��su��[��Ė���Ğ���#-4����i�T��g�v͗��n�y�~L���f�/��vJ'S�&��;=@�ƴ�d���@���Bb]��K�E��B{��T��
?�_�&5
@�a7�rn�$f�c�p5D����u#������_9��:%��W�&�.�g��teя ����`X4Y������rI�S�fo�����|���޿�����O�cU=[�	���^���pV�V����!}�D��ѓÂ�P�7�ǈL�w��WR�0�C�R��q�T[�������l���eѲw�E&
$�y|#+�O�h"���4(Ϣ���I����@~~m�xMĈ*nώ�Q���e�&Zoķ���*�*3��B���z���p�0F_f��-��k�Q`��"
q�E�,V�OG�
6פ�<�5����#m{M�}����#�b`{�+{psn�ʯ�@�M���쐈y����zJ]%\�E���.���X:;�b��F���L=���?�
�"�N������M;����PR����-�,�����߅Ve�BK�C� /���u��D�*����1�
9,�u+��ja��:&��,&ق�K�{�p� SQ@�|��76����F����Ĭ�ť�E�M�V���;�%l_�.Q����yr�![��5Fa���m�/���NasGF�)ČHI���yu��%�뇌��!E�w5���$5:)�p٭�L��l$����=EDE��r.�gZ�ùl�?���S?5�l���I+.˪������,�E9����e�!�X��R/t�3a�{��{�G�bM�p
�EDb�@d���X�H)Z[yrS�$?c5T�L.K r�%w��5@\���!�>f��k�?{�a*s�r��mڮPŴ�����	�(���:��HF�#���Ӱb�?^3�'���a��q�Xc�����:�Zl^8�vM��?Q�-�A��۟�̑\S�'��A�|� ����׽�j�)��M?Q%Kne���<!��K���JJ�j��h�4��{ �F�&j>��\q��걐x�y�ф.��j|��ɥVU�+��*�i��Q�ʿ�)D
y��""/r��Q���(���+0Ô:��w� �NȤq�c����'m��6�xK�B�eO��QР*UwB��a��(���oyYa:"�W��ߨ�ru�����&;��,_;�h
�8�	)����䯎�g����������<MOFf�1�f�u�7Z���g`�<�h*���I��OtVȯ��'ZMdfW�����u���U�Wg�F�[��g0�/��[�i}ޞ�"��Ar,\�}wB�M%:�ƌ��*��*ro&�>�o"B5�w��U����Qrڕ>-N��$k,]�Mڒ�,�����Y<��Y�M�ȸ��GY�>r�_�#�C��
~��z�<�Mj��=d���h����c%.�n|>q��,[h��h��$�B ���R�,%��_�aq�O\�X�f�=$sC�8Ie^� ���u���2oqq9CT�Z�٣;�z\tv	�f��ӟ���v�b0��}`%-�*mi�(��J�z���%45��%)C	��8?{~�B�?ϿM�c0�g�N���m�:��A�C��w����ג|��'��:��o�D�f�g��˛s�YV�����Q����Y�����vI!ny����8%Y�^�e_E��Ss��D/��*���hwR�O �S1���;�)��8���OeN��Ѳ}w��; �2&��{��0��(�6�F��l�q@f=B;gs�J���-�!l��"^-�K���h(������s؏d�) _�	���+Ύ��4�`�P/��Y9U��J)_��8sh̸��:��t��3���mzZ�����$��҄X(s@SG�������<�Ǳ9�W�+�b�3+>ĦGlL���X��ֵ��NN�;Bo�����xt�|9�Yeʉ���M����}��;J�
��[r1��B�'���;�\�O��LJ��tlK����XJ"@��������F+
��j��
�"g�]�is��*�je�Y=ٵ�c���BޫuL���ʹ����>D�Jw�;�=X��jӲj�c�S��Г���@�S<�>��x|萲�ķ�ΌB-���|�zuIJ{�9� �J�԰�����U���w���ݨ�'�t���9X?��@t�d+��@M��וֹ��f�B�^�u@2�Y����P0�*�0 ��(櫵L�&�O��؈�+������2��	��4"o*2���n�K%-��Um��
���}��g��݃�;A7]1��b�����|�g���K�uٷ�'����%�{S���#�T��~3]&Y�Rv׎�4��*x�Y~��^�m��S@6b��ι����F��Tٿby~�����oCXF�M�@N���!��y$a9�[�x
¢�ܯU$�ck^��p��2Y���Ht��Go��l��9ۂ�d�V���Џ��*��G�Y!�:c�
���]ڀQ*�OT��.g!�h�C�@�="�����Җ�����$j�7A��Q@��!�Ӯ��E�M4ʎM�)���yۨk`ň�"ޜ�B�@�d0�mݴd�6���N%w�u �G���I�$�\�7�h�Ic��"�35}����%�e$��ZF�ʫ�.!�a��ú���<A�7�g|Ij&��f{�x���e�ɔJ���O%���ּ�q�����x�����~!��B/4�譬���X �c|�"ḥї�l��nt*q�L��6N�@�u!�V���ΊB�;��Dn9���li����Rx�%�sH�s�3V;%t��RLz�O� �������UN�:�]�����[�2�B���(�Cv̴q%���i�'�N�񝵐�7ɺ��& �LG��yB�G���%^��k���[�V��t������1%�ZT�ym�wy��Iq:�N����cd�P�Y���/����z���/ǝ1�H���"?� �>���ķC?�e�\3(�n�B��p�e���U0�qhQ���d���qsj	�@x)V�e��Zi�ѽ KБ?�9Q[�h�6�J�#x�5�_�2��և��_ ���YX8�=Z�%Ch�Ò�����H��lnh�0�Ĭ�|�D8F�)�i���U�Ȳ�X�j�p��g0~8��x�G��c�����'ӗ�_Ҷ�?nE�E�} ]��g?a��ʞ���L���*��y/���X%2D
r�/�����3�@���hN@!�*��������0���#�dQ8Pt�ҹ&~�ey��~���p;A���$�O��O�7�%AJ�p��:�]�}Ό/$���w&������-��/7�5��*J�w�b"I&�����mO��B�\���+�����a��z:H ��t݈�ړg��� ��4H�t�r$�l����ނ�C�3����8z\7�xELҶ��$�6~����BΞ�d�:(�˝Y�-�&�ˇr �e��T�V/��P!N�����R&~��8�=�O0��O%��)�0��qլ�$�n	�&�L������>����2�fM`�K���>��o���B�z�k����>�W�i������-�8��G�O�I�_՛cU��'m+so1p�XjQށv�;��Ų�..CVKu?��""	8�@��If��\-S�L"�=�����FD,�U�,��:(����"��B�
o�)+͠���TU��Z��U:�"��v��a�{�vx�;�w��R��Z=v����s�[2�9��Ww6�Z(@�����!���� yXnb�y�[e�>�=�n%yPW��z!&ٚ'�q�g��,�ݮdz���>#r�)È���F4�W�:�� Gl%��G'`�R�"�r���|��9Ӝ�p��e�N���$Gl�Ipײ�@�s�b��T���V#�Kl(���9���<˙����68�D������ߥSz�"D�ᯭ���1�$��5���1/7�Zk���˅��D��.�,G#>�R���G�[A�a������wM��pX��8�Ϗ��H�f�S ��I��J�PI�����H,&t;
�Ҟ�X~�P�Kx�9/�)[��S�Q�˾)G�c�(8�J
��'���-N�=�����3�����B�9��\��:%B��1��&�WߛJ%:b�̈{;Fw����V44ZnLh���{�i�c�&�����iO9�b}㞘��$U�Y����!-�)竴;�Ղ��a�n�}���a�2iaR���5�Gg[��prl@W�X<2�z��'�|�E:
����E�����EөϜ����!��8^�;]U@�Aջ4��4��M\X."
��dI�}�C"��xI��j�\�X߅��_	�Z�Q��-�~ұBc��I����zV��Z��"��.�U��-F��cm�kb섕�Wk�������1��n:*�)7��l��isxF�\rE�K����ݿ�졏�}��	]0	����^4T�|
��z]9tv���_@�
���P�
6���3��c��̰ �*B�[�H(��)�@�I�:�Y�Y�݃h����6�,�2����BD�#��H�l���b�^^����}b�h!y�Z�\�"4DAq�= E��\��G̹B�wI��	�7��u��8:l]f���$��HD�Q�Rc��VG*�>�1��;�0�c���f�!9*�q' X�͔��aWEK�/!��s�`��d�u����g�o��ҿ(\̊��,ۆ����s�s�F?���b���"OR��<�����Ϸ��E'xK�Z���%Fy<O$�m0���'C���t�����df�oSF�<l"������rf�M�+�2�;}ĭ�ڣ������7�DцM�ngFmĖ!T�B�p��5��Վ��g�$M�d���!�������Hd�~L 5b��{�2/?�6�cX�����P��:jq�������`�@}#o�V�c�<'CG<^���Vړ�LR+����K�����v��\:��@}
���ػC� ����U-�n&|�Xlv�39��,�5���so�Z��1��x2��y��U�Ma�sU�?>��n�%zn����Q����Bͫ����4�-��⃚�mV���-�;���Xmˍ9�q-�L>xo���vh @�}�#_�-R`������[�'��%��+��cΐ���{@��R����������R�V"J��J��MI���>�7�*�H�OG��1���w`��q�Ȇ�K�F���m{��8Y[FC�J�x g��g+I/C8����cx����a��O�즺��Yo���'WUP$�O�A�דD(�z�	���9��飜Yf��:��^=!h�>8l�p�h��{L$.N�r����՜K���.~.[{)W�70��.Da*{u����'l�M���57�����Nޏ������%7:H״�eUEUܒ;P?J�i�+����c�}�jdq�h���{?���{(���cJ�@q���1��0T�����=�Ey{d�;������I�ؤ��34:	��8�H��8@5U�ew�0��}��#d^0��#��!�,UP�=d�P>�(o�Df��������FPT�Mv��DG7�yc_�S�a�>?���s��j!��S�T�ȱ��W4a�� �{�PZ��i�[ڍ�	���~=#�6BL��$2���A/���@ƣg�︊�6��7��Z�[��*�X�[�դ~�� Ԍ���=RA�+�"�j��@��֛�?��P:9[�z�qG<��ᣕn��A�7?�Tϝ�&	]��r��KU-9�ekd�4���0<�3T�,4�Ы�
fS@H~\�5ο�V��G
�2��R���v2;}�S��-G�:סT��*Vi��o�tN1Y�C�ǿx�Xl'vzr�����.�,�4�/<��>�x>~�6kֆN2�9e�,���"0�|���{_ P�ʡv�D;�W�L� ��ߠJ�T)7�X
N�G��p������L�}9XǴy��إ�bJARm|�`q�u{T���u��]����9�2�N�:��(�e��W�V���W��97^j"��xzB�݈i>�=�H�(�>������7Ͷ�E6Ȃ�,�)!������>�2��
��6CD��Ga�~ٚp��5?�kEM�f8|W�ߛ�j�JN���4
��'�B<�@��׃���\���R2}����i�S��$|S0�xI�;{X�;�1L���e@��9\(�w?�F��u�dP� ���������Z~�T���v3e�Y�i8n86�C^��*��<0��8{h/>F�Q����h֐ņbG6��@O��P�m	G9̾s�׋=�T�C�Z@z|9�~G�_�:�ϽoW@�ڌP�W`sq��:�H�+������k�nU�95�K#H]y�@S�\��96T�_����>�w����V�����ָ�׻��0l.�0Jw���C@�xY3_:$�h�-�\n���.q5��v�xI:���fyY*�tJ٪)�øY��z��5Uj�HQ)潞����<��k����J?������I \|m|�=-h�������1�<��I���8�z�6i�_�Y�վ�������GL�H���+�kÃ��K^S&X��T�� =��J홫E�)�iQ��F�~i��s� �K;�&���I ����/e���G _��&���ӈ>IJ}t���x|T��s�ι�H�1l:�5N������A���5���?d;=��8���Ad��c%���Fs�O�8�u����p~�-�N�+���2*��J(�{���x�~�-`}=ig���ua�8�cu�^Iv�.j!A�uFA���	B��+�B�\��Q/:.L�G7	;��N� ס_��������o��t3�~6䘘4g^�i(�'V��kvdVN_�Uc~^Dn��{L]�=쏷�M0cK�X����$ �B�q�'�&n2�7����� 2L�h�Z���#����Rh��m@v�,� �\A�����8=�����h
�\-rG�y~v�B�A�T�$j���m�[���u����Ų�E�b�̰�q�<���YC�d���(����ʸl��q���[򺣐�]����0��0p�Jxm#���xTd��l��Ѯ�����z���R�_+#�ރˇ��A<���e$���lV�ҍ"�K�@�YB2oD�	_	�����8:1��0�Q����O��j��|��H#�$k W���4�tU��c��V!*`���0Ҳ��ʴM�����+	�^�W?)�vf�/&����b�f���M��1Y9��$f�INQ�ޱI�C�(Q�ơ���.`���U��A9헐f}<BK錞�����w��� ���K�6�=���E0���L�xL�3�G$sBu\�xo����" ���xͼ�c��^:,9.����0qfE�V|���j�#
mƞy�@�|���h�a�_�*�m�0g��|�(���c��`���}� �АB��p�ů��~���)?E���'�Z�mN�����M��O�!*��d?�
	�>�jl��9��sc��X/�=�{����r�dϷ;T&�؅{��aި���,�y�f�R��X`�� ���?��D%>��l����U �_
V���o�R�e��H�˰g����{U까|��([u��"�0J� Je	��#s^�>�B��z^I������"D��� #6rbq@T�T����� ,�N=�ln:��1
9������@J��rt5�h%
�0��k`ç�yvH@(�N��Ǯ�oɑ��6(�JW���TM:LC���'�9��g�E��B�
%ZMq@ /�T�Ţ�*�i6&�a�a��� +���i��^42���Lq�!�=����55@�#�f�:ų� �R�*v)r�9�XO_FtQP�	\�k&3/4�������}�*����!B,u �I�ӐB�p��ҽ���b�$�zT��Yqޝ�_ݣ��Жo�y��sh ��#�b�B��d#��lҍ����<�菃�����
p��aO ��b�FT9p�21���jo�?�"��)W��ղ����?.�`�B !y��K;w���U1k�[��o�.��]���zf��i���V�\&��~�=�5�0$�G�����B�%���/��<FC�6��=^Eɚ�ӫ^�es��a��[��jY�z�n#M[})ӡ�����gH���U}�nn#'V@X2v�twpP�3��҇���1�H�"]�A��n���B�b��Ppi���u#��bb��D^��n��_�r��-�a��7�����礹���
�(-�JJ���TW�8�^e���"<�f���֔�81jN�R/��w7� P�kH�T��ò}AAcx���I9�����=lo� �X���g(�r'�5��~��=7?�E���*N�u�m�<�X�0��ڸ�Ը��M���K���(6D�M�=5��b(�ٔ(@US���5����K.�JLx%Z��B�e���i����#�Ř�c�نۍ�P��@Z4ob ����sA�1��U�� �V��nK��Ų�m>����Ԡ[��~�-���CRES(�19>֨|%��"@�X�«�I���nv��s1��h!,t�r"�qG
V��u�u�0>�V��m^!��r�t�=Fϭ �.5�k1��Dכ�TVAǾ�<��IKEO��$��P�����sy�O����S����w�y.��e�Q�.�Z>ZDf�Z)0�5LO/��%�J��^^�|Wz��|U0����܉��p�m��V#�f\{?�U�7��r�t�SMH�Y���d�6�\�̩u�!�'���-�\��m'۞�~-a?��#��!�������u��p+��/nVZ��w�Q�Wؖ���m������<�}�L���J�s�G[��Bg���^p#�D_�4q:ې`�A��e��O�hVl���0�>�I�ЫFV|������~��l�ͅ��a��k���/l�����>O�k�y��\���O�$����B�i����2|����3���F���Cͣ���Sr[����tC݀�x�ӥ�i߯})��i^�_�솸�S��(b�6Ip��N;`��E�_-�΁�l;�;D�=0���)��7_��kJ7L��rsI�ܸqD���� 9Ib0��=�#�������Q��S�F�� A��*H� �:swT����<$��|%lTԗk��ޘ�����jT�;oV����T��i�JZ�,1J������L<�ПΞ��=�O,��KK,�Ǝ�e `$�y�ª?1`���t�����~� +KT3�������S�16�L�6�������.i�#�rġ�t��ku�^8d&Mٜ^ *���q�@��P�U�֐�~�J�1N 8T�WT�{��X�%�0��? 1.�+��m�%v4�<�LE�"�j��Zc�X ֨�]cji�B�A)i3�=����m�`#1�,�UD�R	d(�6�R�x�i񟸔(�5�"7;l���f�{U�ɬ���hS���&KR��|���J����>�i,�T[�D�7#
�0�������~ux��
κŖԍ�d˪�F���a1r:qP�ß0!��_�WF�h�U%�[�4T�E�9�ӓ@Ȁ�s�!�\�5�v����|�DJ{d��<O@�k�=�;��y]��su_D���ѣ�07�������0�}'�e�{b.yTp��]�Ɍ�!��6��4���S�
��b����2W.c���(_C���$�s��H��f�>�Uy�T����A��X���#�%a�B3Eqߐ�|�w�3~9�'cg0I������EUKM4���P���Z�����k�j�F^=�~U�����?3o�<i2����J�)?�O!; :&1�)�UI�G{��#ތN�U��n�ý�R]�2ô�#�)]�F�_V��h�%ȘdLD�wIp�Qe��N �]�ZH���F�&�Z�O��b�ݔ��
��?��t�
�5���$���2KJ��A��C���Y�ۦ��J�x�Su�q�/�#�EwE�	//�s�rb!צ����E��33���v�,�}O��}B��c{�fA��Υzd�Y$�L�r�=:u��q���q����MԵ�Ħ�/32�����u��M_PX�#��T�Y�!�����'j�]e��G������edgZ�mYH�(��y�{���ïd�;�	c�B�9L����ݵ�89ٴź��k�@d*���B j���U?�ýv��dQB�A��	;�d�i�#�o#~�D�7fzܔ��^��ܒ�y�n��3��U1����'�: P�i;[�������!`����"\�s��b�m^��F���"�4����S�`W��:3�7�]�
�qnW�I�����J��􌦞č��H�FP�OF*�ݩ�Zcm^����[D��B�z�d�f�#��'3't�
�J��B�A+CP����|;���+�Nb������$i��̭���~m��Zz�őY�� @CA�t^��-1�Pc�/��dWt>��7�xR��$��G[j�h|`Y�$����߄I��)a^�oc!��G��_ C�mH�cm�:��1y:1��Z���1��Q�M��3 ^���Feӯ�fSVB�Gw�ل� �����Z
=jΟn����s��0�Rr�X!�x�]Q�C����"e�{5����,	)�uI!�tޛ�T��00�.�}��Q������(��!��e~�G�ݛ~�a����^gJ�:�ƞ��N��a��🸱8~U��1��3��0�*�Ⴠ���䭜-h�8��R���[�e[��f3��h�J�}*F��X�0�4��A)���]���f��¡WaN?*�1�=�mu�U+�ݸ-2���� ���j��^J�_5�7ʍ�t�n
�tBP~A��׹l���xx�90h��hƛЂe��G�{��s�:��%�+l���%�Ӡ�$ZA�H2��i��#�nӴ"}�]>�xN�4����>����N'�v0".i�sC�[�ٝ�U��p�����[9�I3�F�ۺ��ɲx�"Qf���m����Xb-�������D�5��J��Z��}v�7�Ǫa[�����=��be��<��������4��u(�`=�ǋ.|��1��+3�,�~��%%��v&]礍��?�	9�;���J _�~x�
u��B?O�y���d>���h��S�㓛 �T�ߖ���R���M��נ��W��l�1c��n�)*2c�=�b�cN5{���D$UE����ӏ'��}jR�B��,Nn^%���ݳr�W����p�%�	�ya�c��`�=vG~e�6�x�@�h�$�O��g�;��,@�^��R�`_}����lC���������p#O^v��k_�iϒ�����0�i�h���M��2^��ذ�qJ���*)��n W���s���tOmlc����35՗*���u@S;�bJ�5L�ѡ߮-W�c��X���W��%k��Ia���^��������u�yVD�	ds
�d��]���>K�	j;�(���歸,1U�c⪢Yh>lM���I��a\�C��}p���C;�d%��/���a��z���H�2��Wi�Kc��@�k���)�g�p� {?���ƣ���@-k6!����L&ߜ�.)5	�I��8�eRr�ob�S��� J���Y�%8U1wg�s��X"҃�uvܾ%Ք�"���f|��滜���f��5���{��O�݉�� �T�*br���dN\!��v�&$�)ckj_�fx����PT���R�*h�9T��R�S&���`[��K���{�^���?���N7�x,�k��8��D�{Ķ0�-��tG��Z��ߦ��v��K��"ߧ�
S�O4|#�����̈���+�'<�W;6[��X�MJl����DJS��u:�DαqhZ,�q�B�=��E��qߖ�ޅ
r�)0�i�j�L_O�3��E��a��+KQ;^c������K��������6ܢ�[Hh�_���莼����wԳJqzhL��4i$!ނ&���lR�f,?3�[i�@4�J��u��ݛb�.�����.�g�&�+%�p���QIF�Iy3ħ������3&)N"N>��(u�e-P�!��j3M��r��N�peC�u��!���Mב���J{abކƢ�z#h*f���!�N�_�B���6rj�*^�J�ܔ���jx�H�ڱ#����u��drlִ����U�w<�3�w҅r�)�UB�J��8�P8�B���1T��T�5�C!q�ȮD�x�,a�w���m�bD��{C�ɟ�k�lӓ��XlS���^��	��2��?[Ć���>m��S��x�rLξ-2�*�J(��`�J���7ǹ�e�(W�ۿu���]	�0R��Iఛ<!Ɛ8�`����\4�c� k�G���He��m�7�W��ғ�zk[�k��CǓ��2�u�dd:q���B[ �#;�F����(�f̍�Q˅�8���K��;��[ױ[��Qs*��}D�˝k>&8�3[��?��4>�����W��p{Xsd4t�v=��}�{�Ѽ�nk|YcV���<��ú`�g���Bt��C��Q����	&�@�GEps���-N���"��i��K|b�s���K��ELYH�y�#�3�`j�9Ș�U��J��;����"����RM$Iʤ��l�i%\%t���
�P���Ln�^k��2d�$�$�]���xF=��(��YmFr�HWɥ
q<k�M�p���Ê#C�=�2c�B������m��#��w|�Y���{����|W"s�1ݐi��i�jg2i�$ʐV�ܥ%F�����{���J�VP@Sh�c�<:w-O�ob��@�~�����;�݌��"t��#�R���s�<afP������Y�`pZ/+6��O6�0Xh�M�>����B�����Kɋ!65�)P��0�&&ř^�i��a�ءU��X7��3���=�xAeJ!����ҝe��}<5a9J_i4��m�ѓ�[]�4���3�b�ુzH��C�63��*ǻ�� y���ꑮ7L@�Ws
�:�~���&���I§<-�` �f+��Dw�x�d��n+��2�����)瞖��*��By��X�(I�Np��@z����RAl�dLDϯX[{
yT���.�c�n�<��&���I�ߨ_��M��r8q��'>��]���`@7��W�U���{|�X��t��4r�èDdi�k�rP����آ|�p���?�hB|�3�C�?�3u	����Zx5�S��$�yNO���$U(�H#"z��y�X���wtd�z�wz����7!��tx]B�I$GX�zr��x-]�\��ce��`�I�h~�1]'�vq70ʊ;V /�VE\,�:��;�Ra-����)SX֜�˴�;kQ#��x}hɸkYa� �*?��Ro,�`,���]9�kC�U�����0fFp
��~@]c��S�5��,��)�hr�������g��L/�Ox�L�6����5Q�� ��gTDg�1�1�p�����)�xO�{���Y�
)U��UPÌ�qJ���*�Q�|n�����}i���@0��&ǩ����܀Lf�WВR��ᵝ��cb�I�2�����I
�~,U�}p�w'W)��Tv�̼�o�tp�Jv>�c������+[�'�Q�1�S���)���Vt:cU^����!#��b��g�'�I�wh!��!�l<p�Mw$�9[�b���g)�HoM�z �p����%zQd�z˾��(�]��RU0��r|y��(��WN�f�i��=�y�AMB��ڝp�;n�|��i�	2jh�%���J>q�q�wg��k��t@Z��JO2���k�K���H�^���VT	��Q��!�\����iZP▤�����������bx�@�/��U�;n��׭#�'ݝ�jkI)���9�3t�;����GH}�������q[,�::���SG�P w����H��=��T����fW���S�~���Z���ڕ��49.��v�q��aS�S4�9o�̉2���mU(�ڷ{_G�P����gиT|� �U�������|Om<���Mu#oA-u_�w��� ^�~|m!��x�V��#⻱�Q�u��v �1/b)E}k��݀����8�
k��z��iV�E���g��Ԯo|	=(e�dn�b�S�9�mT"�[��Q��	��.� ��ճ�ib �z�q6��=���:�����e����˕�>#IT��ѭ��mX��AĺF��k��\X����	ڳ�r�v� т���
�$�0������������l'৏���զ��h��\��k�r���a��>&J�e��.�1fX�As�﫼-�s��B�$w攠1	~:7ǎ~T�ĺ��L�˲�|�>R����j����H�r��A^C4�=�{����n�P����x��峐`f�1�H�ŉhQ��N[ �>�>iؑ30.��ub����LtH��ܘ~�9��	A�ްyཟ�V�lmL\f$=)0�[�].�}WL��..�Z9��5	�g����|��0�1�Y�|ۂ�¸���[���(�]u�U5'��v)�j�������������wr��
"�kg4#Rv�����9ڵNz���󚾡��\Y�%n�N�ivq.�߇i�S=
�O���4�
�KI��V���̦�&3�}ߨ�j���(N�[{�[�=���r�?L@����B�9��	D��{ab+����u���*�NOt��A��D�������ݽ���I]��Du��B��4) !�>'A��l@���,���L�S�k�w�Z�?����*D��=����ZG�����v�3-L�7���~�?ǐ �n%<=
�H�>�+U��p��c��f��F?�dզp������q��F�$Ÿ�'�ͺ�Ԗ�>�vi���t�8��M�N��U1�J;�*&����3��!�q�����ʹ���ň�b��N�v�ѯt3LH�G�wQg \
�B/Z���F��*�e�VYՍ��g�5m�xO�����A�V�J��Y���Q2my�(�"8�ؐ�頹4>�詻�_h�3Q��Vű�������H���|��gr�@�0�m�u�\^*.��4X ��?����^:.�SpXEh���i��|����_���݆���k�$:�ٮ�B�¿c���b����*p�f'/��n��!)��)�@Tw�˩bwo���?(�.�ۀH5J=��v�?ss8����q���7ƍ����i�	t�B�~*�;��,L���g�Xk27�س"dQ��� <���-�S��0 ��;�n��b�-�Ll7߰>:��X��}P��fv� )���pE�)�*y4��va]�d�Y>����	{����;v��	8� ��=��!ra�M�׻(m�;4��-ri�T5��̳v��Eo&_���|,��\xeVB�������_�X�����(xj�,=�Kx��^�'�#�|Q�,J�~�X�O�~��H��i�2��e`�X@x1���sV��2��Q \Q�����մ��L��ðX	�8���)�i!$B˱[5;�<E1[�\,���N����s��a��X�űTv�ΣX(��ִ�H);�+�;����z����A�!���$�Y�_u�SY��0`th�XQ&����ّ�Nc�Cc�i���8�<}�=VP6p�A� &�J�9A��d����J�0Ǩ�U��f�<p�g�O{8��	#�n���0�c�g~��r;2&�i��IF
o�`f�$k-��v!�b������ݢ���M�F�������>'�K�o��Z,���'��������l�N����*�I�k:)J�[�.v��僾BM¹$:%��Rmg� 4#�.�11v%2��_�w��3_D�n}G9�Q��F;գdK�a��G�ٿn.
�P+f�w1�ug�w���\������R�d��T��|`��Q��w=�k��T8���*��a�IPѶ^�����]ٖ���F4�uRTtEo����!h�6'�bu�/刕�y'HO�$��д���G�ym�*"m��)h���q�}pa�B
Gs������ ���e�:+����uw��U��[V�4S�q��S�*�D��cKr�ײ6�kI33N��o J[�[��!ғ@5��L����a�h��t��)��'y�3��\�Fn���l��[/_�?��cP'E�-uJ�f�p�`KM�<(�7�Vw���,�D�W|�er�J��~P���h��j�
vVY��>0�1)2�T��/��)M����g�;Ԏ>�u)F��-+�Oz�=��"�<>y��V�~��x�Z����^Mג\O#�5�uR�CT9G:dv��q˷�q�K��NU2������\��^K�1��}U{�>�������^�a߉�����2��9�L��)� �F�6��L�j+�:'�HD�&���ٍ��7���	���j�u��a���0pG�l�ΏcR�n�B��`Հ�t�}\xa.o�d���@	��#dgnZ���竆z�o$*� �6����|W� )�V�W�� @�ލP��C����_���#���P�PLӠzeb)Q�10��v��4��՝V#�Qt��)��v�q�LF���GƔ�'זʕһ�_f�f��E��5cIC��;@�ssJ�S����Z]��0⃂ 2�6 �{��;�Y�2A3R��5g��Od6�lg1�16Z��%U���{�-J����v��lN��3�8E�E*���չe��#�~{�/3d$��ܧl����gd�#$�tfѹ'���t���X_���)�4.���h̥��0B��mX!��Tlt��0��'DJ�]�HZc�8q����LKc�G Z��U2:E6FnP�1>��j�~�7P�)g��0���ps��$+Q�����fiFǝ(�!��Ŭ`ͷ�2ZYF�I���X�!k�z��m��x�&�{W���J�9[����+ɵ��f)1����?�d�Q7�O�R!��"��;-����fLl�Iut�H�lܒ���V�;�y����i�s����)�'cq+�a8H]
��9IR���Qb�6z@�M)��M����˂J�����)�;�D,_�G�
���I�-:A8J��Yd;~zOk��n�,#f��wHƬPE�F���f�.�ð[,�)���}B�������LPh�z���/+C=kn�ɚ*�D���&V��>��z)*��"���)H}��X���,�9�*9J������mk�gYO��#�n�ݠKB��&�1=�b��ͷ
f&8�P�,�A��_�H��aO��ri���
�@l���,7B�����j1��3�b�ĺ[��*�����;�6UA(��`�)4^�F��bX"��@?�"g	��鈻��^�/�L��p�# ��x�R��i	����m�dB�k�mZ�n��(�ϫ�{��'m����58�M�8vp�0G���3�D���7�]E�/X��Z��{�ƆT�x��p��M�� GJp~F�EVV�;��3H��U�}:(x!��@����!�=�E���2+��-���?W�NK�Ԭa�S��}��hÚ"�Sq���$M D�OJd��-Nߘ����L>�Π+Tm���\�&so�"ہ��	��9އ�|��5�/eZt�	U�������M�M�|�)���d�w 9�"}N�H�0�`9m��vE��E�񱬆W�tA�����O��4	 �و�Bey
�4	VV�LL�9mO�Y��p�H��n��`�Q�u1���Y��ʪ}7��͓[R�*�x�CpῚ�l��k�p��`�N��ҭ>��羈6s3�4d���u��І�W�RdK2��TS3y��s�b?����`	��+;b��N$����Y{�F�x;�<�F^�-q�jj��r��H�h�i����	�!���l��h���.�(BG�ESc~l\�$>�KP�uEqe�Z��{�[c��`;��M�� �}	��Zo��tD�g��D�����Tj(�Vݽy�Z��Wu4�+��]M�1�ٺ�1/��Nێ�z`6�&����2W'_B��9wsyf�
޲���P[�"��Z���<1�\۫�69T�'ĥS�9V?��B-�]'�yZ��C����ryv��Vq�'�,����K�K��()L�/$�>;zx���
�wD���S�L�4�r#E��r���c&n-��8�e�S�ㄺ��0�82c�ð�)u>T�mE	���91V,oYR�삎2�b����A��޳:`���	�N���F$~h?1S��e��T��HD��5��!ϣb���'�6�ڳ�1�������ip�c�+���Hz�RQk����f��/��� a8<��$��2l�`9R�R0���0�������w7��
�x$�~�u�V�H_*���3k����b�.�s�^�-L����)E�E\P1ğ"I+F\m���{�C
���9V!�A�{�0��Q�W�w�vbɏP{�����z�o�F%xGU>h�h���2��ي/=3t��0�m�����X��v`.
��>���d��%�~�s��B���#r���E�����3�pݶ-}`�%%H�O�N��wa��lМׇ$�1� h�t9���p�k�o�)�~�	>�G�c�o;��@M����jU�u+M�릶��҇��)�!��+k�8v�/5� �K.QLEOP�峈Z!f)��<C�|�,{�?OqXM{F�F�B,4MI��
ٮU�6���>$U�r&�OF�����g9��P^�Y���y��T���Ԅ*7���qF��2M2��5�^�����\ږ3v�@����i��(��N��sfN�5٪�و%[��(��&��]���bC�-6�T��R��o[�����\��^�;��L���Л�&��<>�����2���i�F��8�i&;� ?^�"��������證�j�0uQC�Z-	=Y2�]Vύ��5q�\ o�%I�Y`��a���=��
�R���NA8�7�a1\@F��A�cӟ�RdX�^��b��j��y�"'���aD����O�eu/�b�ak�ĉ�I�&I)�	BuX|}��{2_�$/�����)u�yay�Cy����m��80)dc��$O[A�GU���!���K�
̢��BLX��L�����qfj�5� <�ɉuT�� �^`��Ss�
��}^2�gҺM �I�\CyE���顟rʻ$���qֱ�$����5
�U��R:��%q��J�z�{!#���OԏҒ�,�x�J�b?�	��f��U� �.�%A|���?��E�D���U���H�o�1L���s��Y�g�~z���7:f��cv�����J3N����� *:�󍙁��Jw��ϣ�'�ߥ�h@�Wt�/�ŧ0�nd�iW�ϸI�s�Z�@����{ZE/?�� ϭ:\x̴����.���я	-��{��X�+��u�O�9S��.|�k)ϵc���Hɬ�Y�	�Ȁ�
�}���xٕ�=ȱG��-g��)�y&ۄ�]����X��ilnD;�	A]�*���_[R�3
�>�d�����ײs|�V����׆�ό��af+^���K�.�l�p��l�eE������j���p��?qh�-O�?�ax=
s��fϷ-�� g����&iġ51�-���U� A�N  fd���E��Ï�w�@2[�y��py첗�Z@n��k�������bY79�SU�t��K�R���þ��O*سvF/�����id��� ���Rz�"� �_
��#�V�\��r�>O���ɿL��i��3B砖��(���)���lQ���qS8��z�q�����w1��iٓ��<�N3fհ���
hg�ߓ�X��R˕h�I��6�Cg&5b��i���<��H]Z�G���)
�=�c��J<,<�H��C)�v�[ء�o+^=�MU�������;îv�t�,n ������l����w~�,�<�ׂ��X���nsx~�������5i�&V�Rv���y��P�y�uZ(b!xx�'wg�����2G����f	'
|����0EE/���W�"����%*�RJ����~�t�}�d���A�Z+E�ǋu�?!s!v�2��T� �D��K�b���Q��P��E1�Yu�wD̛��PД�+c.|� ��r£	p:����%���7t��a�Ő�r�82���#�Es$Kj.U�h���4�� ���l~x.>.�d�\�C��)�����F����%�a������`3;�H�>��O��#�$b�cO#3��Kf�ױ�.Wy��2i�Z�дڲ�����։��^��R�=�v᯲Ֆ+�F�?L��/�_�=;y�Z,Eŀ������W4��
*��f��4�U���B#������c��fR��!|-���J�{�ɪ�.������F�,��|�����/���L���S
ˬ@�0�_�z��P5FGf����M;��0��#���n�n�ⱇ�w�\0pe��Q�O��F���1����%Z3�C�T���<( َ�+�+�6�4�X�ɭ�)�\�ɺ� TW��6��,K�z�ﺘ�8������Y�1�P�$\���bc��7Ƕ.� ���1dО��ڗRV�"�k�f�_�X�4���9�����'�.
d�-ŋA�|��n�ܚ�8�!:M��D=iOQa�a�՛�,�xP|hP�'j�o.�>�����XJ�0�_�p�Pm�3���^ ����V��2�{!���1��ĝy]���f:0�M�"�`T3v|��?K~;MI�'��af��!�*yr��/��וH���k�Ҁ��m_�$	����F{�*���~�`�":,c����M�ߎ&VB�A�6�}���M/a�n��[0[u+kj��af}��a?~��!x��󾕐�c?D�.�!���`D����H�����4N��t{��\�͗�0ϒ��0���nT{���tŌU������U���(���/�}^�Y���a�Q����;*�dKڷ�����Ԥ$�C9?����<p2x+&��zai77�e�puP�����\����dU(��F{6}�Y
S�O,9�.��iꦼJԛ�w`IU[)��D�7�7��4�d"������B��q0�\��ݳ���B<�B>��ӞP��#{} ����/��dQص�X�a!BC壘�h���ċ�f���J-k%��XbjU��S�-MϜ��ư�)uUo�^��&B5|�$�W��ao8�>Yy�)��s�w�L��8xV�:m��_b(�V�I��U5��0��mu�,z}�� �q���t~��?g]�O<��u��v|@H��ϴ�.z&I�����A����j�ZX���!�q��ە=� �ஃ�w�L�ж�I���&\'��u�tҵ*�1uk,���yۖn������ѩ�lW��3t�ʵn��eO�3����K7���O�;�	��I�����?�y..�l:OF�
_�Ћ�5Z^��n`�A���2y�۸K{���SP����^�O��d����+"Y����Ybl�^E[r9�ǐ�_�xI^�,��Р*?q��>f[dQڬ�I0Fj��@�7}$CZJ�0�	�1mI�S&�*1�H��)��4�t4��k2��1���eW̫�ӟ�(��1�b���b�N���}CT����g����JZ@�7�q*�CAZC5�	o*׸Ŷ�Nd���@X����!��a,�����e�*w�t��z��k�M��3�@�5��R;-5��Z�~)�Ĥm�	��ɷJ���
U��m�/jK'��P/^�I��&��C8|4߬��^*W/�g6c��47���/��Q����|�|$���)D6I7��zQ�u��?kay�]�-o@�#?D>���}��є�ζ��a��"�A���,į�(�Е�� 
^CFѭ�?���ѓ>w��xE�CE�������[
�7����*f��g�.ׁ�D��K���ǹ($�9-T�`�ל�[ZP�}��]?X�y��&��?���8;{�1�1!���I!�H��v�3�F%�X�>P8oҁ�#	�7�A���N�o�Eϧ�WyN���V��bϿ��h0�t�B����F�Vb3�2XY࿖��4�}찏����j4<��[b���%�*��)�=w�	���Sߕ�S���������֦��&#�&�F?i�<A.�X8K	��JKe�'��v.�ki�ՙV��(��PƼEI��LH.j.=cG����aR�3\s������;�M�����U��di|�?���yk�/�Ac��'ׅNE��$�6԰���t3}1�@Hd��lŗ�8���Ə�։&����y����v OA}��8!r[t� ��j�������{ⷵ��]�]��z��VQ��Ԩiխ
3c�˪��Z�|����L��; �]2��>��<l����o3�u~J�H�M�dK�-�{
Yf�y|�e������}mH�]T�OP
��HQM��L���Tt����>Lo�N�y4��N�
=�%�}�=,x�0���:��s��_)�T�����ѬH�C����-�e��"S(S�>��'�����vYI4��3��������K�J⽌�\�k+ϱ�B��e������-. aך8����v���$~�- 6�)�]��K
N
[�ɨ�h�@���W,�p�4���ߟ�0�VQ�ƍH~?�Њ��7N�H�tԴf�㈏g��O��<o^{
 ��܂�1W��<@��]�o��~$��
�&03�A0k)�n�����$��b�}�}O"�T�ը�0�/|k}�����pJ���8���.b^��e��i�<�5���W�M�3X��@ ���	��Y�[E�&M�-`������n3�o�ؘ��5t��XN��1��i�T|�s�5�{��Қ�d�avs�*��e��N���F@�*��l�Ѥ���?��X_��z%	��Q���!߀���?| �MI+ ���J�*��er�cSC�׶��
�}K��6���p_G���4�Q�ڶ�}��?���l��ʌE-"[˩G�eR|Νʙ`�J�טxT�φˮr�"]^���t�/\�2y��B�^�8�퉝���8�Lt�U�,cv�oD;�2�x^]��>_�Z�Xe3T�C3tW��ǁ�����.�E?=T'o��j{�]z�}�Gͼ�v~�N�K[|�ب(k��y���舂~�]vm�b���٦��#��0�M�X�y�?tW�iBon��Νqv-��O�G|�'f'�*�j�Ļ�A�T�IU!^)�?����������]ޛ.����ݡ�����
�b��6VV��`����H*� ��Ҫ׿�_�����{�`�5W�w�|֪�IU��ӁP�}�y�|	�>�����e���.AIBNK�<�HR�spq���l�p�B�������H�Z�tͺ�@R��7���8�i����LYbE�G8U��tt1���S�֯����<!-�j���k�e���.~8�r]O���^�)o׮��"�&���x�[�E���B��M4Z:B��s�r/KsG���c-�p/b�i���-a�k>Ɯ)p�~���V�ci��R��:pm���	B��V�/�?.���9pW����>!
�zo�>��B�j�1-���t�sQ>Q9��<)�Ȍz�_�j��0�M�'�>�l���d�v�R�cc��t�ٽ��S��W�����6d��,�&���=xF5���=e :�Fʂd(��̃"w�$��g'p���Q;G�� ���-}L�������J�n�a[Zk��%C_�,z8N��)�[EBT5j�x�U���y���?���������P��$A���w4"�f��JC�)�gxH4���RHT��=��|Ij���4�;��^Ԁ�GTN�l�Gdab��q�`��a �)mR`��̱fϺ��*�?g荩;�=2x�x�`�p�r��F�3���N�	�JBS�e��(�2k�Үz�?�ؽ�V��"��ꙑ�����ܩ��-��t�d\���Nx�����6�?�� �f�Fߥ�" kD1�ܠ�����z�.Z�<]�n����� 3;/F�<g�L4�N8Q;&��/4�����O�s5��;�����O&b�ȅ��!�nm�[m�g�-���35l=v��R'!|�~�4�|a(�����d�ڲ˜�K�����>���{��Uju��J�$e��� ��!6�ܱ�|~�?��T��1ٷ����������8��`��Uܵ�k����@;�N����X08��Q�3i�#�rM!��x
N�<��ͨ�\Q�X
Xf��'0��90��_���6C}fd��!��6Ĵ��i� �xG�6��/���p�!A-���+d�s�	��f��A�"	urI)��v�N�U8��f�2H� ����8o������f� ������')��6s�n
 Pz���i�p�,.���͢��r�+͟�Zߨ�����<�g,`���W3َ����l' x�QE�cx`Pb� 9���#�)�P�GY��bZ۴̠����l���r�����d��/~��|~nI'��Hږ;3�i�8~ .A(�l�H(`q�� ��"2�$�P�ʺ�Dh��X�mk�o�cT�6 ������8n���3��*�G��0k>�j(;e!sEO<䨄�dRU`eX��5<>���%Qϴ-��g0������#9g�p��p��r5y>�D[t=�n2�ԯ��+Q�Z��W��Z �21gv}0��?�b̞���q[Ʌ�w�׼C�1OT��$t%|\R#�n��+x{LQ��dg��x�� ��	��)�v��)�u��#�Tɀ����f����y��w�r�T���Q��� �lB�ጞҫV�,�'6���Q��%�,o�-|��n괙f�3���u~�F��0�H.(l�ל)y�ķ��1@�b9�4M1\�.0nj��I\K7�,�+6�`��\BNKy��!�`.���ޱ8���y}�J��cB|��v���r�{����#�ћi�ʾE�;Rj�Qˊ��}d!r���#%)ꢳ���ɲ���ҀaV��Ģ�v.!޳Cc�4��hB��$���`�'���+6��%f��:�3Z"�YN@{b��ަ�ƹ��<6�M�o,ٯ�Μc�u��Xr���Z�~�נ�PP��5��D�9 �[��2�Q�Z��~�jC���gm&��)����DN�
�zT�dc����E�ɉHZU$K'������-�&��#�y� AE�}J�[��y�0��"�c�Y'u�qC�cto��&����[\gLJ��'�����-����p�:�Iqk��	�Io��z�7��֗���ZvY�<�O{�zA�|�8=���ِU^)�n_/V�3�/$7�3����ϽL��s���TV3�.xmڑI[�8F#�2ɴ0x9aNNFj,6o��5\(*��}��TU�Y#cY����z�"nZ'B~�{i�q)A���M���1�rB?�p�D&|Y.��.��i' |��2�����ƈ3���:ͦ���4@`Wx!]0��ŏ%\Ҙ��bQ��N�X��#7Y�6e=d�++L�<�$6�o�kQ:h`-J�#/�ۖc$(�^�h=a�ܹ%�y�k�;�����o��Z���\2���H��������<%�f�c�撧qS��'�o���5,�,q<�W�7�ay��$��޿�_�^��^�D�l�}��鐚��b�AIg���/�,c��������zČoS~/p:!�#�E'�r�X���.	�jJI�?�(�>k�L�-�*�9HM�_mYѼ�~�**����� �?�����q�Dþ{��A%�t��5���C���E���HlP"x>E��m�Y�A����Q����lB^Wo� � 8dC�P "��_��8W��޵~��P�!5BՄA|F�1�.O�U�$Xg,!-��l��@O��+~q��u�r��MN�^Ve�F@�I�ƻ�03� vXmw�,p�~m{��<3W��$�z|yQߍ���_Z0wLȨ�XmX^Mo��D��+|���^8R~�b�9C=~�cH�ߝ&:W�����h
5�m6�~�a��&�B��{��5�?u^u�#�-Jۭ�.e�z14?(���#�	�5B��0��,�$�3M�7��LY.՗���ЭG��5��B�vȷ���#>������i�lg�Q�4�?]m��ه<,�Fr^��cm�MBO��W3:wVp�}��f6~�*,B�}�9�;@�l>�|��p���m�tP3~�B�7�7'^�F7T-��U�.5>��י��*�iX7�<���(����|���S�8g�i-��cWtE��A�,j������<?�A�[�u�G��/�09Xf���(NWr��}Jvv\�0�*Pn:�ő��B�.l�8�TV������*���->�X;���)r)���O��+_�f��*>��{�v���Fd���B��[��; sk���/�TԞ���ׇG���/@�-��7�<~�����t+?�Y� C�Þ���>���\��*Q�I�:[�'uS �Џ��놨[o�OG���]T�3���p��-�[����a~��p<�R���K�<9��W>{�L!�K��>�r�:�� ℭt�Y	u�+��`��]�. �Oj���<&e8��Ss�a1�S-� �)�FR��5c����yLO�i��7g�a�7�@�u��6n�}�0������^��=g���[� d�h��V��1�����i��I����IF =���%W��O���m��'�}U\H��ݔ�"~Y��}��5Q��iS��*�4
+�jT/���HN50o�	�6v���!�'�/m�,��X,o������*+h���6����!�j⼊F)IX��"i&Y�+���gDB�bWu���0U&Ŕ���Q�����6���wY�7��E�$����P��xz��fۅX���=Y�IQ pY�߼*���1�5l����cP���U9��r`�5V>սE��G�Puܪy�|�e�%�;�#���Za��V:X:�u_��@�ͽ�Na*�%���|[�> g8<��a�����Vmtȑ�Ҏ!x��b��%{�zDDJ����ej�*�z�ˮ��kv���B���l��7�'"˨E��~<�V�^���bb8��bl1�s�`k����6%��YtoT�!=&T)125H�{`�A���K��K���zX�p������<z���J�B�]��&�lZ�������':������%���k���T�)�� b��;��Q�#�汭���o ��Բ��M�
��.o'�J@b�A�.m��@4����q�������C!�%��5��$��=O�F��' /�F�'X��ePϭQ�S˟��H��Հ�%	D�	�g�L�r5no}/�R�����ȃK�,qT�Xj����?e	�"R�0�]���`���jblʖ��z�dv���Dօ�T�N)�֞���޾
V�"I	�G�Q���63�t��"����¹��gs~]���/
���>a��l��dPv檒dS�pn��ڄߔ����p�n0������q?�V��3��1�6�F�Ns�[?��08��L5�;�solD������*m����7��Z/�ZQ�Z6��5oiU�$SR7�v�}��ɛ�� ���F=[oJ ��lfbp��.�׬��G4�����d�U&yvS蚖f����vW{�x�$�@��S�0����-��1?o�T��<�%�go�U<�K~=�p$k�ǰjà�(3�5d۶��z^���K�������������#X��*�v'p�)�#�zR�=�$$ڤ����*h@�h�ݳ� ���၄]�J�
�/,��<�;&�I��z]B�>K7���Мfy;�Z+p�Jo��X�)vyMky���M��`9}MblTQ�j�D�� >��]R�2W�f��~~��i��t�h5�3B������O+H�^W�����Y�j���ҷ�/M;����f��M�,�q̣95������) ��"e2�@$P?� DWl�H׷$�:R�}H�V��_��x�#�O�k�C���}���`�2`Wt3��K������9�;9�����jmhS�������-GSE?�j@��%��V�x��.��n��}�G�f9�֒��!Ka*n7X2y�,~�� �,DC�k��G��d��Ƙk� Y�9���򁸞�$E��>�������X����$�Zf��.C�bA$Q�E�7�a�vcdH�����@��`v� �h�4��$���,�[���c�(\��P=I%� �DNq��l�_i�]�KΙt�	v�E $�X���_4���-Y���sN�����̎�ȯ��m+��A̹n�B�f0��7�^j��*��gl-ܚ%�8�?��<^B��'��cF�9��H����*����)\�k��R�U�9��V��H���,@c\��]����6�!���)�8��6�xd���vV[>��X�_����y�ΔZ�0�w���D=�k𣛼a����уɷ�У�<��'H|��5�L�L]���Q�
J%GPdel8���ڈ���D����!
๲T�ȼ�����h��c8 G�p]u��t%��--��M��Y��`.ni��e�;��9����8Sb�g��/��C`j8a�\ /�Gh�['9����m��` »�T��ߪH{�
��1<H��b(�t*몞1nS�x���I0�oJ~��r֍��Cb�Wdpqp$0�O�!
m9�+�x��H:}�v\ե͜wp��Lr*��	�����u�oZ$���gn���}P����[h取��*����p�?�({Y�Iy�6���¾'��́e@��z*�0 PI�/83[�ǟz�ܫ�5p�,�e�i��F�~+�c�IB�$���+O�J�E�z`�~��fLe�z� B{C윖�y�2Ƈs^��dF��~����N>������Z�:�,GV	Z�� �E�2�������%�ߕe��%����~�!1%�G�&k��'�Y�D,HD���)��U#�)4R��[�w�~ _�۰��(�-.VF倰������;����'� ��@���FrxBk����VT��i���$�'�h�ĸO��$�o6{�(���,T����]�w���r�x�ZmRb#�z��@���@�4�.��\����	g�ҧU?8夵M�J*5"	Nj)�b��s�/%��a�����q����C�M�H�6���t�ᄎo�GU#�[넯w���F�D%�k�sQ`	�[Q��)JrbFR�։�E�j��J6ܗnDlh	Ƈ/�^����є�ݾ�+�}�#��)�D�/Ó3���-�O�`8hn�*72o���MA�h#�&��N�.r�(�[�O~�χe������&}��8I�z�c���.�c��������}2��FX�H�jr��YJE�T�Q�F;����>���o�%���2�-�f�Y�B����urљQ����
����1=Y'����Xm����9�h<ls�9r�G���sW�x��.g��W�˂C��N�����\��ꛏ�p8�0�VS{���"�I�N$l�3�T��L�P���4نf������0��4׶j�M.J�@����)�' X���̾��&Z�w_g��
��h�#S��LӐJ�O��؄;�w�ػx���6�pA��U5��u%�B����%TEC�c��Uk[|2�S�5���CS��z�Վ�Vi���W4ro�^� �z�����E6 F��_�����I�$��@��T־�phK���2�!���;w0�"Pv&Q�ۜ�M�u�2]�y��@z_=�֩������M0���;��HI]
�T&�m��Q�q����Y�8���R��҆�$.����i~<�'|�Pߘ�V��h�d�1O��Z�!|D��L��$A���s�먟?��W.cQ��a>�b��q� i�6�µU��k9�x���ELeT2 L�bu3�$kЅ�
hǖqTu;�-`N����{�ݑ�R�����y(�>�ɼB���O(�B��)�3{&���ښ^Fkd��E�F���}�.O� ����D1I�;��C���Q����c�I�����'�������=N���h���(��Ƣ��Q�/Ղ�Yt
^#b��%8ٖy�~ck��k����ado�k�X�7�P�8�|'�ث�2t>t&���6��X,�_T�{{�(`@Q�,���$mT�(�L{��BGx*_fR{�Tu�)O�צE�K�Q����{��H@��3k���o���ٻ�gw�D��z�@�)ӑ���;�չې��E�Lw�܏[Q�xA�$��fxOZ��b�`����� O�&��R��<;"-����p���^��~-FrI+�6=���?����*��L��YxuxN���O���%PAS�j�ۈt����R ~��K��۵/W��[m��X��q¹N�ă)��E,�����gC${������B%�[�۝���W`=(5�o��4�Yzw��rX/뜘l�	�9\A��*0�a�+S�i숨ع��è2��HI]�Y�"P/�o]ߛ���[hz�-g�©�z�&.�o[��i�)|�n`��\�(^�{�+u,8�cK��`]M��[�� 4 �n��ڢ0��u�aD������pL�6�wT�%����(l
�]tVK)�e���uE��*FP�#��%V+%�^^1%'9��J�}3�u&"�!�W�F=p���"��8Nwk. 3:�m0��5��ч�E���Kpw��"����'s���(֝	��8W���ʢ���:ڶ5�'N����,�CZ�M����"'�i�	!,������h֋X��|Y�\���yo���0��SM(����D�L�?�;�d�H	�S�O��݈ $[X9�-�����$�fج"$Ɨ�qJ����[n�A�砏C�/"���F)���^�#<	8Vc>�duw���T�;&��*n���]𚐯ot��0a�3��Q���Q[�"eS�p�:K�4ٙ5$�p��ˑ��o���?؎��(NA{�8w����N�!��1���Y�ɷt|G�*�)i4�\�̺�|��T�� wW���]5��A���F�A�U2�M0�����3#ꬢ��<��W	��ݹ��r`�����~�jI.��y̭�������P,�k�zH6F�&���q��G��?��|wX�&������O�@�����,^r�2ٱ!d[���N�P  *��Y�:=KgiI�������'̀䁅�\+f�2$�o`O� �#�)�}�>�fv_E��)���)�qep�gR��q��v��"ژ�$I�X�S�DE���a�,ɑ�7k��|�Q���.�AE����Ao�������9%�%���g'���b|r�M�0RA�;�6��$�g�{�4bi�O��j�4�Jʹ �0q7�3,�j�S�vxִOuI=�iz�ř@������\q6�$%�c�D��b�	/��c<xU �C^1D�{_woS!�i3�ar�jy�J=g�.���Ԩ��ǥbE2a�[�k����H�4�|�)�Ҝ�eYi��R�RZDmR�b�Qi�OVe�M��C�l��OtP"�U�1���P�SK�0�s��ݒ����	yڣ[�� 쨯�j��V�-�gę��u�˻އ�o�MJ��q�7���	�YĎ� ��=E��ɲ�P����[
�Fv�O7��3�{��d�8%հ�m,p+�Ϲ �`�$�%�N���"J�����%]�$0F���*q��@@�&= ��uRK�6��?cnœ�����.k爙��Z�&�+��06�~U1�Q��71A�����m6�х
Yp��O��߬Z�_� �"���БyG��,z�/GkXw/k<Dlh�ޠ�TW?��K�1}�r+xm�ղ*2L�$���H�iy�c>�N�6Ntg����Y�/�k
s��b���Z�o�5&��D"q�����ո.ѝuB@�q��k�9��&��2ate��	�ʼHj0"Yg@qu>-[��:*��E娨/#|��-3b �U>2��^�<c!+g�BYI1z��\HO3��iPS��\��҆� �-�60�.`N	=�
�-�V��*ݹ��Xmv��t�*�f�D�:y�t����%�0_���0HH�#���0�P�zݱ�o�\�����=����7Qr�gT���C���m��+��*,݇�;�h\�uPg:���Af�sd��?8R���k������q$J�b.�:=y������U��"p�\~I4 y��1Cm0 �&��-�@P�>����I[���H����w��S�b�Ԯ�&��g�fSk�����Ɂ<�����G������d���j§� Px'����4�R�9K�"�|��B!y�g���6�	���;[�8hM�U<?���hF5K��A��I�r�e a�ؘ`�8���:/��:B���� u%9̎\1��H	�ħ=�����Q���a��B�,S�V���-���݊Rm�ѱUj�ˡ�*��IB�'�Kz	�&���S�|�)�;���`�C��>'w#Y?Z�0��4O��G�����އ��iS��Ԟ��ZE3�/�	�tkh/�o-��T��8l�;Z9R,����iy1`˝��:�7V�sW����%U�,� ��d�߹��{�!��9M��:��I`aכA��K�����Bi�U����-�f:f�l��q��분�;�pα�1a9�6��ř���Df�s�ڌ�DӐ�S^ƿ�.M>�ů�tBhP��ͅ�G�� �ku^��.-�% ����T��G[I�����pc"��o�o�8�����7����[�b�IJ����dĽ�]t�&]�&�q144|��`�����`?V%�V�էT\�HlBej�0��HR�������ƫG�b�j�`�t��шg��	A�>��}��i�c}��DݻCr�3_��9�j�0�͒���##��bh<W�2��%ա�!� �L�Z�{�R�<Z�2�)!�,�}�:���l-��A��6�H��<���$a��{��R�' �q�,&j�|��ҙ$�W�#�7 �S=�4�� ���ֲ��-��c7��M��YZ���F�]�	��B�x� ��L��z�k*�оg����2�lF��z}�EW�4l������P�)HN�1�Zn�S�Pb�l�T��U���X-���b{z�\�ߝ��5;�yP[,����cQp�,��C�Ud��$O�@1�)=�'���n�5BX���ׯ?�ȍZ�@�F����7:���|#>��6� xiM�b��3����[�&�WuP�neJ��y<����7t�rcY,MVx��T�X�	�$ ���YM�")��ѥ9����#��ҟb���Z��ܮY����DF�+c�O�K��h�L��_~���IA�MJ�E�S˝�+���%5�&�r�4�P2`�!М0&����;Y�6E��k�����F��K�p��f ��vb(Jw�N�*���x������n�/Q��C��&*͝n�>wY�W�O9P�G��֍��@xQ�M,��D�wpZkR��װ+���Yw����y�[��$��:�LW^�,�����0*q<Σ5�W����`w�I�{����7��)
�x��!�[������>�1�Ҋ~�&���2�c�-�
$��6X����f��v+e�4)t0D�Ղ~;�G�n�6�dkZa�I*6�fOz�������F�3��xA4����d�����$�0	ﶻ��8g2��؁��)�����ٞ2������:*��a� �H����6��
�gϤ��}�o8�&��M�Ҍ�4�Tw�y�{�b�hu��kb �X�C��Ye�!\X�y���b��]���/�-tP�h�X��1\�?�n�������$���Ɋ�ό99�K9�I��o�c�U����*�0����f��Sr~����:����1�&�׀���� �G�
�p��z������%�4`�t������J5���2�LT��Uz"vT-���c�	Q��I�G�J}k�b��m-�����6x�|� �'�6�aX{1�4�ߟ���Q�ϛHLĭ����|�:UP&�;�B�ǛYܼ-[X�*yV�� Ԇ�ę��g�6�Τ�X�9��^�~z�$C( h��4]�I��z�<ޚ�q'"E7��ۇ�g�?oE���I���1�2�k�p�C�v����~�8��XA���o�S]brAmϑ�#^}�e��u�v��#�*P�l��}��0��˹�n�����7\{R���KPr�����r%Ot0�H��C��es��3����C�)�Ygu��2��mXH6����T�Z�?r����|$b���G -��ٯr��\��@[eA>��v�3�=�ڥN����6���5��}���B���n���'͇��@����c���f�ۅ�6o���h�z����|�sű�\f|���vj�tP]G�$�1��֒ۄ	���D�t{�TIk��2�AG�՟��b�:�޿Dݨj��28|�3��ſ�fɳ�N_T�ki2�V��e�g�Z<����]�@q59�:r�WI�x������<vW�9.�9�^�@��s$fD�*<!�/�v��M�|����9l4��	;"���,�ԭ�7�~:��N�BH�r�2�?��|eP0S<�X��x��+��Ȥd	)v9&��X�q�("م%
��#V6��c�E}��2zc�K����V�	r>����. ~ۥ�)����q���2� ;���Ø@�- Np��$Ϋ7�N���n+�DZЃ�o�l#�E�Q��L�|����x&sX�D����-\s����P�?tl�Gtj*��[����+�������>J5�A�PAȟ���S�½=������	}q�mUP��/�s��|��*3�#�zr�I���?ڮ���L�����)vNY�i���gʜU�_�8�e
��.��R"��' �P���A���/��(k��x����6����G�w��P<�c�����x5%Z��_�15��0Gi�+"?����c�Δo�����=vME���A�C�㙕�?��o��R�ʪ��2�����+�F�^�U�_����}:K'��$�V�Mwi 0�����މ�v�C*q2rGVIe�M��+����Y��2zl-�H�� �8���p���Z���{ 
\�<�D�V�(�&�6�+���h�A�yT�$N�k�G�!��+�m���=�]�#����s�ͭ�60|ܖ� ��6Ҩ�g��F^��]0�zxN�i�'�}�r�hxИ0��L�Q���]#_�����#3�gk���%N��I��{����U��si�@��p8)��̥�q�-��,�ws���Y������Μ� jbx��y6Tҹy���%$�!�6�\ȱ�UK[3E�H�<y,�%�^���-��V�M��I�4$#�z�~�{IKl�@�@c�ɷ!��'Fl�I���C�ۘ�%����7%��.�g�0�)�Ӳ��k�N�
(;@,���!S*�bm9��p�z^Ami4��)�:��K=V;�ìLd�k&���܆{@dd^$��Y�K/��5�Xv�r�G�5�fHI�LWL��o��I,�9�9PP��y�d*�,/�������eT��S��]j�B�N��9������C �.��TA�==l���i��=q*$�|.�f�L�6S�ր�O���̒%AI<�.��g��[BE�w��i���Ʀ�2��6��NW!�W��P\gҵ\�gq�����o�b���<|dYq� ��{u������2@+|���<����uC���Xah����^+�d�6η��ֹ_RP=����m��c(�"-�e�S۩���ʼh�W� l�v��9�ُA��1"��oM�͋�J?���]�Qn�x��ǩ7����#V�u�]��M�z�!M�i�(�%-t����]��l�v.�Ge{���n9���mM�`���f�cȹ3�����nN��ѤC��q�@END�a�����|t*����lzE0X"���|���_n_a�)W�퓄BϙD�8��ÎU/��o�7�#�
�Фn�NP,G�]��%%��<4��x.
��ް��=���U�����$�HUI��,����R�_g�(�Y����I'�e§ ���96J}o�"���:s��[p�P�9���Ep��S?��0+�NX������ ���`��^�9ۡ���K ��9�[��23��F�p+##������0ڱ����A�}P�a6mHV�A �UD/PK�"��"��-A��$����-�"{�Џ��
gO�H��V��k��=����j�����`s�_��ǔr�!�}>�q=A���~׊T�F��#N?s���vL��&Ҕ4�9�(/^X��^C�M�K�3�������������*��z���~Q�ɋ'�L�]��n1�![���x�޲u��uʄ��,N3�~�[qL�Hk�=��OOE�