��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>,M�Kߤ�I�;�b��v;-j�f��-1G)zC�!SRa��<���9��11�)�)�4�.�U��|t��-@3tt�s����}�C��)%^n�素�r]	��Ξ�����-'.Q�R$��
y,���DJ��S[�<Q��ŵ�Y(P~9�אb"V�ｃc\8ض���HOT�����F�G-��%{�xP�,����S���j����V̠O,1(7�*�l�M�eHo�e���˞j�W������k���yzl
T%ĿE�"��-#�Q�F��y�]��,��=ϰ ;g�{nȼ��ZT.�{�	�Au�5�Ic��A�FdW�s��ͤ���	W�$���oy`ޝo��ǧ�jv���uL��A�ʛU���<4BcS��53k��]�bjwz/j[�k|D��5���칵H����Ϩ�:��Zy?���r'Q�eq�q���ˆ���I�IB=�(�f�
A%���<k��ٝ�`I��~@ކɅ�v/�QAr��uFds����n@�f<5s�_�<�&-® ]���Q��.��ܔ�k$�	�2��Х�M�T�2iS�����I������rH�:l���ݽ�d"����~"<��\�2�������������"��*�;qp��cmU
s���Wy܏��% �+.E��	��!$���|���Iʰ���G�sE� x�h�ߙ�"L�m[Ø�0��,�j�(&� ����u��>�4}���{h�y�CM����9GZ2luBL.3f��z�&��z�����31�8�:�B�y�M��{��Q�]E�(5�M8��4J~ހ��⟟$#Aj�3<D���9g2��[�g8���ZģL*ruҏ� ��Z^�� ��{5ܔP��[f��Ѣn�DY���ކF,�<�7��SRÚ��?�M���U�7ce��ӟo���Fj~��p�E���~���� i�p�OA]�[g��p�:ޤ_�,` ˸:p�.��X,'��� ���0h``27f>�u-����P�Iy*$�W��h� {6���!�����d"`��`o��չ2#� emҌ�ٍ�zL@L�����:�(���ᇬ8���(�U��� hM���|��(a��`�����rj���<����"����Är�z!M������ '�ҝ�L��9�c�	W0��ö"3��=�x�� 5�o1 T=����I��x«ol�q<ǁ}����?!w:�؈J�%D�W�;5H�$�s�T�vC`�
�i{2���xן��+��{�a,:vL��V���N�'� ����x�w��P�] ��}�T`��Ǩ���\�H�Ъ�|,RA�#���y�d�
�MpY �V	yk۔�GZK}4�,���~Z�=D�Ό�۽���6�ޣ�K�=/��9�l����U㘔)6'Uc��g0/�����R/��q:;��T�VG�a�Y��Q́&���q��5�i�P� ��	���.^��Z���skJ��C��I�
\ͬ�,��~K�%2�A�59�6�����f�s9����1�w�����G�����yE]9��B�@���]��|wM9�i9=i��;t2ʠ��u �\f����2�`?ۑ��K4̶R*k-bcI����#<��-��y��^�FS��L���[��/�K�[\3�N�����t��.t�4C�V}=�}Ҧ�QI�pZ7��fw�䙱�[��{�]�6�������o�����0�����mЙp��n҆���("���p�Т�t��8m#.ܴ-Z�꼪�b�y�ċMv@\�^z�QJ=aը�ߓGzM�%O�[��+F/lb��(ac����bzm�6�ߟ�0g���)����sc��^1+�
2�	]AlH���B��m-S�f�ٽ:�$�3q�>0��$�1#o���fB.B*>��Tl-h�}�`�d��D�}i��OL��\g��$2����L3���N�ѽG�ὠ*t�@ ~2J�*��J�m�11�9�]�{���6��s:�B�ք����ji���<�b^lr
�2j�/>A�UUy�iaV������_/�yk�aD��,��Y���!�#Q%̓�ŝ8�<�����C0���qx�C��0ɝ��'�y0��y+4D�p≝��/�;(<ؐw6y�]�����!h��Q������ꎫH`�ԯ��t�@O�����8�|�O�����A|�y�=9ɘ�8(�Po���ѱ�=��nd@��$V{?��]׺���)/u�X>���Drkf��¬Mo�r�G�V2c_E)K�8N�r`������XWZk���W�0�&��`��T�����l��.[A��l�� �6��Q"n�RR59�8XAf
\&g	|��Bє�C��M�W����_��K�yp,f�se�� ������%��{b����Q3?  ��JR���wV�Q���q}�tG:�]�,_P8�Y�Z���A��bP%�ZUk�JJ�PexIq�Z�s����]�Bx�~�fu�з�Rv|���~w���0�7Y%3���-����dΛz�~^�Y�yǼv��e�+t+��b)k� �Os�I���.:��Ud�/g��
ў��<G�b��섐hf�,c�S����Ã��9����f�⭓�;��Iۀ�^/.�����~l����}F�'��}���
D�r�@��:Bxm���O����c]���c��K�`�����K�s�X�)�V��z.Ϸݢ���!�	P^�W��Z��[�>r�,Z8�î�%MGF:��k�����qU(3�2��ZhE&��!���`!R���^_rFh�u ��!϶��E!(X=�|Neg\���M����5��R��T���E�ž�2�Dy��:�.6�qEc^���i�DF�`��mk�=c��q��i�HB� ��c]r��[�lc�@��^
�I�I/\3�e�ɱ�q�	��`�!��Y ��[M�ga��%�-��4A[y��l-���?�"O�漆�c.�-�
$Ќ���V-�>��:j~ �<����4ވ�rp"M�6iJ��rF��{c�13�+�K,ǂ��͠{��]����|8��3
`Xf:ηIΟ�6ʦ�_����j�
ކ��#�.r))J���h/��Ɯp�}$ ��=P��1�R勲["��fuc�rJ��	wvP)�N�]9?���YΫ�*��p��}�T*^ �z\�0���s�Ԃ��4��e7wdf��ȌeI���z�z���m��,\���!��6I�)����nn6�@k�~����/�����y+�'<�2��$��[�旻ZH((3���7��Ⱦ9� ��?����Զ��'Q�#�<�K��E�hU�p$dEe�
�<@e�w�@��b�aO���W�+_5��K��3x�+Ci�5>N�C����32Ʊ:v��-U��FZ��!����ppZ��;0��0�@FuqY�qZ+3V�7*���i����U���[F�]~�w.�VI�عNӘ0�L���3�����y��ʐg��vGlf�%�8�ͫᴄ���ὁ׊#reJ�\L���*`��m�yJRN��/����5��/w9%��]s[TS�(���J71�tI)���f�b��k����g��4�.�E�\�*����"���h\�ELQ��/���1�'��7��A�:�h
}M>��q*t�t�f
������@%;�A�rF=a.��Ҧ*6�	�X��c5%�0|��=K������}�������w���Ov�c߲s�q�^i
�lHz���9��s��fݼ�(��4	,0r�B)�Í\ǰxĽ�����3\��܍�9��U%+�9sQg���]���i;70C�>��k��ò�(b,T�A�M��{m�ܥM+#-��.���?�gOHF��o���}���3�ϓ8�ҧ�V�*�D�$������V�7�Yh}r�e�˿�(-(>�~>?UڍM˝a����Ux��q:�2�8�*�ڹ���4��4m��-�7��x�XȦ�v�p������謧yԀ��X�3�kn�Vސ%��-�Bs?��(4�d���,�oz���a��Ew`�(L���7�Iu�����J�w)��U@1���_C��\͒5E�g*+G��o+��*b%ӫ�'�����#`p�&���?¢��V&��vMp��bL�h���h�F
���-�Y�#G妬����-W�t�8�G���A�qZ@v�ώ=��O4���Q8�k��%&�J<�����V �8� W����Q�3���L�������yB:��{�s?G��&����'�g+ Xi`�vP��蔳�1�n�X��d�a�1@dRw���֖�9�������X��gmA�"�Aٟ�|o�Ȑ��(���u�����85XvKJ��O��q�vY�w�(j���",K:Z�']�I�+/foF������+��B�#��Gc��F�������R�����oi��T�{���NJ��D��Aʂ���[��qh�L��8�,�8'b�����e��t�_�g��k��e]C���q�[�*�&Ql�n��]�T������ȑ�5�S��j���3�	�(i��X�s9X}�~`��a袟���1�ܸS���)�q�}(n���]6���W1�7ԫoȥ��]�����q#T�&�	ϙ
,"&��A�u�<u��@o��(�D^�<V<��ѡ���m,�o��`S�in�(;��mXi`�d8���k2r��b熠�A�REf�<4�Y���9߻��Q��+G��kF��s/�-���m�[=��k	X�H�_�E8��\>[O�ͩ?��j�������0F���LHy�إ�겊�������=��*�]�3>��K�<p���s��H����ɜ���=��٧xam.{�H���q�kN3s�����0/���d�L ��k�zNjx�z��P��R�����d���ܶw�]�z�����b��F�6�n��/��H�v֫���RpZ��@�or�s�̆gD�2���1X�5O���o�i���F�*I�m�t���͚Z6����E�C�&wB�,����F������f$%ޗ��~����n�gLP�i 7_R�I��#��`��D�z��;X��h@��^0G�h�&a\�_��-���i\y�aD�xI�]�Jc,S��RZ׺�/�q�� �������LTJ�>��"̌��,ူ��)4�z�ݶ�:!*��H����"pJ\M7�#D�f�z���4q��|������+{����'+�׶�s�ޮ�Ҫ���6-H�@�b�hu���r���u!��n�QHț���3���BN��,�W����G{�>�:|�v�?�|z���x�+o>P��w��J��ղ��hX,��>�>^�D"�:���Y*	��U���Eo���!o<�s�����}�����}8Pw�wu5�aε޷�� ���-��9�!�U��d��k��ŋ*��@���mdH"X�_!W��2����/�T�ѿ����P�Χ��E��}��moB.�As��ܱэ�����IY��~�4u�&�CA%�҉]��I��v�P�������&�>k00�4)}y]�UH ����zW� D�P/�d��a+W�G	���3BX϶iQ;�	���N�h�W�t�5z�5�q�چ�V3.ŖUgn`і,�1b����9l��K�a�H"���U]�_.�*?Y�ԕnh���i�2�}�wr�`tZe�����p"��"U�R�M).&[�n�����	$�n0��ڟ��ZG5��0S�j_�@R��dr&D"�U��Y2s�����6���K�_^���%��rz�?�^�J |��T��:7���
@�ߪr=��{zyM�`�O���������ov�CXh�C����N���h�Ѷ'.۝:����������%ԨVg*@��YsC��K�Д�A�`I���5�F��1,PlM��ЖĬ�'@Jlݤ\���$���r>��#�0�����$:>M��'5��g *<�wv���y�݁���Gl��2|�Jh�������W/�I�\�Ź-�zΗ��S��:��G��j.銦%���?�.{�g�*��5��T��(6���8ryG�=�D�â0��ƞ0�.����U�p�:���*^Յ�dTia<��Ӗ�t'qdʑU$�lc:~;#�_��V�f��'D�l�ի��kn}��Zo_����co>������w$�գ�<ͅ�~pf68+r�<�PJ�ʍ���#!v�b,�����.J1,Fi����(A :"��7�Æ���	�܁KT~05���1����Q��R>���a��w^�������$��8����sqK� ��Ǌ��<�`o��8����|��8Ak�{�)6F�}5�?��6��{3�}�4�_0��V��_zs
U��sG�� �{+}as��	)�p�4��Y8�45)�w��uy��|��/@IF�=� |p�߷M�y
4��p���JN"�FO�U�M@���M�;�f� eC�?�<�d�j1�t��z�jmh��Ca��H�!�QK�X,:s^݄\0Ǟs�(����J��_CȲ�C��k# ���eF�z��\�I�{S�;O�NIχa�ť��JA��o�Ԗp�i���+Դ�.Y]�ƑqKl]�"�6R�^������R�x�f�w�$�?wib�dg���/g&m��EK=j����37�x�)�iT��-�H�u��5N8�іs�~�TJ�;�B�����'���+�
�hN�TB%�#���K��JqZ�җ>t����%~�TV�I �z�j-D_����at��/��S��f%�	��������cA�.�	z8���u�'+�����r��ޜx��|gu\Ll#�&F^�C�g��c�u"�|�>@�,!̅�f���/�e ���ӏ��������Lg�]P��c���?]~�����몧E.֑i�f��+�v���XW��ac���AX>"��1�?c�"�X~�B���5�zlf>��)�ZF���}m�_�<��?c9/��_(��6�x�0�&m󋖜R�ݸ��"Řǥ��Àh���qE}��d�h���ß�򊣘 �B�//�e�����c�)��GA2Pi�$�}���� ��Ã�M^���79��Ϭ����1	��7ܤH�O��w�ЇB�����ۍ^V�4g���òR��?�iѐ�#\��yt����\d`h��Ox��DW�!�}΅���#h�Y�g���ZjZC~RlW��(x�#d��~?��1\�Y���|���Q��m"�c
�2Me�6���~��+	�����Gg����1�UkԼ@������	��@v=<��*+��'mgg�WH�F�ȩ��)4׼xI͌�¿s"�c�(q&t�7��E�q�>�G�_,�e˵Lo9!�=�\0��خYmyakӌ]x_�V� AC�M���Q���ɥ�摇���;���V�m�c��a��O��f���!>�,4K�$�Z�����i��I>����
VG����v����Q�R<]�N��0��O�?������1pd������1��8Ϲ�A������K����
:�r���P����G�g+��j+Į�d��ԧV�ŻqH�T�	 T2�O�F�Y�]��bF�l8��o��7lkn�H���9��'ћ
����y����Q:�6�1���"�
��>��w��/[�e��lHJ큔���a�9VDZL�p���4kq ��􌬐T�w�Uas�S("�S��M))�8�v�G���B��)W�T.���$eg�vЀ-����Ǯlh���[�U`��])���/%x�M�zb��N���}��Vk�e�<��_C�C��̰��� ��QiM��^�����xP��L&6_m��Ǘ�;x>+��;�m�ª�=#��4Ru|�Q��QR����b5�����Mn�u]�ˤW\ڢ���˥#��E����^��5Kڔ�Ȁ�U �#��z��ZzS��.���r�R�p}I=��D�lC�/�㷱Ҧ�,YkW;�u�J]�k�_j!�3}�R@Ꝇ#0��`�Usbm.@
r�΃��*��#�� ��WT��3�d�ȥ�Ɓ,�H�hnz7E���x%t�?�rRd�O���:'O��pnB���m�Jv;����T2W)���h	?��6�2[8<��~6n*��>��Fvƛw�����$i
�RU|~�I��'؃f70�~�7��:�F�ۦ^�j?r��p �!�%�p���'^�Wy�u>���7h�g��^q�����.�dx�.,u	w����0����7����#�ͻ�ū�`�Wn���_�4��<#P�S�]y�8����M?�r��"�QU�^��E��d:�x�sw75��;0.��:�`*Q����	
D`i� k�\���n��Mg������LM ��1�S!Үѱ�>䩫m�U�Y��D�:!��{�;���_O[r���WIb��#hX���;t����kV����A�s���]c\�r�����t����m�I�e��t���D�ɶ�u������q&��d�m�igU�
"�N���!䃅�ѿ��0t�F���_7y�6����nb�G�K�lήk\����FX��l�M-~��^�kw��T�$�ȵ�ɚ��?�]̅>c�����h���5+�j�#	]6לM��Y^�|Դ~���U�P��ӻ��vd<�~Z��1{'���Hم����5�ϾC��`^���:��%�/^� ��C�N�MLB�;�p��zV���������3��N���@�*�V%�Gم��.�0w ܜ�b�iL1��Gtoȟ�֫�g������'ib�9褾q=fJ�0+�HaZ�8b�x���p��z�@|�]|�d6�[?̞ъjW(ŶN�M/��AKo���m�n@�i1^.'%x�Ed/��L'��}�P�OOj
�"O?r_�&�(�~�B�c 3 �^L�Po�*}+�%��ږ9ݡA� ��@���>|{�/�������ɒ%=eA*Q~�-�,�״W���"���|��I˨���3��,0����5_�-	C��U��q~�`�V�&
��k�?�a6�i��r��
��,5#^�f�쪶�FN�+ͽ+1�]�s2�m��{
��#��ܓf�DTV�]8�����/p��ď�����Ug`/1��T�v�"r1�{��J0i�Nsr�| 	��f�[m�d����ꑀ}���Y��=F��V0Z�[����$�_;VYn$�z])��Өͫ�F�)fO��~��֎�[eU�
�����H]=Q��2�>���83����b���j#��+�$(X{����I~��ý�-]�#�mv��Ya�(�Cѣo����k�zl��tmgR|[�3LWv�	m'2��Rj!m=��VſJx�|Q��:p ]��~d���������&�>��K_����h�N�;�˧�P��1��G��,ñ:���z�wsD��QE�?4+���ol���s�r�V��=)i�-GǿE� �y��ذUxK�^�CV������86�A���a�����x����[爞�b�ߟ����zB&��Q��K��crZui�q��|�:;\lI�J��_0�M��N�<) ���UҠ�̶��OC��Jr̧7�g�v
9!���LR/'��M.VwFh��Ǔy��F�Q�M�v����l��@�OL�b��L)��^�5A��GlVO*SzzƊYK;cmv�i	��	I�8� �9�SIp�mLVl$�t�+��Zc��EhY>@��2E�0c{��=qJ��}E��'z�|���v��#���ь�@�:��(���$Вsl�I,�|}ۀw�ؙ�2�GwՁ���y%Ӌ<��=9(�oP�tё>]�d#]an �T�� �В��|��d�w�.�o�b�;��?i३e+n��2�������X7�J��F#�_l-�%���E�')�E��j�{�Z���� ��&r�P^z�)���b^�EQ߁��������a����O��mv�\�_zLC�~�, �N֬��m�U�J�	���QO��Sg/��(S�(k��"�������ϧA/O$t6v�&�j�H>�qO����_�U�BP@5�FQ_�,�^&��@����Q�����-Y&@�.����Bw�:>�'�u
0��Op������Pk3���jN�%t	c�T�����fN�{ͣ��;�~O��Q����X�oE �_��ȣ+OS��� �����g�N$2���|��D�!u��~HF��z��S�U�
��a
E5�)^����{ĝ$�J� p���G�aT��*^��و���	cÛ�KE�����a]��'PJ���@��/nj�O�Oeٯ���f�i��I�[�z6���\k���M�[�{!��!�%�)�?cɻ�]����R�cEF@���e��v<BUnkL�E��� n`�Qk|;j�=݅���CjU�
0|�p���9��[�����"2�������T�9eCV��r����j��<1M���E�����*�$W.X�T7�&��Ĭ%����([�:�n����1L^�PV�dW�`,����]��9,i�<y��G���c�+�k�J`����_bN�!ML+��u1�W��
�D˔�^TMc}ؓ ���_��'�@~��s��"���rK�*NG�2��7l`	���\@}��
���5�5����Ԏkk>�f6�^����
b�1v|�W;��2����ܾ�����${�֕��;�IZ����HM�+������N��:���3ָ��䯰ux'D�{9��ho�$F��T* 2���uH?oH�#���D���h�C�倪4��������zR���������Q��3��cŃ�u�>a��U?����Ce�q�.�<��q4p9�����jMl���h�~�{�*LI�\"��ѽ�V��Ҟ��(v�|���T>���Y��	�V����y�2�a��}j�35e2s[���G�D !�$���kF|k�ⓘx��GN#�К�,��E;��7�ˌ����P�8~C��Xy��57
�G+4Z�QA@{��x�9�-�q���?E�Ŝ��5רb˰�g|����'��뚺z����ͮ�Ӻ�>�����(�2�LZS����L�/�{��Sy7�E��ҫpVV�U��1:�4D�D