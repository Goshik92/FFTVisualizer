��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�K����]� �h%o츅��Jʤ�|�w1 ��"������]"⭛���]Ul'�q�d���C�^jds��'�vк��gL�ZU}�#�}���T�TZ@`��c4U^80��)I&�r�U�T�~)��7;��	m�`�~nӸz�E�����2�J�q�D�ԛ��\�]�奆޸�a�X��ޛ�����{L~�m�ޮ#Iu}�:�WVA;��D��&��(�嫋�m��rӔ��ˆ"�L��-'��1���6�6�L���
��9�{���y�&�9�gi���!�G����Gqz+d�6r�x��ǩDi�8U")�r�xF�3I;��R-TJ��ߥ���"��׮ s�ȿ���B�C�"�9�2�z��3u��a~0ݟ>$9�w߬�n��c�
�n(�4����P�=��Cn�"PUŷ0�19%��'o���a����|�<eq��ngY���"��R=J��M�^.	V�O��Id="xC��m��b����j�6*�Fᦝ@6~�з���2!�n�_�B�/Pf��p���� {ЛS�U��?���y�������'��p2�vC��݃h�HR�J�P�lj��'IL��"%�)D%�iT�B�k��G���+��3��j���>����*��ĵX�{����cizxE*ڣFI�Ǵ�׷���/���`;��j�$�L��\����^.x��y�I�8Λ�~���D`���M�����;���.��6�ʈh�޸���X<����1�����X����(�V��Wc�Z�7�\D1Z�ʵ�Y�]�kA�{���Qn�s I:������u�X&}53w=������x�u��Y�P֪��Ox�U]�{��e]v�'���}*�ŕY%`ėđ
t���z�`Y8����MS�uZ`9;�Vi�}���t��ga��&��&�t��j�9
�0^A�ٴ��2+���4��rv����㓎�yX�� t=R!�㲏��F�1�r�dL�{�}����,���C�4lCdି�ݸ�5SEV����"@ A�2=Y�!��5�[o(о�cH�kz&��+_�ɂ�Xbl���T�ynػ��"�^ESH�w\Le�<��	#���;`%����́Uir��ηF�|q�?����bl6Q�k�Ko�.��@Ji��5��5����g�g��٨H�f��xڿ:$ @F3t��������ӷy�q@l;c_i�/��3��ӡ��3������x"W��4�mvp̙�[�e.e���ט4��03j	C(�{�d������������r����k�0�<���u2���7ά�{?�:H~x8|J$�W�¥��˵禲�*���b�#鎄�5�2��s�UBe�����P�_S���[6_R�������L���+��햅�g����|�xn�S�i��m��%|DA�^
p-Q�3,��\&���L�3Q)l�?�9�@����:��u��6��9śCɴ�/4�f4�T�3�d�,L~ R���8��÷�]�2��OS^�|#w�C1l�Ԁ(Y�c;�l�h�{�m7�5�P��}��Ǆik�}i&�=�������@홦�����	�"Y��m�8C����gU�Z�k�g"+�x���X������N�����G�b��՟��6p1�]�p��K��f]T����2R�ǆ�MS�Z�ʎȌ82��[�`��Ϧ�B���<w��"�>ဠ��T�N)߿�����,��)��B�f" ��P�,sa?fK)�6��A�7i6�����R�3e���"y�c�}���{��վ�oj�㇑a�̗�hd��-��^����K�� �Ƕ��e/Uu���:��|4�Az�V,��q��˟��r��A��,�B�K]u�(��,���H��N�Q���O�ROr@�[JTc�F�j�%(s�ɔ7�����wet~��}��`O|GY��Y�^w���)��A`>h����Z�~�91X���W\${p�j�z�X��� ���3Ls�|N<|Չ�4�.M�c��Q���0mp=��Z��_X�*�(��8F�=���^�i��U��Z"	
P�bZ����A0��A؋�~�i�eB��Kԛk~��+�K�A1�u��2k���@3�+j�R�]�K^l�֗5�ªs����kw>d�wi�E}X�S}[}G�z ��p��u�2�ը��1���0GaC:7�-�L�Vb`������V��&���l)��� ���J>�]s	S`E�;y:���W'�@|�qXo�k��
"^�Q���ɒ���Ħ N\D�*�/3@�%I��.u�҈vs����\�[P�x!|��.6 �]�[U�#��آ���Mxe$���C�'n�w)�*�;Np�u�6(rjz�/�}]`F"��ݑrSY ���ۥ��.���6Db�a�NSU�VV�j����j���6�qC�Ĺ��uFڣ"�쵺��@���)�\��#�����dx� �ů�&�6 �p��a�_��f(��+�.�v���w���:.՟&��3 s|���6�����YR�t���6��_� ���?n��'�L��e���m�;`�B�5����M�R_H�����w���f�ڻ׳���k*�~���$���-��l.�����4n�Q��	�>�2w36��C���;N�B�L�Y�m`
����Ŭz�-u93�6�� �VSp��`m�K�z��+*�b4�̠ߡ�T[��vZGb3H�h��#B}Mi}�Vp�e�-��[��mn�W�
�(�oJ�g��(M�f�Kv��P�so��3�H�Ϩ"ZfR����3�d��cd��a+�V�M a����9�>�n�@f0x�*���M�ݐ���:�azJ�с���yI���{+rzy�byZ�ΗR�e��*?����ٓ�m���i�j�o8jf}'�k�����N��:����6�`�&�s���u�]��{
'2�_�t�e�8�J���v� Wz^*��2��!��z���D��E��=�@�#�7ڙF��
k���t�9�S��Y�z�f�C�3l�#�a��x���iz�U�j��~�6a%�77�t�dM.�������	n�?R l[Y���N �15_��\�^���x�ʫ�ع��|�^E�F>�ܘy������߹w"��̢5o��9�S1v��i�\n���N���8q��^�73<��%�-��1q��s���gkm�?J�YZ�
q�y����<��aȥ��ˈ�WG�E\�+���b�-M��x*l���rՃQ6?�J�H ���oDs3< b��S�����O�v�b��$�3%7�n���nDr�R�~����O�Jy0�]���(m"��/5�1���F� P���Ւ1.�f��1l�p%)V�HX��5z����W*nxG�{��?��i�ֻ� uyG����ix�$��������Ŀ_Tѱ��WeYl= ��Ȁ�����)�ZV�������{C}LM}<
�J��tw��?�14�&E�n��-Q�6��ĝ:��E9���G������`4es�pv9.�)G��ҍ]I�	0�8�K�G�m�@?�H8lwC!	�hH�F;��%-�Tx,���S��W[�i4�-F��w�W9�f��pv^������E�5����1?Ł<���|�7ZF��-��?c~�������:ԇD�y;�)z"��IPd�wx0�q�����`��� ��Y
%ʌ�ȟ�K�$�U`����b(ƦlK�6��&�+D��$/:����Vz�X��sd���X8�����l����JmRи��(�Ǟü�*��O-�5��N�;�L?��,,�II�Q��>=�q�)kvspn�����Pֆ���� �g�wu����.,�:�h�DKI\�B��a�;�H>�
i��Xv�#�-iD���'צ��Uȥ
5�4O�iO�?����\���C&K�t�p!Wa�3͔��|���P�eT&g�(���tz��c3��~˧t�t֒��b�Ij���mc�h<�q�?��j_x�!+�S)�qm�SLb�]��\[�W�:XƇL����J�YO��Gx�my�4>�w+Rw?����U�S�N�ԏ���ۢ��&�e���~|$MdƱ��rç�!�}Ah-!�xw�`��D ����>&�w��`�����TW�r�8�UFO���H@(X�����s�_�}�Z�;PN��X�	)�܄�/D@�@K�Dvj�`J�Iu�h9��At�Lm�ŷQ	/��W��p�02H�G��u/��vf�08K���A��D3'R ć(�KpnL�3����E�v߳������=�_v���z��)C���ȥ6����Ԏ9'�E�G��>�e�ܗ����Ǎ��-��i��5q[$�0kv�l�5T!Ŵ�ً~]���'�⪐yc�nwa_��7u�����= |݊�#�FʭPk.7;:)�R������\M�A�U�� ,i��]2��RC."3^
�D7� ̶�P��t�Ɗ0Ks4�|��N�Ù5���<��_��ՂdIE%n�FC�L���˗�[?qp
�N������lΆ,R�b�ϣ�z�Vh���<R>w�ZZ;@���	�Ҟ�&�xG�u�%�6pH�#�3mle�Fu���	�%��n� �NX�G�Y3d�EZ~"ݼ��n�1�,�q9+���7K�U��n�Z�q�\�{[��S9�B�E����S��$/�]щ�=�t�v#:p�Py�c��h�z��Rze�prx�~f$'�\��$���gGp�P��>�'C�(7�}B�"ԽhC�9_�QZ���/�d�PK���l'u������p��rx��,�Z��)��ĝ>�Ă���`L�b?�*fU��Ti � ze�#W3�a����0(f���;U7�\�Z�#�� ڟ���jg�@iu���f���O��47��>�-R6����͉�� �]r�g=���N��'�1�Ǿ��^�6*s����̧�i�c�,��oqsՂ̋����l��8���0��yy�>�U���L��`�U��\��s�w���a"�2�ց��Pb����9�U����g�[\s��͠V�LP�?vJ!)jsZeB�Rv-�������eI�tOg�N9Wg�Z��$��r��W�OG��vl�: eE�k��Ru�n�S�*�P�wr> @n�"���[��@�~_�`;5D��r�P���U�P�[�Or;��s�^�W��zc�Il�n�����I��Uͅ'�ȋ��Pӛt�{~�Jk����f�n�œe����8n�Z�E�)/Y#m��$8d�{���a7 ��7�M��|{	�Ӎ���;A(�Ty`Y�B�Sd�~!޷�=��w��r�����o�����1���:q��fG�}�.�a����|�F��j�C��]���Eu�U@z텈*�/��I�K��7a���l|�&��&�ބ�$%�T�<k��l��i�/�N1����������+8O�^��|���]���4;w9���K�)Ao�W��ϖݵK��F�����w��U"���Y�c��\��^^ɫ����݋�W�4q_�xХ��<���@ =*(�Ҿ��j���W��u�����<�,�#��e�q,�Ar0���fq��<l"���&�CˮB����;� GNG�H�(Dq?W����JxX׌e]��P��ޙ8���Y�-jO��ӻ�tE~�k�Ht\_��L.��I\���H���I��>B�buq��8���j��U3@q�u�����s=�شR�Ib�;Z�BXy�~
(g����uf��OD��fj4xJd�l��ŌٔTL��s[���x�#e�QXl�'7��Ժ2�1bS��-�o����������u�]oXګ��ewh!�m�N�� ����RĂ�h`�8��r�V��x�Xl�M��q��䟯�s�h��ʷ*�-��d'�?k���\�]w��~$�қ�e�����C'��$�z���tc
-duѥO7�m�C�������Y�0hփ�ׂfv 4�gumz����NA1�s�gOn�MS�ͨ��n>;կ�j�����3� Ko���M$	��O� x��VC����h����=�X�VO��=�C������P$�����~C)M�on, ��&����H���ڼ�9��¯���á7�q�t#��jb��m{���#v��VO� t���e�̱2T�ː�*��ȑ�g��ci���ū�&�=�EPSu�=�_�Ɍ��9G��E�N�D��7O�[⚱���k9m~çl�a�MĔ��S��;��O���#��i�QΙ% �X�"�%�3Y4��R'�����Ҟ��t!`!�~Fg>=����ROCjkn!�e�k}Ⳳ�06��I�B&Y����$��0vm��S��[Ek���NX�g
��%��Z�'��jR����s�q���y�#RH&5����r����h�UUɽ<�Lx��պm���a��(��,S���c�G�V���%��:ʢG����O���(����:�$�4`�~�
q��0i�%�N�aƠi�Q���;T�u�������Ԓ�òI����5k�,�����&B	f0%���ϐ��YYx�s���f���Q<���]�c
���Y5�I�)�����Mh�S��e�>
P�G�� ��zH���"@�R �+��_�� �h�x�qz���Y}[C7{�
�@O�z�.1Uh��S:>�-o:�TY*��;�Lߤ(�,�&7{�1.���]�e��}*ÀN��dL�+Y��SdP�h�k^~��6�h6sj����W%���ځ|g�'Q����ҳ;�{�R������P��H�f/���Y�Y���Hz���"?[:w���;I��X61�5=2��;��,	��]�P�c�
�B�V����ӑp��ȄA9B-�r�ݪe56ڮCB�