��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|p�n�U�d��Lx����D�~�dE��!oC0���ñ��t��!����ε���}�V���2��˘�8_� �-��Q�r�eH�<1v��b�qj"|	s�z�9�q5�|��,��x��"�Q�z��Ml� �(�EVU���+"ڽ���,�=+�������j��{zh�К�{1&ě��d�nF�� w�ng���E0�5� �O�>I~��o9�!u��&?۸׾)i���-��/� P����χ`ya~��(.�/��a7_Nn��΅lRT\;t���?$)�����_�5U�B־�zh�a���$���bL�K��<���*��.�6�
�x�BG��h���C.������Y��xg�"/�v~6;���v�l�c�S.]G햵�Q�}ו�
�e�2�r� �P��]�Hn&'����=�\PttZd�	y���bLO��"�;�!�L�@x������� 3�]ʧ��g�4���f��фE�ϵ�۹����.��#7��!ƩZ���W-e?4Y�T��dĄ������PN��w7�G������R �H��V�+a�^o0��&`���ah��~C[$֞�x��h�7�r����;�r������9�q���۽o8��6��K�L������a���ބ�ղ�5/�A��FeU]�,~1^��](6 /�I�Ef��
B��:y���$I�&5�7+�Z�n�,�\�װ&��P��0��(�2X�����?��9���ofSa� }+=N�ڼ,w%ֺ�	�k.�h��'�m��� �A�9���Y��S���:����(�S���gM�̓��\oj�����m�HԼ��0'@f��,����.Ǹ�J��B�<o�;UvcL�3�zj����D��>y#���V���y�����E׵�fP���OS�q�0�!�����[q;4���L@���ג2l����L��-���\dp����I~�V�a�`��P���|�Y	�M43+�w{D%G��3_5g7�I˭r�.���EtXg"x%<��a+�Wy"^�-�~c�1ꬹ����᙮�Jş�Gʌ�#8��^E�-�t�����R�N���TA�)�Є�R���B��	�e�Y�6jA����ɍ����1��E�D�v(��77�N�ǳ���AD�7���u�L���˰z@f *"��Q��mL˭n%�䭨(����^%�ӘTg��Ic�T�r�b�3��c��5��8�}�ʍ@a*\$;�6TSa����ӄ8��3��rZ?�߬C�� 8ӄ���j�J��C�IH�.����z �!q�X�;�%�q;�טR�}�֓�]}`��y��7��-n]R���`�#�b�y�|�.�!5��HR���-�@��g�i�j�6"��*�KN��������)�-!�׿
��5��)ڌt�%H��*;��E��r�U�A�Hd��I�yj�.]�?9���Y��Ğ�.UOcJ܂�Q2B����7��j��Ҥ��1��z~�o�E�R����z�{�,,ŏ�4��<���v�����On���h0g&=_��x��kɛ�vM7Hi�;�{&M8�������-�N�i0�ji�XZ��s�S�#�5�@<�d�CE�a��:i+Xm���i_0�-]p�M�K�:�h9�c�0��9�Xd���d�����U���5
$���;ٯe�-bwF��pN� �A�㮢1{��#�7
�����|��b	S�4���(ڕ0F���(fTi�4TcB��;b������o_.o�7�[��ys����R߂} �-�d<_��@���ǘ��Co4����)[�i9��Q���9_w}"��?Q�����_��Ed���%���WےQE�N�!���,1+��(�9]�C'�F�%����2�tPH:��4���u-'��j��"��̄�D�(����҇:�6�^4��% E��F^e�2�!u���%fg�g*/� ?���0���P�ˇ� ޟx�8Pd�5?C�t�͛;B��n����c�qX�_aW� H�~����>\���8S�K��g�|�T�JӃ3+
�&K���/�x��O�su�U Xku< oMJ��%R����l! ml�9nܺ�ѦL��
ZF6Zo;Q�ޏiҖp�FRn�����_��s���b@��9�G<`���+�$V�?�uN-�T������wPU;���H��S���2�3�Q�_v�q���y�p���@}-+�Nw禥߶mg
�Oʉ'gn>s!�QzSw[��cmt0J����u	�����s�1�2����H��e��*� BC�[�Qxp��R�zF�Fbn����_�	��	�JK�`sEWZG��k�`�P��p�R�(�/M�������[	4�E�X��j̽ǐ�v�7pF͋7S�U���4�y?�4X�P�ڏ_�zp�$2���)�'8
�m�'�y�W�-��0 �Kg'��_OF
������Ͱ�!0�Ў���{�$�DsW�e������
˯����/e!e�1��l7�_j�6
��W2h�&,<���E�:��w*���k�3���u<�4n�����P{��aV�](A�u_ﷷA��<�A@�_�����<�Z��Qm
���}�P�����C�|��g�-�q��M�!������;�4���!_�'��#��3&�$-��(�,�lńmN}^�R_�G���.I��y=��|���|-O0A���q����a��d���֫��='v�?��u+b!]Q���F��.dk˫����*�,~�K��+%��0����͞�U"�M�u�Aa�(�Ä�(�Tṿ�ƴ~��SI�����B�M$��E�0�>=�RX�F�}9Ul���W(FX�O1���+M�ӝT�E���\���e����B���..dA*-{+EJ
8� �p%UU�P�^Õp>C���J����nLr�@��S�7T9���N�}Qqٖ�h������hӡ������eH�fmٜ�F����ғI%m� 1�&!c���U���t#�b}
➙�c+2C��Ա�1������
�u3�9�kPK�鱮y��H�@�Ae�r��X�d [�@#,]ٳ�����#� �[='SR�k���Ļ��WG�g0W���F��>�
��Zm}� S����&�n�o�;���.�s����l4�K	�ٓ�c��$�ّH�2^�4+��-cXݷau�R�U�h?6�t�N�ç�m��Җ�tt�����>��Z����㜃9I���;"ᥗ\�FK�dd��h��¾���1���F���	Nֻ�5B��0���劇q����9BO�7�q)y��D����\�4��>ӗ����gD�����;%�m"�э\OW����ৃi��v�o��*�Ъ��ݨ>kN�pY@�<��]1C� ���-u�V����B�lG�
�S�Q�:
~����6�>����5�+ɓ�wEA�;�Ժ8@ţ-����l#6��NS�(�6�ճ���ӜPu��g9r�z��MY��hdb�������
�r�:3i��`��I��m�_��b���>��ӛ�(q*zy�^�@c�#����|]�JK��|5��d-�W���՞`��zW6w�S�ܽ]��O�Y)�V_�?���زi����6���<W�?�4v�wG��l�����	H�H*Rb)�c�$�N]o�!8*M���c(��@h��3H�#.�ceЅ	�rc��林�I�v�j����0��lA��;/��	K��i��5K��Ĝ�J���@S���f��M5�
�~N�5̪�˽.X41V�)IR����}�=���c�|���َ]��J���4?}A=��j�4�t�~��ڧ$fG�)縅�5��Ř7i�ޚ����Ou1�1�W�]��0�C���g�S(�
����I��[�VWEVCDD�AQ��r~�@�V�\6��ܖ���gr^'���{�ś� Ml�r����� �Q!�u�kob�?��=(A �#��'ݍ�Vo��TTNӱ4	`%����U�9�wH�v:�&h��۽ӢI9���C��9�'7�ҿ�e��Jƞ�u��sSØ��\`�>��^�Wƹ6P\����A�V��;4��h�>Þ�������F`�u�8e�,"������٠6S��f1��:I3=;=�!`�{�!h�?7��l�^��!Ԧ�K*�G�~5���.��촬p�ݐ���!"�3x^Ȍ�3�g/)�7;���|�����}���w�7�`��_���S�[X'��R��͈�~�v+��THh����H~�v7����t8�4���G�����}� ��\���P�)���)���7���j{%n��n;kA���v�\8E֦=����q#\˫6��Q��<���0���ه�(����B�`�x�~7oՌ�����
p7�(�etw��Sy�`����;�H[��ܸ���V�Gh��/n�EhHVZ�A��n�@��E���I�GG�� ��Z���"pΕ�o(�J�ۉ��aS��Jf��D^ʿ��#%$?]�4�&�t�K1~�e�M2��dz��ϖ��@K�n���}S�>�	lC��XW,�DzhGl�8B�[��i\5�pU߇<�=��eH~�����=k&ӃNc�ð��2�} �k�Ǩ��
�?�=���La��Oi��	ľ�] ����"���(�>�Im�?}]]�J�r���Ò�EI:�ہQ�ˈ�S��\���~S��fp���X��7Zwվ�."�&�D�_/�n[[$�V��e�6x�K����p�#��9�P@,��=�D6�rn%�S��*iR���s�g���J�|\!�
��,�5�>��ۡ��n�i��ȺO7�����ɽ�A$����*D�ZZ@�ǒ�NG �&�ÿ�0C�П���3-j-C�_����j����U;��3m�:k�	sɂ<�����I�!��i	�}��e6G��[�H��N "&ҡ�����yCly�x1��Sg��-�9�ty��71�Ε}�������b��X�0;qm��.���	�ml����G���J���><$��'3N�9�jK�^k���f�O�5�4~�l�ka{�CD{Ɉ�ZS��AP�	���>����{d���W��o&��Z+C&�
��}��}�W,��]8͒��Ke|�����m̤�qsW4C�sx�w#̧��k�Ӓ�\i����	X[����C��-������=�f��Ź=�[����T䫯�U��Dɉ��?�`�tRְ�s���,E����}Q��h�oiUƗ�f4�]��>�\�۬dt4�[�����9�N�6��6�ńtU&H����tt�K�2i��.Y�x�7���B��Y�U�m,�k2�R��cO��� �0�0Gm/��äQPo%E2�y��d�Vnz���U��u�o�8y�SM��1L��U�q?i�'f�<�<tu����3�tӂ�)���� ]0�S[�ĉ���\vPq�Q��i���ܳ�M��6���ׯViEL�ϢSώ��^H�{�x���,���ɭyG���/�%�\�������I&��g��9'���/�]8��T�7������-q�H��܏�%<��qs2�����)b9/Sƀ�Y����J)/z�Z�ު�xL�Z�<��Eh�R�;5�Օ��2�<͋�ŗ�&�A�2�E��C�	T��㘈�Ś��d�t| K�@�y�D=␎x;�f;T�EA�p9Gk�ݕ �\�/�&.����=�EڝA��l����� y���rR� ��#	B-p��^�j�Km�o�C!���|Y��'�{�V�O���*�>�O��v�3:�|�?�xXzG����.��{TYn�JwB���U���-\dr��W8����VO����9 ��L|��JE�y8�7�5#}\�83�K���A��I��ړ��C���5�-��d�6�������rE�)~����p����/����jP�Hz%[�v��k�O�T|g	�Gj!����`�o��@Zf��-.��A}�?4�,��V��z���4e�J�?�{|O������K� �5��/�w�D�%�����9n@�����%*��%��.�.��m�p�cX����z����݃eO(Y=�h�ʋ� ��_o~2R��r��1�vRº�Mm�3LJ�|�(w� ���j�vi��-�i���0��'G~kEDB� �޻�%.R��8>i]5�m��ܮ�x�r(P�W���&i�^��xU��	���B���v�XB�Y钖_-0��it��76�D��[H�M���TV��tf�4���CdJf�����Sdΰ��ϥ�X��Y$��&E+� o�����+R�,�i"�I�xc�n�chHS���#��i�4CT>���e��v<wr��=�����&?z�����9�; �Ơ.�n��a9�gȮ��RVc�[j��2�}	�4̡�!˒�B1y� �KZ�(�=���i-�5�3gi����Kv��:�w9A�1*?J��ȅ
�lȫö�CS�����&�*��H�*Ԥ�#�	���AB�<��a�펅F$�둻�j�t�l��|� 8���,��;�iκ�l�O���<� ���@��=Ž��F:�D.>�u�ԝ����|�6Uu�>���+�2��.���d:U��rsw��0�,96�����B�°�*N˖wv�#aGA����`ԯ�A�������(kт�6��Z�?|+��G�Qs�i���`�cZPBG��<T'7�k�Ti���4'�㾹�_�$�B �Z���4�ΗO�]����2Cv���S>f/�A��N~h <�?X�Lㄤԍ2F��1��ۛG� O���Q�C��H2�{mJ}D�0�Z�K����Zch��c��D��D�ij�\��̯0 �W,�� W}(�`�.�T����id�Ŭ�E�-�pt�$��\%ڎ��Hf�x'�ѽ�͏��/5	�6�J�nz�bJK�:��������BO���Nn��������)�n�����Wڨ���(,=�k�j8l���,!�:!�=�2�]�?P�myaa��;�jߝ�t|G�o���6j�dv�X��?e�6x��
���O\t�c�`Hxg���BSx���A.�0��1\�]A���ܲ�Fо���
fD(N�-�1��|z^f"�Gu�__�S�`��y���/5��끋�����g$�NM�en�R�}���߷J�s��g��]�[��f��uN|zU.��J���c�Gu!����Y�Tf��	7�HΨ(0�M"
{W�����#�2D")�I���MR��9�~��o���lq����#�l��{�����U�_��E�j7l�A�C0�$�Y�J�Z�}�ѻ�i�����#�WҪ�o�����f+})�6ɩq�h>����G22��#���֏�l��`u���%Q�M),؟�
`SA�����q����|~&%�&9a������ u�˨6�m�A�Pg�n@�DPT\���΢B�M���ͭź
z���.h׳��!g��������nz�y��(�7[��͢���k��݅1B�{��N��Y\k�.��L�Ⱦ3X��A��5�tr�ۙ3W4Ɠ��P��H�2���7&����p�� �ձQ|��*mk����q`�uS���<�W(��7�?H~@��cI���Ǆ7y��ܽvL��4���)O��dY��P�{���4P�͉����?�����F�=�g���Z-S�����`.����e?��糀�#Etn���8o�:[���]�s>���������B�J����3��%���	��������ⅎ�
�eq�B�R��:*�fuQ����|Q��ē\T(Wbo�;�Z�LS��06�M���b4ά�jѫ��R�T�*��CD��W3��:%�	<=.��	��b�	�����N�4L��b�F��Z�7#��q�<'�a�(�F�h|%����sgTb��ە��"��cP8�Q	�/F|�� ����h��8����;����U�'�'u�	|�����6r��&��>Tq�,�KH���2�U��Բ�z�qPg��g��q�zh<.�G�Q���1���㤋@��]�E�50.�i�j>��c�~���ݎ}� �8�>
��_��A�����쾖-�Uֆ<����F���Hx�R��H�#Y��c��;�p�1��5k���Grl�eD��9a�������oˤ��l�-P�^���1��­>��5d��.��M�JrԬ+'�Fli%���u���C⦲|?��s1:�����B<����H�F;��� .��c-�O~C�?*y�A�$�o}�҂�.Ga�z�Qr��*�̠.͔���� �XM�h[������Z&��������T��
wU4�-B���J�@u2���� l�P���3E0TS�n�c�m�B�:76�JnB]}�o�
�LZ�N��]��K�AP1sh$18��IcX!'~\st�=͋zA6��z�1��ޜ�[�G�mP��7�~���UX	���S�'΋�+���Ӯ�Y>��7LEj��4�D����~<Ҽ��Ib�W�9ɸ���/ª)��t|d�vtq+*�y�$��Yw�Y�Д=�)l�J�.<O���}�Q'�c+��<s}Ҿ�B�<wQ���0/(}���W�[���SP�gя$��p���	���o�b��?K������+֥;k��\��<�%Y�2�p}�\���hfK� ?ש�Y1(�?z>m�CJ?�{嘎��x�x�sa'3@���R���� �.������a��{��!��{̧kL��f��}���}����ۂ`��DW�K� �gf?�2�T�ZQ��DQ9t�d�P�0�7TBm���ϓ.�Sy�/QW@m����ӟ}�I:wFﰄj�kޔP����jG~���X3 �dR�VL/��I�a�u����_/���gȟ�d�o��RqP�a�����	ԫ�/5ah2UK��T�/�b��b�?�ki���� ��X�xP������(z���@�Ib�a��p�櫌�3w�X��Q�����"G2�ᔍP�bZ�MhǱ�n+�G�ZWP�>��i_��:CwI�ÿ��Cy���,�h^=h�%x=�8�Q�BY!�mCJ�A��W�j˥+�6t갗��d�lj6C���w04c�����g0VZqI��Z̭ק�v�d6���t�9n�p�΄�o�����gD��	��s�iem�����!�vVx��^pW��x�@Z��Po���[p�tG�ߐAd���o��f3��Љ$�2�u�
N�G��c�C��!���.�W\z��6���	�{���t&���e̮�h���o�����vuN���� U�5�[3G`2����vYhS~a8�s�6�&mpY#��ո�j��$�4Q�"��]]�_��do�̤���H/�z���n$�����iN18I|Z4��h#�}�%f�s��"�o��T�vL���5�?kVn`�"�4i#鋱&(�(ʧ[v]�Ʈ�{{����jО?��
�zz�ϕ��z��`D��\UX8�c�&�����-�[[5����QT)W}�O~�M h�E�n=;X��"���<���p��.�I�~f����uJ��J�)�ـ'�Ĩg{`Kj� `xЁZ�,�uu$hΒ~�/��I�?��)�^��$
jP��:��}��]P gg����E<n��A$L0+4+�w�?�����q^��R���z}�s2f�e�#ϥ�N�iVJD;g�@J�S�Xv�g����R�2�kԙ�$�$�����oj�&��n�)�!5�پe.r+��sg
I&����K9�$wz3���R��R�a��uwܪ��Q�6�:�����[U��+E4X�1v�~���4���uŶ�t|��=���*f�	�䐗�EyQ,��5���g`� �G4g`{v#�s�����X$j���_�
��=~o/��5�	؆B�qR�Q�'?�O��>�I;��bI��l�U@��Z!9��>#OyXғ?�T�{xa0� 5����;ڷ��Q��M:�G^��@���hEn�Y��%��� ����6����VT.��9���%)\�.j��ƻxP�"�h8�~��<Q��x�a�LF�0gZ��S�5���K�ӈ�`y[Jz�QW�ק�:�5|l0�����Aqwm^\˞d;i�M\Ff vE^xE���X�A8�4�(�h����������Kd���	Ԫ8 �g�Y���_��ǚ��������WU�r��L�|��9���Q�o��$���0>�s2fFC
��a4�)��x~)��-ݷʒJ��hx��n�������Ķh�� �VŎ	m�Y� ��XMF�#b�yG�)�i����<��3��d�� �]�q�����������4�Iߒ����3D��&���P�j?$�ta9�<m-�"D��F���b�P!�7��㕾��?l�(��¬#�����Ҫ)Jb�\�{X��}�&��!��M��Yff�/�
9xi��^K"C!��u�n�5E[z�~jr .�� c������G_�Im�f#S�쇈슢�Q�ۑQc9b�<Qu�Qr(_uNc�Y�Hi�h�GRT�vt0���7xF���f����hwV�~�n��7�Ѩ(W��gH�k�����ի����U���f�E�$�w~���&�}���r����N.�I��)��!ׯח�3
��[v��F��h�s��=�	2�t-�2K��*��#���[��M�� ���v8�S;�W��u՟����-�ޑ��@�!r)g���ƍU⽗�@Q)PI�UE�I@����ϔ����	�vO ��T�`��Dv'��{:�5W��	�[G�G�������v���a+��*���/�g�.�����	5 X7�m��Joe�%�����C��>�ͩ"1��ʋ��ß�i%��Ld����#������Ԓ���,R�Sk��R&R�.�'���E"E]�%t�����u��>��`��&��n~���D�2ճQ{ۻ�L�������>sd!�I�q]�R-��n�/ݴ�G���|U&;���[��8� Є*6d�?^��;N�9:��~=X'�ǩ� -v���)@�^� }Ĺ�B#����,ϲ2(�H��+.v}�3�ڧ$���Y`���gZ��ꐦC"��H���:��_��b]��)�
H�jdP�_�|�է�Ow���Wj>���S��P�WqƶV!:���HZ�&�vZ��V<R�Z�E���6�GH�c)z�Al����ۥ���+ �P���r��Bْ�%�ϚZR����H� U��d�O��R�GhZ1x]p΢_��4-�&R��rhU 2`�8������ ���C1��%�hs򣴥%S���ET��;.`���:��G�a\<�i˯�RO_��H1r�+^5�/��9��<E{��1BԆ:��>W��d�+ڠ��R qκ�q�m��:3�a�ܮ�c.��m�^�ؗ�ZbWz&z&��!��Q�~}�9������<�Kwbk�DL`L�0��h�A���|Ӵ�@�͉/�d`�1���X� 5���.Z��)�_��L3R��|��Gy�8+��S��q$�{�k��Tpڻz�6��^��x��/��q�T����XKA=N�������f�*�.IH�Zf�2sx����5����YH��V0����*Qm������Nwn���N}y�x�ӧ^r��q����VY9��dO�}`���l
��`�B�������)�Y���.�Ǖ�4G���b�	�ݫ���j(՘�q�s�w�"���A���Ϙ����C�Z^
�|'�AF�����3'� �R(>?�S�v� �k��;IbF��2�������X�BJB�Z� Z�02/���r�f@%��*m��mBgʝ���Z�ya��U�d���`R��R�����?�f�r�ݼ&z[��t��N������{k�Dr�w��i܅L�R�������	��V�?O��*f�R/g`/��-p?;R�S����e�S��J�+�K=�?)ω���ț��0��6[ԅ%���Wq�fЉ�b�@:����������F^�5�~���%@���S+����Zє��W�7���W����>z�ϫ��$^��]<��G�3v��R��O��{�V�\v> r�qp�|��c�pgd��# ��9��9",0�4�T��t+���3�)`0�]j���8��@QQN��F�LguB�V:��Iw�\f�O�t*�E3�/0�nf�U��"v�Ji:�돛����v7�:)Uc��4Isu�2��O�����Rk���:�U��=�ͽX4��[�V��t\)
��o[��!��#5m6)�}^?�Uy<�&Q�6Ř�m�l����e0ݠ��h~�*�]Y���z}�v�ರ�O��)o|7��B)M��[�[�wPND0�~��RY�����d�G�|f�|����[} N�hCb�'ml=1��I.��_��Y��TR����b$~KP�U=Q�"jn��` 9�9N�7INϓ)BՇ�ꒌoWҭpU'��Y^pܘ�9�_��o�0�iL��M$����1Y��r�T7q@1��v=�"����y���'&�T�Y��F�9d�͐���sяl�E�KY%n��&<�_ DT��j.�3� ��:������t�|������}�Y܋��.$����A�r��IibR�F8�7 �Q�Pږ���'p������?]����pƪ<���QV�J�q�$"VU᮪6	4��
(|N�>�ܭ*X�<u�B��d��,N_Eyه�#б���"&��^��jmnK�ed�-��C7��J�
�}�o�R�:�9�*�f��������w�.8���v<.!S@ي���=1 9����(�4����b�+@����D�:�%�o������R8*(�恬u�ٷ�U3�z�	� +�"Sx� <I{}�"-H���
aB)���TD�ې���s���A���'�/!�K�[����?̩��9���n���G���J��H�)ְ��oR��<i(�����z��)/n���DD��>�nP���|�Ew4w��#��i���Yj�Ћ���î].�%�>��`�D,b����$d�rpܾ8����%]������ͽ�Bc�On��0�!<\�B��4�,�F��0h<�}�%a��F�iȌ��,���#��j�ڐ�n"�9���׎�&���q*���;�Yh�{�8 |���Xoa%!�BA� i���pL���v�[Ffw�������;}	8�A�sj�^��і�J#<B�=��9�yH�/�̺�#'�h�=� qW�/����;,dZ�`��?�l��0.n
N�u���Q}4:k�7�s�J�j2R� �aHA:��ï�{��'�=���+������
�L���RRx �����������1�~��*�z�%
vZ�"1�
=p�M�=��7�2�V'
l��pi�~��5!���m>�D8a-��[��8cB�m�0a������0��d�;�ь�,:(�w朱g��o�:E�W��x%� <<_�g?�;�V��p%�2���7�tiU��f	�	&Oj�Lo� �7c�%�'
a��b�`�U/#����T�t�$>�5�kQ�(�f]�/E#�����z����_���ĳ�"�1��f�BW�C���ޅ�� ��� 1��[����D�6^�&V�u.B�#���D��,�ҧ	��N.(NrY����Jxlko/ �6R�������w�mY<��ś��k����Y�n�⢸˿��flN������9o�
�Ԑ0%��r��ht��+�s��W�xn��h�8+1s�.
�����>�	�^rl��((1=��~��:��v�!(^y�iəʉ�
��r�J V㛾��%C&�u"_�q�ޒw����1V�+�厶ڙ��Zi)k��^eݛ���{�+Ӊ�����c_�)�i���Ül�zVtE.��Zcz��%W�^��B���)ϱ�2"p��u���u2����-�t����Y=�ZD[?Ga���lw�n1��mmc`�"�4�޾���ON�&�
1�G���"�9�:���HE�(�.���ꪑ���/��R����@������_���?�����»�ƕ���N4����^7�Az�~5sE�y?��J�}���K�� Z	��	҉t���FC'{pt{�g�E�)gu�;�-f]o�M�مJ�<��S��/���KftuQ�U��Ѷ�9���ޒ��q�����˕+�@�z^uL���aJª}$�3�;*��������u�g�̀�FP�.X_E�YY�㭇f�m��&0��/d��Yf�^!70~�5��9���S�x8W��AoB��3c��W���ޫZ� �J�,k�$����l5�F�k9��.�=�B�5��"��&�W��	{Ϣ��6=;�!I���OJ��
�]���6B�&w%���Uh`5J�gM?F�49���eQsE����!�!h�Ʋ���O%F� �'�Fu"�ż�5��	��=yo�����P�J@f�7_���0�����:�!�ZTDc�o�ĥQ��ż�9�?��-	wu]Ii����՜���&)�I��9�-4hO���ɌeBt����Şc�g��K�7ڶ�����4a�u1�Z�P д��e3a�n��8o\��]d���{�{� ԧ1��pJA
m)d3�lm1چfgI\T� `ef��m�D�!�3�C:,�cm,���V�;v�[�X����l=��ܝ�wzv�&"!�ц�r�s�(s}� ��2�`�M͙#��z���J�@��X�\OD0�`��S �-��Gf8� �+����D�*��O@N�����U:�ruXowp�ws��!�ζQ|��n�˜[�� �U�E��R@U��78b.jB�Li��<"r�������Q��&�,No�bw�d�n m;Dą}{m�2��L�АXl��|}k8�~�q˽��И�m�t���<��L\b��omt�Tð�`m>�>8 �6��~kC3������(��q��j/�X�*���Йao�kuC����lW�0 �F�>�~r6�tc�r�u,}��P�|9*c4��j@�t"��Y͂�w����v����:�΀�uV��Unb�K��Y��������Nָ��ӣ2ݒ�)�<j��X�k�a[��Q��Ay1��-i�~�y}���P4��{��4�X�F���ʀ�]H�%�N,�0���^�� ٮ�tfu�#���7�n�ق��e�JxY�gR+6�(]4�L�ڂ��R��> 	Xeg%d�.Z���Kq_ŷ�_
|�i}��=h`�u*�kZD[�(i �G.Pqu��p��Eq����&)� ;K��d�Y�o����qK+cucIR�m��%^�Ñw��3�n�a�/��V��h"��W{�lm7�����*m���G�ͦ
�#��0F������6ظʑ5�:���& ���O����9&�oY� Z���`�僀��|th"��)�O�B#�KF6�� �$��1*i܁�	O84���U��t7����S��^8d`�y���?�i�(�����S�|гEL��]-�'�>�X �t�����$�@�m��G�$ڰ,3��0�$(�B�e���	EPi���`іt�"�i=�Yt11i�ŏ)�(S쟸B{=7�3�B�כ!�gJ�][f�ěh7�mEO���.�
V.�}�)�i�;��k�jΉ��}E�]��NHȤ�C��'�KĹ �d�s�(`ր[3'��,��(.%����T���Sm ��E|y3�ؐ�sH�nf�ss��*��Z�����Ḟ׆t���!���[�
���@���!�N�.�X-6�̽�/	Mu��#�T�>�ӂ3c��x|�QFo��%K��X����t�ݔ�Ɂ
���cЬ�BF�{�6 �r�])�=og�c��"���t�_�h$/��!yg��$�P��ǳ��B0wD)0���bo�m���#� �d"X�h"��@s��TS��&o�e�7y�JȪ��JDI�;m�D��lb3�O:�vO%<q�Z7i�Bw#�d��)�d.UG>��9®Ń�HBι��U�Q-6�xL8�'�0��*�+C��_�2La���HaW'�_$����~�����ZH�=��I�}d�h����n�!�����g��R1'g�S���}5C�^�n8�dz�یE[��wιa�������-9ө���Dۿ��k� ���X���OHƮ����r�i�ȣ��ʵ��xř�|v�l��"���2�L� �}}��	�)�� c��IRm�h�UI5殶��8	�y���?��YZQ6��/��5,����鏆�Z}��1��,�m�?��"~��Gܡ����dI=j��:�xP�?.-U)CE}�)�pf���l`�Z�^h�ű��=0v����?� �1Ob�%��}a�}�������g%F����G�\*4-����RZ8[�{j���/��e�r��RQ��<�<��]�b.U>i���ؠD��3�<7��qڏ5��4B��p/)����n�E_;�)jN1�s!*���3���JW�d�]Z��C�ܰ�H�>d��\�YF�S�N�a���rM�j��8���nhLk��p��'�@s�5K�7��V%���7�'G�,�/�0�N!����.UEb^`����ܹ��peܣ3��o�[�
�����,�3�xr��@�����(} ��	6��##E��/�l�����Qۀ_E^�7�({�H��|� ��(���>�OkZ|ƘZKY}��p_z��I��pps�s.$��*���ʒ>*F��kChRE���Y ����^�~���Aò\s����å�Jb��?G��s�w��1E%rkd� 8�)�ܠ�S�r�1�8�2�D��W��Mod�^�'Dg�V3�QF�e(jZ�mx�SS;6z�i�����椂]0w%��?���Z���nP����AB��C'a��~\Gn��}G�B����7��0u� ���),�o]^�5U��P��o���:G=��������L�c��&T��y��M�����'��ϒb�tC�^aQ`D5�4��U�U��F����=�R/����ꢚ�M����䆂��XC�dJ'��Vd+��sX �mqەp�r}�T�/I�|k�$��M(��H���=4~|���K��kF�2��Y"�A����~-xۓ�S�;0��+�
V��B���Ș��SN�:�좋��P%ío��Fy/j���	�d>c�a�o������N�B���2��T<R>��_̰p!�f�e`D�'di2�p�xL��|�Ϩ�M�9�B��l$\���O�+��T�I�=�|��< ���o��ٝʈú���W/�n�j�U X�'*:E_�9�~_��Å�����Hi�)(��ɕ�#=B ���<���"**�u7�|k�.,-�|���ai��[��©��D�	0��d]�6�wA�?j� �{P��*�E׾ߗgP#�hf���|dh2g���5�	�U��s�xR3|.�5}�i�G\ѭ��Ҏ�B�e��u9��*A�
 ���f�P!2�=\Wj-��I5V�^�9&�@˻r�}NN�N�����0��6k�8	�bV	j}# @��])Z�	τ����0l������Q}�I�}`@�L�1M�x�{)�3�g�>L<`�+�c�3
��s�\�q�e0�4�����S�2dKFW�J~PN��,LעŇB2��J3���ɷ݆�.fu#?n­���w*����8e6?x�Gf����429�>��Qg_���+�D�7�(^��7KÛ����ky[���u�c�<R&�[�7�M6Y���gh$�I��ݝP���T	�p����<��
�*X>���_�l�\I-cqg(����7��+v_��4�,�^�F�ρ~Qѓ0��{:=����E0���%���Ԭ��,��S� ��х���hot��7��)�'Jz�x]ok�%���
��/�;�;a�#y�����|c��W7ǠQ�$�c]΍S����s>ң����P�t�gG�n����`�exe�����@��� z��>,�D�$���-��"R���]1�0*t��ŵ��!�A_ϰ��7h�ޕ	��	���XD����� ����*X��=�]�m��ff���t��'|L���}8�Q����u�i�iN�r(O�z�����|��"�Xڹ^���]jb���yl���d�y)e��L��������}�k&7@λ.�B:���s)\�F;���?"��C~ؘ�M'�D�}��l֮��r��c@���1�S+D�a~��UDʕN��*&^�Q�}�~��-1������JK��ȫ�3����*uÂ9���O+V0���|��h����fF�"�#�I���qU�J͍��G=P�jz�2G"���eo`�e���[����&� �6�6t󈪃A��M[-r��azkt3&Xw��R�<7���r=�D�ez{�u���2LKR����D8jwN���W��.�1i�0�a�1��e�S	����F�(Y���B����f�~Kkga@�XM�(��S�Y��Ǽu�.���H�h��,&���I,�Gyr��&�^��B�!�  M³����e��
��=�`��d%8@t}�0&��<�H�ݝ0�ԕ�l�[{�U��_o�(��f��VN��4�7kSp1r������������z܁�V����E<�>0�J� o���^@'�h��<�׋���G�z�lW����� �м	sRՂ�&�[),���	����r�`{m	v���fy�3-��W��AI�:?�Uk[�=�.[=�-�\�6���*;�ܩ�C�JE�2�i��I~<o�qW5z�*��/5Y��.�aM�
��L)lH:��%��0���|�oZ�B�w4�X[7���s6O �]�2X2���y>D"�$.*P��)�q�FK��'���`_*����/�(�t��}�Z��n�u�B�m�:,�<lЪ�\��'�@e9�_�.�k�o�W�t�7��-Ӿ������=�,w^���	�GM�q�+�"�����K n�}8����9�Am�o���07#~��U.;��̮-2�p�Y�\���#d��&jv��>sy�X w�J�]n��v����x��s�g��N�S͗Y���n�S� wIy��C]�]���ĉ�8ce_}\��X�� �E�H���@̚VA�j����!>�W��PU��}�['U+?}�hLΚ&gWȚ�F��Q����h��*� ���:&���BwWl���o���Td��'	�ʣ���'p�o*�?��ytP4�����5Y��}��ø�M�ր?�`�55w���P%'̔��2۳�T��ltaLR��no�i-΀�Zl}܍�	���,dqL�n����t�KS�|.��%����TK@�C�=�GRV8CoP�-��&��ڥ�,�V�c4��xYL��~��zDq�B����}dD'�&Kڣr;cy��lk'v���܃���l��d����ө#Z�P���h~�zj�t7w�u��޵��6����>7��)��v.B�\ܤ�0���I�[hl漘�|��[���xb��&dj$�Yk�-����5�pr���q�Pd���0XN������tZ�C�T)�����3�Ҍ��islF�[��GK�E�/�be�M��H��p>-u�v��Y4Rز���^���������BE��Y8;2�-���:�$X?���-_ �YB�m8
���?�c�C�w<j����k��@��^N�|�
�\�����A�([�V뛭eV��M��%5R���$��Ot��&����gUS,�O�N�z$&cȥ�F�����71��C��j����q3R)����\�"�����_%�3Q�UT2T�b�P'�2`�P�u�Uy}��(�|��u�������^a���>T�P�:#|M+вJ����[H''������v@���4�z�a��ȸ�wR���G��<���F-�u�p����3����	�I0�y{����.��L��%x�)������\�$�p�e.��9hjŘ��S�(KW��Go�C�"���$G�1/�k���T�Kc�1�Վ�7�2��W��Z��V�s�O�'#�Aŏ��Q�_
V>�9c �GNl#��.����B���-���O �Eg�F�ƚ�^z�W_�髇~ǋ*K�r���!�X~>[�4��B��AY�Z�(>��S�T�8|A8�7��K�lA��'���Ѧ��$p��\3�b",���qw�,S8X@�����ϟ�i��[�K�4�+�
��XI������������m�DPA}��_`�w���U�A���_�y2�Ь����t��_߬'	i�c(o������ݹ�w�0E 4~╒fO�l��)'�����'n�3T(�'l�?M1�vgI�a�*�4���@�']�[�b�
l#_�Fy�p�����㤛7 �E���>�y]��>�eJ��������Ta�D�<�l�9�V9�h����@�A6<���?��,�M�K9qwND��D<3��B�E�+c����Ra�ǽ��ס�N�T�3*~��T�w
��g��f�d�����Fg/J(!�*�̀R4�Ⱄ^��g$z��B_#���Wo1�Ff�@E[���~�&��	�}p������F]�\�_�1��d�mHNs�!ۥc=���s3�Ȭ��o]y�a�^ĻF�3N�y<����|6d����߀�z�}�����xꓛ��h-fap	V{ 	>�A��G�{��+�[~��{2�i�M5�R��S����0��<�@ŗϢ28J^���gf�|rCv���;�j5p9����+��nr :�O��h��(�u�� !�L�Թ�v��Y���ί 誮@�>yv1yu3�ē,�X\×J��9��w����"!�WˈDuɉ�� N���>^6®��h�H�@��O�#�q%�'AÁ, �~!O���M�bl����xV��1�^ץ�Q���B�	�����
]f��B�Bg_҂�=�U�$=�Gw	��c1RӷuA;I��ߙ����ooNo���|
;��9�t`V~�"0����V�Njxu�3�Ճp<L$�$��դh�"@�f1$U^�al$f��d���`�=L�mɖ�rY�v�~��BaE.��ػZ�Q�[�z��lo�:�I+ƨ�!�o��
���Xl�j�VJ9N�(���'��D`Jk��ڹ��?^-��[��̈́0�Rƴ�-?A0#��O�~%i7�j7�?��x=fguv�iͮh�'	��-���gbq�?��	~ԓ+���R#++����c󾎻��)f��k�#�hl�a9Vc)V�� Pr呔�9T�$jr����^H�@T��QF�g�ୖ���D�ہYW5�c^�U��)f���@����.� �j^C�Z�7���P9���-2mѹ�g��5(�^���
�W���pXXV:���M� '�HB)�q�����6\�(J�;w��և��ӵݩ�y;箍*��oB�o���vX����E���J�K 1W=dF�Pߣw�;o˹�/��>�4]�cȘx��;�#:d�1��^ߔ�6UQ��n��V�<�A^�R�l*�li5��7��̜�.���(����D�ոkvi
�g�F�F-��mwH| ����E�H(�"� }~&�V�I: �
0R/7!�<��z�vy��{I�aN��q��
C��=E��iL��|��%�VO��i�x��S���:O�/�6:ks�e�}�|,i#R�i��{E�c�y����R#J,[�A��#N�3M�C�&�G�O,��Cy���S+�7�(/r`��n!�ҿ������跕5g�U�)�Wp7	��x ��Yv�7�D�NI��і4ة01J�6��l",V�z|�Y�8LƝ��{U���+���__E��A�¼�E:����6�Sf9�:��8�u��O}�Ĥ#���yWS|<*J���`�Wm�=mD�D+�q�ό�)\�KGO�Aa��A
���m���1�y�+�Y�#�̒/) g��I�0��6�|�L�)�l|a�]�����s{�}nf^���O&��W8͔�70R�j�Y\�ZކDZ���A.$)�f5�]�C�.�P��g�������v_˪� ��������
\�*(����T/2u�XJx��h<
��Q�'�?(q�cR��7���<��Y��������k�����FHsgB֥%>Kݘ���N�|r�"�'�"7aQ��P���q�/=��j���ћ�e����ĭ�V<�H�����W��{Q���j���o�9��j��QWYӏ(a�Y�a�zf�e%5^��㢐(ֶ\UH����ޯ�Za���8���Pw��BRX��A��K B-QJ���l�k"$�|�/�`��ʶ]�K���͹{\�V� v��ٳ����R&�N��іs�
(�L�8�\}�c�+�T���t)���䥩��#�)�J������1�a�6��qsoVK{c�\Q���Q���e�KE�e�p�]�R��)�F�6^ ���!&MKh5�7 8-�X�Oh���������m�⡕�V�9��)�z� M�a�,�i-�3�s>=��@�.W�=ȭM��Ya���o�1����̨i��t�o��L΁`^��/���8�W���ӆ�}�;���yw�rz�p�l�Rs�.�1�|��q�Kc���u}q�v$Fe�����R�3ERF�Gp�S�։z��4�߀"�?i��E�~NZ�_�6�RA�H�� �ukuy�����m��S��j�@c��Nu��I�}xj��,j���%:�p�l��c9x�Lޞ� ��{mq���A Y��b�x�j�GŹ-�XQș�E����(�_h�%e��K���d�g8���Y/�0O��:\���k:�s�sZ|v�`�P��>|����W�m)�w�b2y	gx�H�6�j�G5yW�7�YR�����#��HE�g�7��X ӑ#�B�=�;}�OO�(ȷ���(��S�=\G��I�^
���M$�]�\�'�C���76EѨ�- %DH&Y���I�w�FO`A/��T�W{��/q��^�9w-a��
rk��L�S e�e�)���
�&0r�]�s-P�#��0��t?&�0%�n�
�Z�a+L�UA�&��h����pp�;��:�feU#0���z��d��j�"2k��7��hm&p���2t�$}S޿yrw-'B黩��ԩ�[�K�����.z�Ȭ��Ʊ��-���JpDArp�Pt��.�_h6���{c�'��B8h��� Ӵ�Ε���ct�_%@��^�9���}�l�\S��