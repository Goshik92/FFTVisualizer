��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]���t%�Q6��i��`��B];>r� �m�nC�2�������N� 7�۟-�΄e|�,Z"sM�DB�n!�o�r�[�'�F%�i��Ɩ��I"Imm�^ �Ϊ9#��0�0U�0�� ��Dk���i'�>��{���XQ!�%]�,k��<�VѷA$6��`��3����()�s ��#w1d�#=Ⱦ��]'��z�'TG.6PJ|�i�iJ���!�3V�6ښ��&q�s+*�����"�� q�,;�"a�D��y��P~���m���Rj��0R���^Bɯ�Z^[������ݷ�S�<��6��Ѳ��9
A���ī��_���-� }QSBj��U���߈vL��/zS�����R]�5�]6��1���9$��V�Z�v�8�B��:0���3�f�e�j$ԿE�|�K��1H�ʝ�C��;���r�|���ؓNYi��ß�F�-�d��I���p���yg�e��+?#_�q�L _��Ari���}Xi)v�茹�ԏ�(��IG��0($�����Z$��j���)��]"pa�u��S8 r�p�m!�d(����j�|�En��GO�&��J�녮Ɔ�rW.1���w��D����.�}l(�g���{r��V(Jg6�����ġXL��cjis�e9�lΓ]z*W~Q�͙4��/e���6�=c�4�Gwlʘl*�tD�Z����u������޶�NS�aR�J�	��S��tF'ޱ�E��������ȓ1��~ɩ�\��߫9=]z4���U��k�{�0'��t�ʼ���5�'ހ������#�o#����0ɜ��[΋yh7�
�ߔ~�f>\%����EF�
2=*f��{��U��%1O*�Zd�[c2�)�1<�<w^�o�c�J����Q�)j�;�Oĝn�Ff?<�ڛ1��[��U���چC�$Ǔ� N��\)����q>U ��b.�<�Ib$�M� �!���+zU�(��xDcDQ���ז*�QKU���w`&��M`�)�6����be5K��3��%U��]�8�\?}�@^{}Ҥ���BkE�Ew����7�D���_�~�dLT-et	N�x_~�]����[X�o���qC�_Kl���Q �P"4�u��h�3�K[>�fkD?#&bE.�P`��l*�,�r�s$)Ju��n�>�J�d:��a;��5��w�h�\���̰���+����$�·�*K682�S�)^�wb34&��U�X���$�M9�G�	��O�@����.z��F�X7���OmT����Lm��νe��u�j/���[x<�u�ަP�,M��l��wE�S�K��j ��@��=6Iq8�w��7~�/�j��M���*K���#��f5V��\v(�"���k�����xw;��܏����.��y�����k�S��tK�f�8��/�
$����c����UX��9%��e��	Qc49�ͅ;����ZI;ƺ����'��8@^~'�������
46��k����6��t�P~�6��^���/6�3i�<��s�	�w-d�/���{V���*w�)Xf�B#��f�0���!�#�,q���6�wu���;�r�]2�5)�ޢ��+�%��ˁ��y0]@�e4|�v\�5���}���~��,M]��A��&��q�o��`��)�EOS�$s��T��lF���A'!ov�"k�E�j�u�fQ֗/��E��dJVb3����K��ÛFgF�ZX/�*x�_R����9�ꚭ1����L��0ps�df8�&��y�����0恟$z�Xoz�S�'���U��NT��Yl�I!V�O�>��N�+�[�e�x�QҜ��i� Y���:SfBVo�bݽO�w���RPe��4��'bV<d�g������=��N"/16U��9��Ia&�7��L�)΋B��Tm68g��Ia �)�d���:ֹ���֌�l��Ro�t��[)�9�f{�c����O���C��6�18��g��ȓ H��i�E[�j��J�I��+��!�Ϣ�
�YE�P�ڛ����L���^a=H��
s��8�|�W�j�n=�V[�B�p�$�ۥ����o�@-�zdPk��,a�-Q�S!����3\e����N��	�!�!�z�z��=��Z�S�d﫱���h��-�W�&�P��?�ί�2�`�*�Bp^�l�j$&�@���SӉ~������bՕ���ˡ�5�/�o"�FH�1S�.$��5]�s�}\����`�z�#�\P�Y����TѲ�ڛdn�`��z�jr��`���c#��N��^�J�W`�d�.�v0~�?��8-��2ޣR,'�37&��\��e����<c�+⨥(� ^!��?(l�a���6zz�[(���j����굚(5ߟԁ�["Е� ����t5V������t/3Հ}?YL	W�[*�3�SM�ke�:�t�������OA%L�
����w�3����D�~Qr����؍8�8PRS�])77�l��u%��.=���� �9`��?k��bw���E˖��}Q�Wo[aG�ث�N�E�Oz�M�W�h��MKf��ty�<�S���*������i�^�p��_Oz�?�^órK�1�uW�����?��2c���E�����2[����q偼K�\m'��F�>9�ԉ.��ޫ���M�k��1���G�k�5���'0wPJ��ńZ��͜E�D���3@�_]�o�d����?�re�H��m��Rvڒv��{���;���<�a����k~�W�H�����O�����\Vz�6�Ps~Z[z�=@a����"�c�.���o"ʽf2��O��~����T���'k���X�� � W�7�H�a
%'*wډ�md<Q�o�G�?=|H ڛ@~�:)+���y��m�~~�M2��L�*O|4��Ei�
�+C�U.T�?;h&�]L���'��'�i��Jw=ى��#b�8�,�:.����n���0�l�i���`�Q@�P��v���g�����������/��췾����<���b��ɘ���N[�aO��җ�
#�4+r��,�[k �ȱ�Rc*������b�} �i<�g�r�uо�2����0�$L�W�㏡���@�hkYOp�oB��KN'��/u�zS���N�/�<�mg&������
Lc.��5� ��Ín��=KY ��@�����e��#ŝ�a��T���:�ڤm.>��߻�F�$y�y���ز8W��hP����J�Ѫ���zA�4������=,S1��Q
z[�X���Q�L�3���*On�S�1$N���DF\[i�*�U���z�R~����A����LI�� �2����-��T�7�_�F=�}�XeaW�J훉8�h>[�.��@�ؙ�Og�/�j<�����e�~��'��7����D���(ۋX�Z� ��@�Z
��1�������O�\8E�ꄶ3,}#�fy�=10	U���Z.}��I�cj��M8�j?�2��"J���h�a���l	p��V&�i�q\< �v����Am����E����=��݈��կ�����o�T�jmB@���N�����1�">�`,��a�@2�ҫ�l�U<���	��M)�c�|>��ҡ_�Zh�Y?��1}�k��Z�����n�<u���dfI�N}�E�	����_;��l����>�[�y_(A쮌fWt��M�iWo�vc��6�P����k�p_�#�xR/���Xw�b��AF���*�{ɻq��C����3�^���`"t����I�/̟XWP�҉�&
A��ZD��h40���Ŝ*��H�-xm�;y���G���N�{k14RuOgN���w���*���O��R^7�˓2���)}*�/�7�H�&I�Tg^���&�Vu�yڭޞ�>L(��ǔ�'V�=�/ԚAy����V������8u�17�����kbMLAs��`jp�s�ѡ�8(鶱�v�\U&�ܨq���l���zx���V��I�1H&1�OykJ|�b����ߣ���
�7�7�~+�ꛁ���"ȿ^�����m�f��!%��-���u�l�P�T��a�M�| �tH�y@���Kq�u>V��	Z��G.XA�)�9oAP�^eA�#���\�P��y��9Kɴ�2���[x��F���,<u���7C�N^��ne숛�é���qW�d��B&�[5$ئ�X+JsD��z ү�Wg�M��U;����S�q�FS�S��<��/zFvP���^��l��n"�?m�p�##n��[!�:���#Ҕ�`��z�g�o��#P8�N!�C=�%��4adI��&�p�ɶ(�7�~�&�E'�(�.Xi��:�*H�4��5�1�>�Nn]��no��?�V[K�F;��"߿M� (؀v��N�m⼲���y�] ��)��[�n	�X�P�]�X?A:�/���m�>O�pD܎l��5(�a�'x������`e��agw�X;�<6a�g���� Ҍ���Z9��C��L�
C[�������{��6�K��p�Xz ��B��/��������S!
�jrI���%jo���mTBi�.�DU���O=y;�MHKл�?` ��/i�~n����leܝ�?f��؏Ѷh))���֛���^��
�j��n���}�}�}���K6��f�:��]5���tۡ!�)znƎ��;u�<��"i\�C�y�zc1����٫��
�s_�'�Kx����8�.�}����Q�U�ik��1�-C��O>���EF��=���w]q�!���h�+�{`��ګ��E�U9���=J� "a�b���?q��.h���U���ɋ��AA�1x�C]��g�6�*�1��ܘ2΂cl�������l�J|���.mq�ᯜ����[�i�k���o�f"W����8x�"���[�"$1Q0���Z�4 ~�'8x���J ������d0~��j��䧫oz�v�3�J��et�q�D��8}�>}	��?�}B���h��'��%���ոd����<��b�Z�Ek�%G,H�?!n�U�V�cbA%�C��s+��l��{���G���vh.�	Y���7�о�b�G^S ��	�	⽣BQd%�^
W�x@�����v��j��H��DIL&3��Q�E�������)O���ӽ��-�����⩥�L�Z�$��VV��
᳾��,:���o�$���ܧ��in�X;��!�}��u+W;߷���8������pW�iV5�YNU�Wj3�� �Y�
���vq�͠0
H8��`��^�����կ����^�Yp��:��	��U��}�Xc�D����D'�`�7����R2�R.#�=]�� i���　�K�l�d������pⰇV�D
"�ugJ�n��	�V�۵���gG3텈���b��'�	�T�Y�]�M��ݞI�ۂb<)�{��G�%�\��\
P�K��.̫Wdfё��i�	�&�z_�R�1"����=�b4�b_�͙;.ڵ;�/��>^,�i����;�F��,�[��4a�P��)y*�^�R|�:�H�F�hg��1&o3�D[�e�J{�g��*g�a��m�����_�$��sY��"m3!�i^sUJ`��M+{�B��Ql�|��>��-�*�^�%��#V�L��g�K bxL���C���D�Gj	Y=E�[M�$N1��%Vyk"E���i���d��O�J&ۣء+��m���,/���񭿣�3����>�	�nos�K�:��'�wQ|\��\<M��S��S�=��*�-���Orb+W�v�P�� u/�;K�K8�X�R6����Z_c���p���A'���^�Fwr���w�(���?��B�1)��ӂ�h�6���z�,,?��*��"_�^1�}B�nDla�!T�"w�'������\�.�F�����z�%��A��~��!�ЏJW�K�9+���_��GU S�"n��e����=q�>ns�/��Ah��F~ϑ�SYX/��^,�9�F*�r(��0�;'@��F�f�F����h�y��+A����q��JG:�b?�v�^ն�-��ԈE�� y��\.t�����E�,�C��}�n�u�<3/�U[W�9d�c|��	�7�m�8ڤ�YDS�k��K��K{��G~�l�Ĺ
y�1� �Q���BJ�!%���.4�|h[�a�9|V
=C�4�oJ�A���S�Cm��y��r,R�'�	�hb�T �rS���;CLX�.H�6�\������3_?�����ϸA�:�:�?� _7�i�]$d�$�����%|P=<B���`���S��6�����p<�4�Xf�h٘7�V���s�ZHR�i�}����e��G�6�I-�
3�=��U�&�#z��û��C��p5��D��6�?)7��
W�o@�(�) ���^�_�5���n��V'�DRb�I��sU�&&Z��@�V��qy��],&�Tl^L�IO��r
���8Y/Z*M	(M�|b�odt`�X�Waрgᓸ�~D ?&��]�F��-+��	�zk@�8/��%���@/p/B��������+���8���\�<�!���"�;��(�����'FHz􍃄�6���.�}=, �G���q�,vߠ�6�^glD�b���o-�N���a���-nj{��?;�)�R���	_�I�{Du+h#�l�lvc�0�Om����ht���h�w�0U���2]bZ㒉��B��ej�F7Yw�h
��L�]�����A�c�B�z�t:]V��� ��8F"�p8)ӗ�Z�ItC�ܕ�n��hn�VP���mGl��������$S#��r�צC�=C�C��\�cԈ��R��N˶ea�%�4D���˿���KG���p'N�t�<����7A�Q��E�5�r-�lb����p���U���Z�+j6!��{؄�fd��D�>�U�aЈ�t�&�Y��M����Q���=|�����h���v� ;���c���M�`Q�������K�U0.ĩ�wEF���Z��^vE��<��^-"B�%��kS�L�o�[3�S�����ܞw��9�t��j�f49�	�=֧-}����%vc���U*b�J��W;c�@@MeS!i��+���z��%�������\���v�D00�.�i�B~�T Њ���1�!��U?�
�d?��|)�/�2��XH�K�4��S��)]�|�9�H�YG�=�qM	sR��X?�"E�7��F1wY9M'�5���
��
����d���K��1����hB(��o�T���F�A��>�z���^�����׌����i�\�C���.�ƅg�n�H]�r^��6�r�ZŹ�(��>��X4<*oGg[����-�Y�=�-�<,4��n�ٝ+�YfІ��'%�لl��u�ig[���=�a���gޫ1�V���P���aAPm��Q���f�/A vE�]�tj��#��Z�0�5Q�>i�YJ}i��c�p83�ï!#.p\��9������ z�04��� ť��OW/�<@4���Z:C85���^
��A�v��=��;y�ۚY�z���:��O����#u�cnb�6�e��3?�3�8I��,3у�ԩ��20Iؤ����a���K�g/��$�5-��08fVs_]�u��ѩO��̍�s��ܼP�z����۸qN�o��?�>TmN],Rd���~�BD/3��9��a���ې |E}5������h���'�����q1m�p'x��z�050/�6��?'T�R?�t�J�ˁ* h���":�(��i�
\5T�Q�r!Զ��)������bJL���Zg�:Sv:)؋���yL��}�0��]Ұ(QY%f�׭P��$3*4[�7ݛ������	/.��:ە$��@�ux&�	�D��l�J��Bv��F@��_��J��ϣ���(1r����eŶ�9��:�Yx���Y]�����;����9��o\��w��4yZ��6q�D��������:hr���%�\9�6�]Z��~D����a��k� _�����s�����3ݶe{C�#��
�����m?���=ρ��q��s��=��#��:MX���
�<3r��_�w�з��_YY�s�!B�����)�\d�e&����1��@��"��9���"�0�?t.ә��	7 �1J4��?˾S�v�v	:v~l��U����튒���Wx}sI:h|B�q�7E����_꘳��8AĞ�!a�7	H��UQbR�u���m��j2D���ׅ��7�rD=����!��ɖuׁa ���Pr�C����e��Y����%+E���.N7�#�k�C��������/���Ί���{���I�D?䔥�oQ��%��vkPƊ�1Z��e�B���F��y�e�T�,H:�5X�7%��y�J�0]��O{�CD��)�S���)��^`�}s��Ā_���T�mbk-�<�7V��:�Ѫ�
����©��;Z��f���@����D�6��*8.�0�&h�&!���5�����E� �&m�IK$��B����:�:���Y���B�R1>W7+�^[q,��M�<+u�j�6U��gƜ	,�ҳp��o,۬��+���w(����p���~xo��L��צm��xj�d��r���V��cg��\�u�Y7S�fp@�{D�8_P���D:�l_��?�8�d���]�*�CT�Q�:�E�󃚁\�}�
�Hۣ����R�j�,�y�xx��Jz;����P�y)�m�g(� �I��N�"����꘵�GM�틳nt��7���u]8���=��ZD�����0/�9F� ���-���;9���6ߤ��5���j*d�c��ӳ�mB�����ZϜێ��*�m�%��`k����N���U���� ��ϽMѽa�%(��I?�����ɫ��d����қ:.�V®Ӏ�Y ��D�O@d��_��v-�aE�	�U<C�m>�.����t��̜��e�sYKڟ,y�z)H�R�gyђ.��EҞȱ{ğfHI{ڝ���.����#����-�9}�+-���K�"<���z�}�_��ZR�y�y��3�ԇv��7��A_��Y����1F��p�a�UZ��������Fhy������|Q�F���k�&��N�3i>D��<F(� �o�h�xֲ�t�X�]r��M�����f����bA��6��ק�ƍ�b�gR���Ɔ��c�W4�����,�����F��|[H�$2؍jc6E�z���Z� A���ۣ�!8���\�����Z��R�N?�&��0���G��F��LۚǕ*�����#��B����O�<}�@=%���5���͌M���C�x����6�t�jb��z4�ɓj��JF�9W,���K�]f�K{�b&�7w�1c����:Z'H�?����\�0����8?�8uG��$�8p��b1e_�*/��"��((j�c��z)ߏ�2@	7��"W�Ê�	��H4���<�x8�)e�������0�b���ж�~���x�aO���׮�3e�j��S[�ܿ�:z�/�!�8�{�b��"����C��:�Q����MP��ӕ�Ϲol����;�I'��$׽�4M�+�FH�Gr[��S��Q�#8��mY�R��-̡�3����eS�$k�7�D�W�6˻�1c�oH�	#~���K8�O��d�0<`�����|v�zI;Aαʿ�s�ݴj���Q�B���6${o�JB���cߎ�i��b����p���&��K.�Q.�YC����k�eB��q���vN�Б��a;����l\F��t�����{;���b���^�w�!6v�<�|�����"���U�B�Z�g� ݼP�(
�l����F謣���OO���x��xҾYwF�o*�8�������u5{�?��,���q�A͔gC��ep�=|m��:当�6��r�"~H$Bփ?4�cI��t?/6^��"��$a�,k_Q?��!b���M�E�OfeK8g�Y��hrem�����F��Ec??�F<"V�J���x�Z+�;Ѣi�"7�j�l*b�8{��72���(� ��V�D���?��
F/k��>��.]x��,�����.k�cy�Y]�ͬce�ʂ�'P��#�FІz2����� �vo�^�tN�FU��+2pK��E�*���_͡j=�E���0�`��d�a��C��֖��L)�����m�=WK�`*�Xv�@�N���A>I�߯���b6��t��p������ŉ!�׿�<j��l�	^P�B<Sa�׃���E�#0�,s���y���/��0���I����(���0D	�I764$'z'
}a%��ҿEqb,<�O���<Bڱ\�lϗ��-�)-h%ߖ��x��J�L\Y��58��lM?r�ɟ� ��zv��yV�>�6ҝ���x�Lص�J�,�N��i�A~���o�7ʈ��Pi�a�."b��;p�l�=�P��n�
�1�?�vmRxK5�-	3=��|�m�n�7��Z�ͨG�c�x!�Ͱ��6`w����evx����7���>ԁ��E�S�L�-'�e��y�>�.*W�k��Z�r�ְ�#�"mm@��.Is�y�>�0ղ���h�/���o!x�r&�8�D%�%��6�@��{��9��b�s�&��u�NLR��ϲ�exC"b� ]�]����o��0�_P���M�{E�!��.>H`�~�)Y�v+H�F$�c�Z��$���uXtqB���gx�OŅLܟ���h�x1܍�j�	�G���*C��_^*�Si�^���?��^ s�y}���?�YK�V@V?�#S��m˚�.��j��:ҷ���[�T��Cf��}��:�"9��CÒ4<l�a^C�A���ϸGjL���s�q�1���RD��(�k�a�[o�Z$}s�%Z�O��6��nu���4p�b���C_Y����D�ؒ�³�Z#�m��ŮI+|$��@�T$����_�̢|�E�����������C�+���LᏕ.,E�8��	�\���Z�ܘD�dnNc���� ��=U��̝��m��iCr�Vo����M���ˆ� !ό��
@G�]���:�U�㮯c�7}�d���׾C1ȭƼ3��
�E,�����E4�(�l�C���3��[���'�~hحy	��Jd I[��1b�}ԭ���g�cq�6��8���f�EC��z5L�{�*F�������u��=�j8�A� �vJhВ�8��Z�+ e�r`w$!���5fC��������ܠ��e��9�Y+�3PVƜn�V����s�'���]����;���WYqGX^�r�Y�ǅ��)��
շ�i_͏�^/�.�s��
Wo��C.~���4�!;ZlL����3M�Y\5\���h,�p��3�����
���Q)@�%-���l�������`�s+zI��6� t�Zs��x�/A�*� �[�a0���C�:肹t�����(2��" ��%'!�KW<�h�B4]�
C�#�D�������3���B��X�u�m,�J���;ah����;j��R��Ȃ�m�D�6��k���d}��r����L��G���?�Z֞s��؎7��G�	&�#�5���P ���~��BD���3�C�����]#�,B}�YudjKF��j��6!��m0���f6D�7Yaڶ��ϖ�-�Y>&�(�,uH�sd�9�Z���p+����nd	�o=~t�#�\�Ī=J��FQ,��P��o��n9��!7�YN ��H��>��l!EQ�kg���",� TrϿa����߶�'w�xngTqɓ��d��A%� ��C"s�a�J���ݠo�E��c�Ԡشf���C�QQ�fGW��5/�r3r9L����	/���^��$d̀����f����5[���9��NP(נ�u��/ad�ZjI͍��	��Nh�Lbi����E����Ĭf�i��ޅ�6�H�B��wd�8���!���ž˾CX�o#�J\aOf���N��Lߗ48�e*o�H�3��k��zA�"�;	���o0k������Z���[�i{�x˻ï�֓�k��[5�/2��#靻6�t�uN��	��ݍ&��<~|3B�)�D���A���
�H���}�E���a��Jy��}�x%#��
b����ou��az�65�A�!غW��-��YՌ3����}��wm62��vrh�'F�ĸ���~Q���9��g��n_r2�pH�!u��x	�n��{��{�NfV-�}���DX��"�hbk([��ľ�POK�o!O��I x}�>����W�+��#3~��v�}
mү,�I�P��FmW��4������f��[ig�����Qz��m�Y]ת�Ɂ�굝��64tTf-�k��x"�~����.W֝w�k[�J���,�MӍ��[̴����Q��&#[��N��k���ٮUQC)V���-Lލ�59C�<�x,�b����!*��Fd�!D0f�����,��n�'GLe�CM����q�0��lq��A�P���R/��I�y�G��j�f���X͎�q^�����Ԣ���5+L��FMGd�5���a MY�7��0��|>��W�O��xV��
���`�p�0a 2ąU��i�6��0~E��v�ʨ!G�����zU�O�l�j´f�xNR8J��2$�k�,d$�/�|, �
/��/����Q�R�
�/>��z��PDn�A�|�D:�����l��pa��pgO�F���+^@l˴3�!�%��X��t�-LK��W4�·d�k7O�j��-�]'���K[-���ӲJ5�m��t�+&an��S��~��J�%R�%��R��eAv6��"Ir�c�ha4��]x���4���x���`�^ ��;9�!7-#h/?j�Vu�A�8�M&soVDu�4؎�SZ�)+e�Pj^����t1�m7B$<J�vBܰz $wQt['�Y�1�ؤ�����5��ix1�tj]&�9�V�7ɬ����2Z.�'����'iH��8�@WGe�{TP	4G�����V�zي��C��tNé�ii3�SH#/s�gYHdM�ȅm�K�b(�Ή�>�4*r7�n& �����XMD�ZV![����σ�&�ȥ"�-_��[F��s�_�D�o�K�: <��6�N�.�#���Qa�vYr�i-s3�O6�����Ch�-�}D��k�e�k� �F+N���2J���� ;�p�.��r��`�]h�����z�𶾑�>����{4+�y�Y�g�Q��K�M���(��K���G��*h����%�T�u�N�នR�l��@�D6�p����7+��6�X��ņb�_�x~�wZWpP��y0g�.ږ�X �\3�:���:Ix������r�Q�609a���خ��6AP�)�"���F���2�����>��n]`�����::']�M���Rt�4�L\f�է�oaeEQ� �}����̥$�u*wp\�8\�] �#f��Iڊ���]�+J#��H͸\�"=cyօ���[�U}�puŇ��6S�l����C�u :b?L�y(��������݀�gi���EG^�L7��\�ݨ����tHČ}c��&"K�;w!	�|qG�\b��C�3HS:fl^��ao\#n��Q��0�~��&ܸ��so���1�39K��)2��H��x�]|w�m ʨ}F`��U�w�~��p�ڷ�2<Ƿ-Ƨ��g��,�$��5T@*(R�Ϊ��
C)�Z\��¸Ok\�A�-d���]�~�U=������r�^k��:΍���EM*�bol� �߯>�~?��9(�Pu$	Ǧj`H�@.��G��=�G�C�d��t�<F
�t��)$q>8u�Ba����vr����ޑ2�O��fg܌(��(f������4�BQvD,7Lc\��,��$k�&(b7��:��-��1�,���`}�J{��I�1/���g�((a�C1�HDd�X��pIY��G�`إ��]o�E��ը�`�JWo����E#k*�e/�_S�1����^��ᷴ6��/��^�聆`�$@���/�����t;j@D���뻌�ʑ���nsx����5}ᬭ�=���->��k�9�dfd�ר����
m��y��V��Bч����Y!����D���|	ԙx�KqqW+"�(�v�\b�m�2�W���\��u�����~��zZ�����.2]F��\�7����E�=L�8tG�'��cg���@�L��Ez��3�
���څcZu��sErW]��[��L���.4n���iVn�J��,@�ny=���A�Y��b�:�$@A�y�r�iw�ɳ�Hq���67��8�R}b�"�|0[d�4}��]c��+�~N|�KjAEI���qJ�䖹�p��߽I��as>v����B�$GHP�� �E��A��kA��1��k�o'gH]�����dx�pʌm	�2�݉u��B\6����aÿ�E3.�Ă	�|����M�����H�]��ؗq�Ny��CO�Z��h,�IL���P~ooIE�MʩQ3>�)U�2�ץ�*�MT�K2X����'hz)|����JE�Z�	AZ�X�`�p�2��y����S�c{=id7*��5+�^���{��������uIK���rkJq�7�c��)X}峯k�W������&���M#�&U�3����i� H�ۑ��ǥ�`}��X�	d��>�:���
6�&X̱EicW�!z�Q��CS]�̺��P�R"�������Td!�>ڇqI��TLD��HM�2��L@B�;�S��H<֥Si�S�[m�xb���j�.�������C@y�G͸Lr�k�J9@��B�N���q�bq0
M��NB�ill<}`�x.���������
-���Q^m_��?��4.1aDb�]���5��!�-o���x�@���֦�>�qq (nߠ�Z4�7I�{��蝄�������JM��
v+���C)4��km4Y��3! =��j���69��Z�۵P��%;Y��d�N2]^�`Ѳ�>��㟍���X�2�?�t�4
��Z���m^�S�T���m�n:#�_��h&-�MZ����:�W�+9��PI��m��ʺeq���@�T�����GG-c��?ڝ80u���Za?Uk[��+d�{v����/� �' Q,o�6O_��K��uy xw!cs�9�)1�q�2cS�a��ā�QR0̽��O3�D��� \��I^|Vh�F�~���+�L��".Qhǌr��-xozm�X-V�v�?���%!/SU�1��4�j-��z�Ԟ���
zl9�UMũg?>�Λ2�%�贬�W/qy9q��<�,��4�y��Kg�j9�M<���Ħ@8F^����2Dk�f�l+U�^�b?N�������6#ǔ�FG݈q%�ua�i���t�+a�oo|���0��ڣ��X5[�F�Q�S
����^����MYNXʮa��<v�E9���]`x��$z�p������\,�ݡu��{>��T��{�w�Q��v���X~�_��t��:�sy�jyt?"I������G��20�kkN���p��݃�0 :���!�u����hR�%���Ͻ*����uͼ ^����5�Y��J�frRo�����*MѤ�KҶ1���%�/�"fkk1��������E߲��9])qR1���oUzQ����}T�f+1��Lp��m<�7�e�G�c�K6 }nd�(���<ރյ�AgZY�_�U�K�u֐��,2���d��6q�r�xJ}�y*OCq�B����}
�3�׻�%~|u�6��Y��e�:�&~�e���:۫jI��c��R?_p���Aa],I�1�B
J����q_�p8s[��d#��(Z|f9Tn!��R�"}s#�6=(�=b^_4�?0F�8�7����c��D�oɞ�2��{�	�+6�Vq|�D��aZc�=��l�G����e�헏苼���r�]�D?�D;6�!��^�����8e���FN��1д�H��<]qt�޼�g�d�hts5,v���k�^�U�)�f
Qu����h�AklF'Z�ټ�R|A(����:���fp�%mM+����G8�,�OF��^W]�Y	 50 1{�&˼ALESY�7�d�����{w���L��^V��}O˧n�Y�s�Ы"o� ʤ	�8�����-�~=&��FT�>(��YdX9�(c:e�N⃮
���|��^2���3�;�oW4x�3(���5� kF�%�Z��옇�Yq�$�����N97W�_`2���U���o�a�����tu(��~p���2Ǐ�דA,Z��%���u
me����[������a�����u�Ф���5k��{�p����$M�;¾R�	��=!�L���<Jh��o���o�=��٬~��tnɪ5Ѷ�u����q ��_� s62i���$�)�g'�A{R���H�#��4�	�^�fB��&�1v�@���ws(�|�׹�j��5���ۻ��)�M 3�ߐ���/�� ��Dq����kz��U�j</k1Bb�N����9�gb��6.�^��i�tn �ӗz$�r�-R����+�,*��%x�wy�����F�����<a�>�jw�aFg���~�"�
�y��x�����X����	G~���q�V} '�^���!��5!��b^e{~vA�����ր�n�V8�qg��,�@����j��f��Lg]XD������fC�[�q\B~�b=X2 Β�e��I�'�B�Ё��R���r�
N�eUi�6�֥0~����%�I�L�-N`>k�{d��c����uz$�ݖ��a&�G�V=K�i��-^>,��y�(ʔ����v��ա�+��а�:�L�[���a�����-f�8�dè�O����̬;F%��$S�l����M�Y��� ����� XD��ܡ�S\��gJ��w�G>�(�/�h��&m��U��U�����K%dW��@X&4�bP�.��ޯJ��Qd)v�ñ"��)������d.L;uF�x�B�S���v9%㏑�둁��ʷ� ���&�%1����E����_��^��<�X����)o��$��­��⬙���u�a���,#�,�&O�����N��h��)�o7��P3ib8 ��鱱�v'YHBv�GFr+9� |��#�����CUZ�V۾kGf����t����|�
\�*�9�/���J�Ѥ�D
�������~�!�z�x�er�)j֗�cn�7$4��U�ԗl��3���c0�[#L�mȇ
bE�d��r_j%a�e��#Ar^�Jp�.���wߗ��[i�+uW��_�o�Ϙދ�%"�����K����7�G��oŀ��!��:�C��E�~���M&���$L��T-�c�I�,�3-d��7,mJ>�-7�-���Qr��w1�B��yvOs?N�bx5�\d�!
�e-��*x��i��)R�8�-f�Eo�S[�m�:G�C-|Sv,�����j"F�RL�<쮼�%��<8�l��0��o�-���<�N��	 b��z3@�=K�����m]���	/����Ϥ�jd/����0p�u}}^=�h,�����2Mݚ�`v�Z_YҒx�I�e-���)zef�1lCW&�Lv}��4��Y@>6̋�fT�M�o���j�ad�@dt8q��K<�
����(��T�_FiB�P[�ѐHO�6��؃�Eِ6�s]���)���l��yݬ1����#�V�����Ş�5�*��*������x�Y�h�ϼUmt�?.ܩ\��>j�;&�QX�+�x�T~�߹�e ����YD�����H"T�/"[�X�Kߩm�S6/a0gz�E�Gm�C��tF^L���G5��ĵ�i�ُ�=8�l�ћb����RR�ȧ#���	Aj^�h�(E��ߪ%���{�H�qrvg |sDM�ֽ�b>�Go��݈�b$=��h�lZ[Wl/�ys��")~��#j�]��SZb�9��Z-~y�ES�$���CM�k�4��\�6T�H3�9�A����k�n��>� i=��l��,��ʕ@�F�kС���ެ�0���tb��}�n�����囨U���Q5���j��[��g�؍�6D5Ct���9��A�&�#�(�Q�{]��:J�G�3�\�=d���`qrkƹ���+�x�������.�k}!���:�!KK�l�h1��Y��ށ��LROy]h�A|�ݥI_�n3��fjz;Q�R?�Ghk�5�P%*+șvQ�S	qډ��`�zJ�qށ��Y3�O�=�H��^����9n2ѕ����W�|)���n�ҷaR��fz[Ik~��^���0�X��P�|/,���i[u
�� �Ոቁ����NM'$�L���P��h.���熭��6���X,��a���zĹG'��/9���Tt��^=2�R8��P���z��St
Na�8^��x��\�� y�Œ�6�57K�{�P> B~D�	g�~�H/���<"�O�z���SJL�UmN�uH!��Gٺ2��x	��H�k�#�[K�s��!�)��{쥃F�d�t�X�6�y�'z��۟�5;�k�(�N�(۶�Uҫ�(9�U��P��)�;�6�
�M,��� I(��	�<�����T�'�@�I��l���]{5Q�go�52��U���k%}����0���=j;2�3�I[_*�?�@G�*��./�αWхX�PL�ʻ^��:G�S%n�JËN*3�Z���r�)`o�oW�LH	'Q���X�	�O��3��OE�<:$�|��V���C��Zr�Z�|
g�G1�J��>f\>!�~�F��v��@��ȸR��X���gN�,,���o��f�DO;�9�?1;{щ(�"�v�cc����P}�����UY��c\�W�`�N�vܩ)4���������<�IOǳ���Z�)���$��-�)%nY�� ~$ּW[��"��;�t>�)�a���J/����m�)�=�Z�.�AN~BF�+�4��H��6��tg�j�q���K��Ű��C)�|�yvA�����ǋ��Q�wqf���`̗R��R^B�(��䮺M&~���1�֞S�F6����/��T��1v�S�; `���2�uorƅ)��t��%��=�����O����,g�&�X@q�A����C�䲺�;��%�OQ��^�fЬ�("}�o�W��m�yD�������U�ծ���572�/0�V�f>�T_�ܿ"��.[pE��R�Ǡ{�N_� ��U@��r� j<�չٝ��U�β#���*��Uܰ?#�g��;Ŀ,�@�.��`O�e����k�A��ɜ}'��1��՚Խ���$��c��.;a�}������﨟��>>8z��:@��v=���1a�CB�������Eu�BiK�鱉{�	���\h�l���|�5�uţ��i��ĭ�5�S��n;>��h����g��Ѝ7|{�F���TN�#��9����{>2	�o�V�u�f?ޣYZ9�o,�@������H�9�Bj�@�ˤg����,�ӱ��No�>$��6U�Q�C�I��L�O��1�B<���?OL<.6�%�/؅��8�֯�� �CÔ޼�fkq�cTଧǺ5x�,1ݒ��vl9���M�,�ø2+̋b.�:�ݟ�Vv!�Ǵ�� 2'��o���͋D�.�[r��O7dv�����W��-�ԙB�	���O�m��j���}H?mh?�_��>��58[V$t'XH�q��zt˾��.
R���o~�'�ejzV��<_mR�?���y�8@r,��UF�G������G�7�^�g-h~�36-e��tE���ܺIcMݻ�4tW��������R�0s����ʹ!N��E6c�@�#��C�\V��^!�bp�Д7"���H�<�~�#�����)�*{3=5x;���QA�0��w����9�s��s2NNQ�гU�����#G�_�?6,�g"���=���n����E��>�:��S[N�����0��h3������'ۻk�9z�1ʡ�1�%���I�ѝ9����Ϗ�N�*a���n�f�u~�4S��>��#��섔P=ʫ��rSٹ�I��8�n��A����f行Ǥ��5�c4�����7�9���+��a� Q, 5d�|B72�~���!x%Pl=e������G�C���r���eGl��� )�����[���oʵ�,���!
�489پ����{����a��w��P��?YU�6v���B1�.��d���(�}f�s����is�%Z�0�Oo�۩,@���޿l�w�\U�,S���[�P����h��9�Ao����iK��ƻ"�Z�F�qc��b�6�yxc �l�е}�ؚS��}���#9py�.#���_�'�kT������rX�L#�I�i�H��uH�K~��U��B��M�&�n��� ����r��l;���'�Rv�;�e�VM��ˏt[W�&1�v�Vk�y��wi��M�iP��A���C�G���eeB��h�F#����;!~u� ��-��U
ᝪOQ!�E_�=��?�~*�-J��W:���nE.��<��h�T[�(f�*����}�>��HR��]�ԭ�J�w�ŗ}�$n`��U��l��qL�3���"��
����^Q�x�ёJ�葸{W���~씝qŭ���J�0���]y
�gB�ѡ�F�֪b�a���k�}:I@�ԺDJ�����*�?jw/I!���a�_&�l�pQ��d4$on�(��<��W 6ϯq�����iJ
S�����Aw�:��	�?ږ�YAF���j"��+SDE�:c�36I������ ���0�<h9q�m�58P�wa�Dzk�]LA�����.o�W�f{��<���w�Ugu{'�A=�wH��<h�����������nu�=��I�nU(تmx��e�{C,�/ħ�.B"����[������$�V׮�(I��*`�)d��SP��pRo�`��?�����y|�I�P�4���,��0�Ak��WB�u�<�� ;�&9wGi)�-��F�ݨ�����Ǫ��t���~�A�{v�}�.�jb�"�n�$Q�XBF��n�L'��c�U�V���e�Pr�B{��o���4�����6�.��8���çm�ֱe�òѤ0W�Y1Z���)����U[%�^��r���Á �L=��Uݨ�Ƕ���n�(̃Sq^��������@�
���a� �o��[y�	��)"hŲ�e� ��*?��&�ee�i�a�L��}е(vp��f��:z��m��`x�n��
4+�����^GF��A+ޢ����������Z$m���+t�̣%�'L��J?�|��<Ylp�A�)s�{����>������q��6���^�"�(�vr`�<m����l���*��j�2��<��#�+X1�_�;��ˏ-@/�0U�����MP<c��7.����� ��ɞ��3[ٹ�؞�]O�j�b�b��SC\���ē#:r���}ts�iK�l���w�����+ސ�4#��Ȃ�D�͵�������F�#o'+���z���v�J�����,�����l���#�������Dݶ�Q�Q�"�����G�R���?�(%��֕��_s5�M�=���ߕǦ�n���o�Ex����aJ��2�(�ӏq��ƕ0G˓�D�ܚG.�����"�ɂ���+��xS���Xc�j��#98P�)&w�)4��X��oܾU���󛒤Em.]_�K�\��ҡ��a��,���i�7�e�0T�d�@�pY�.��\0�^vW=�^��dp}�sj���_�^�6О�yO)�de�F���%���/#�o��M_߲T��T#���jӲ�K������zzF�hܓ�/g�|=�(Xس8�ء�vUFBZP�|��R�jip$���Y2ǉ����Tss�Ž�?��� }��g��bm$�t�Z&ϤY2��Լ+v�Ԓli�x��'K�f,�^U!	'x#���#� �6����W%VWzʦ;Y��\ �yBm#�?m�«f���tkf���DV��)5��-�	� <�t\���n���@Ĩ�I��m;�t1����w��&I(`���76���i�G;����\�Rn���c.(B��LC�!�}�Ov��
UF@���)�1��	�(k�l;�8��Th��?���|�V������wR;d�:v���!GIxţ~� n�8L�n���j��q��/gBr1,@��մ�g��qr(�p<�8S�G���3"(���!b��[5�f��5vn#��+�[u�3��t�^�>�#p��G b�����g}�9І��nD�6��<y.�u�ρ��~2�5I�>��"�Gz�R��й�i\^�iL��_�+k�O��.%J�c����_V｟���6�_�H��	��A��;R�U_��s�S�B�5���z�T� !S�����~�L�Ĳ�Y�Cm���&r��p8u�JM7w�6s�!N�:�8����9s�F��|��� ㄁���:!�*�j~�����و��9��A������C瀏�ɼ+�pX}~���+"86z�1j�7a��򵰇ٷL-�A�)��kݵ+u�HD�����;��f)6֧����#��1��c�hX�B���6} 4b]�D��ǂ-�	��p	 +GE���ݯ^�"D�!#�^"ǋ?�w��i*v6���EM��o{X�r�d�Af�4��=թi�au�H�|H���ɵWȻ����n4$d���V|8byS���z���� _sU�\�NX�r��7q�r���s4���h�Py9��)��52��9��ٸ��atH�"�2l�_c7kt6��T�a`��w�'���k��o���?J�SC]�k�K��EMGT�'�D�l�-4�Ɣ	ޢP�.)��j���[X���!�����@9�:Gـ����)L)a��.���-����m,���[��R'�٥w2[76����\�~�5�@kO�e��}fˍAН
߇���Xq��=o00�H��FGc�r=g���U��G� p޼��<џ���Ա�SE����N���l�nEP��J�����!NZl�AΑctp�%(�)#覨[���Vy�qVlG54�~()P���U�|�m<��(]���h7
?gRK{�� Vl�s�ﱸrSٷ��l�K���Lv��a��ޡ�@G_������ű� �Zri�u��h	Z7ԁ3K|H�6�[���9K{�C�ں�O\��F[꧟�HPq�����]}߯��\��%�W�
�Id?�nl!��3��	A�����q�*�[�v3�r���ӪH�l2�f������Avl۰�w5ȏie²������/�f!���Mjt����	�	�j7I2���Ga�|H�m\�hjHzٜ�f/apt�`a-T�Al��Jk����}	$6�f�$1?Zpn!�L�Vf[l�S%Ŭ��)���ۜtt� �[��@X�&E��A���th�(:�eu��U5mo����P;V�ާ��`r�ez]�>�(C�C5�ޝ�W|��sc����P�a�&~�{�~�ϲ����d롁��O���<���e8,�4[�%mT����e�2q}������i��w��^�-.�hM*�/�F:����z�D	���Ӗ�l]�a�ȂQ9H5
���X��t�tre��<sNC�h��-H���K�n�����wn�ܫ,�B<�r��@H�%��L���x�C!�A�:}z�Y���6Y2m�����˞�8rPօ��;9����.'���q?J�'[Au.3����<ǫ��xϲ���ouz���������kU�%Ӟ����R6h��eZ�.|��;�X$6�x�q�R�������� W_�&bJ>��ÁA�N嵹.�k�S��j0�n��$�������w��  N�]�`�q֙:���òhې��Pi�z*������LfjI�����M���⑋�',V
Wt=��W��ǧ����Z#�'�4Q����	�nF�v��B0������ �S��G��,S�=}x�Why��+Ј"���=
�O	z4�������:�.�)5�I鋸&qc;ȹ���;J���.�l�B�Uc�d7�_� �5�O3�xGH��y29�W^d-���WB�����X��*�� )�xE���{�/��ܞC9i,!:d`���jR��ZU�Q��FY��ԇ$^x9�b�/�)���E��q�6>��S�I���.;�.FI�?�����g��.\rhY��2��n,������Ԍ�O<��ٗ�����S�lq���T�ͷP;�x��J|��2z��J�y�>���|fs�~�Y���|C
�"֔d!��e �c��M�y�C8��׫����RJ��b�U&�۟�r�BmDK���(E�g\JjJ6u]��&g4N ��0;�c�61R١�/}��O�IM��J��J��wF���X�3H0Y+�,�fÊ!�ʸ	, �j�Ih��G�j�l�rJ)H����v���:d���ūO�CȦۼ�?g����Z5R��qR���F�'׌c��ΏG����Y�ۣ�����ڨ��ݠ�f��`U)��2�G�*��*��&3&���t��&�v��Nl�6E!R���sl�w��W� ���@A҉n.�Y�i�hg��Ra[���^��A>9_}��[����I~���x�Kښ_��>��|\E@Q�����
M^�9��wv����_�7*�����7�HYz��A�/*��͂�E�e�ו�����ۇ@?@�,�{��f�ɘ�/�:����;�ߜ����ݷ2��_f�4��2��ahO���5��y�q��,�-�5B	/2��z��`ZfՃgr��XLX@;��*g fZ�]F�R���D��x����;U�����1�驍�����^��ʖZ60�����2�@|E���yL�)~v���[����1*�$d�Qψݧ�W��U.d��^o@�*��uM�8S�|/���5GK���ΓO���c�WT��$�ge��.�W١?d^�5<�
K�ԁ��n'�J��4cmh�����_�� *Y4��Gyvl�_�Qޒ=�mqgA���{��t�M�����l<�?����.��vG�S.�wD�ss��!��D�R����^\��k�x��`9󞂪�� [5p�);��?xqy#t��x*��">�dVc#��1K�n��ş��
G����aL�=�d�{4Gǋ�S'�҈�B�����3��@�ȓ�@��V��C���hu^��=n& �����uA�;���O^;���Q��M����?֏���z_��4O�=�N��'�uLZ	��?��s�i}/8���n�m��w�wQ����8$�v[�UA� �;��IX5�� "�0,l.L�~�c�-�w�d0����~���q^�����eʌ�.�/����_�j�r�xIylfE'ʏ�ƚ�=�}��2o���b� ���GY�-,���v.E̱�{>�z�khq1*� �v*�6������xأ
z���8�I��vx�l�r<0ؕT����m4I�1��/��^= E������g���F��%����A�41�$�4�������{)��|������3 _��2���u���q�xǄ��+5���R�9�֔������@exThY�{������3YD̳>�	�c��UoI�i7BHR���{oP;�p�xC�4(�aM��#�i9(�gD��G!�ay`��#?Ń�nBUH���n�<�&sİ�wb�d��;'i��:[EE6%}��6�QtiF���U��q����J��ӝ��s1F�L�����k��)���؏w��1��$�1F�����坯]nP
	��?��K��U�^��Gq��.��ޤ�UC����*�qXm��%��sݓ^pL�_P�I���Ķ�x$�dS%?��y4n�9�h�1lɞ��{7ݯA>��h�I����U�l�A�2Ԛ���8/|AOr�vAi��!ܱ�C��F�� @T�Iͭm�)a@�N"�*�V�����$�S�#�	nK���ԇz���َc��=�p�Y�Zڒ.k�rO���!��"[<�V[� d��~�\��l2�m�h�ٛ=<R��FuK<�@P5�|����}����GA��$,y3�ra�(8�~�#�0C�5)i���v̒n�[�(ѓ|�T:7oA��M�e���U>X���w_����:~:�;1zР��¼�F�S��&��=�1U'#��F�I��}�>�;��[�Ys���_ ,���h�e��
�]���t+]^<F�����_���n��L�U�P�)]i�&d�3��	jc�%"��\-.�Q���x�	_c��Q��r6��Y�9������F�_���$�i�ʀC�g�=��?eR�ݕ��1�"'�O��/��,\6ᎋ@�j�۵/>q��n�>��/X��!��H҅LM�7�$r����'�is�B1?lb)l>Y����FG�e�h�K�!�UC6� ���O��6�=���<��A7�D{˸.��S[*@�cj�EBt��&֩1����l�JO�I}a
v�ܨS��Y�h&#T+��o�����{�D�|8�I\�t�����V�2��cK����އW���~[�fյ��S鹹��re��d�`�zz!�N��� �Re5Q���9� ��Pƈ~3���Ʋ��&D������
�g��Vo��5���9���v���"�B��_jۇ2�)��!�4�ғ���]	�Y�>��6�w����CbPaqH|7uu����I�����=�d3�.M�!�@�sv�*�z#lvc8�y/W����quH�J6��k�j�nF�2ie�����7��B�8�bj�uW��P,��D��/���Xc�pBE�z���v��7[<y�:v��oci�s9
��@R����x��B�����2��Mj��cyjx��_���h	S{e��o��h�E�I�'s���U�WNt�ݯ�TN�>Ϝ
��U{�l��8���6�h���g��ND�̊I�$zƬ(8�
K�@�3��Qu�=*^�(�a��^�>�ܫ��r �x�l���;t����ϒ��~���uj���{8���޸��6��L%��nfL![x��(wֻa��l��	
	�A�h#��뒳Ү�]m�.�8�:�N�aS^\�� ��P�RE�<r;��X��BI*��"�']ź�PF���l�{#s+�!{�G�1�V/��T�oq����u)�4���, �#���ª��F��c �_+�:MA�d�u@�u�3O�Ϣ��s@U_;s�����dгb�dh�S ���kV�'�a7�C8��G�В���o
r� ��i�D� KmX�+L��!18k����V�?�.����n�����cO�#��9��bYa9���t_|�QC����P�͒���e�!4��(���<V�,��3� /���?�A�.C����q �(~�X|ӉE뎫�$�:<�I�S�T�q���[|҆�����y��w�>U�����C�a���9���=��'*3r9�=5h�.�\w�tI�6S����1|q.���*H��΅ OC�w�֊q{��`��Z��ʞzKr]���.׾���O���1)��C�Ӊ� #e���K��d4$��'��u�F�$]���y��w'wr"��Q��_���g2t�H���s��YYnx<ߧ�;�+����4o8�A��8�-׵G~)�OD��T�����3�5�8�b��Y(�rH�N���[g����X�P8�(f0�¾i\LѮo2�N�k�fy�Ȏ5	�5���~f��uK.5&�������ZU�e
d��]R�q�XKS�z�V12ڡ����w��\��˓�Z«R:8ٽ��Ǣ��@�7,{F��i��i���:���+��IN?���JrDAJ�3�ʄeR��F������A��8��Z��RJ����y���~ȓ�d�2|����n������\�p�7z�şE���@�vC2�=~��pn����یxħ�۸[˴�z�{|�T/G���Xw���z;T� {���#��������
0v�>"��V�f/=��+0q{q7�/�����_�/��@�l�(ꃧO_Y���Y��Ծ����K�3���/�f)�v��lW�� ��3��b�C�!�Ou#�� �)2m���w!C眘[t�>�I�s�~BL׉(�ZI�ZpV�B�t�̍w��m3��h����o�f�E 	�?8s��Y���}�$���[v@�˫��\�7h	�6U�9�Cq�5���������79�d�^���^C������G��ި+0J��n"���
*���s�ꫪx�!��{�cBb�'�\�ʍ�Jx���hF��\�"lȽ,����� SEK�6��cG(��<$��$��4��58t���1�Ec'�HX��)��lU)�ʅ���O
D�M���蔢��X�^�|���;H3ᗈZ���U4��O�hA���վ�}�܅oJ���Gf��E4 :�aݗ-6;�h�w����V������Փ*�^)��o�w�B�)��탵u��.@.XN�$�5Q'N��-g�e��k����O�i������\L�/�5���p��'�t�}�5�\���.!��d<ló�Z��t=ٸ*%���u���gFG">��/����^���Vܧ6A�uumm�X�� � D$����l��=�Rк.~�G�+�d|ۯ�C�!�+���8��7-��!�v�&�rd���n�����z��hp�z�:�Qj�8NZ��Zu����`��8*0h4��0�*R=�UU�Ľ�?R_&o��ζ@��d{frO�F$ů�q�,rN����U��_[>�o�B9;�>+IT_:i.er��{>��j��emf�� ��r/#�JLF�K��%'���5"��w�6��T�7%WI�Ҹ�.�����"^�]�S>���(��״��< \#"d���m/�:�\f����,�l�Fctp��5��
 ��r��#�� �}���{R�s�#���Z.1�e��Y��������W�e���K:���LV^�0tn42��U�|'E��D�z���O
 �<\������P�&�)!��[ {OܡU��U!@᩺�$䠫]�CL��غ}*�Ϲ5�T�����i{S�x><#�*��׈����D�Ȗ?�!�\[w3J5X�謩�:g�G�WSړ�"�l���� ��&=�۔�{�Z�u�o�9L@��I��f]dT?׼#�·��`�֯C�����0ֲH1�?�|�����9�b(�I^��X��`"�s�<r�w�<wEp&I"�a��1�E�aP"���SmD]�ɶ�iE�����+�k��S�RX�,m�����DN��66�n��?��1:�Ģ�?�GƖ����1�P��9v� �EӬ����@��;�.�t��f�t�r8� lڡ$��� |,����'}�k�1j�m��gP�h �B��w���nvB�f���ȼ@-e�8�)��e��S�-��K�V��Z�`�\:1�e�w�m���uG7bo�v��0D��7}L��a�E�	ݢ��(�DM�\���Vy� �Z��f������=i�`��ʹf��U���r2��C�Z��˗ԫ?��G���>-��Tߓ��h>A����NjNf�m���]�J럾�->�ѯg���aM!4~-�<'K$�y^$��H�F��N�����Ç�25�Y������}*�A����WU�j�L���Y���io�6N�:����7���r��0[R"N�l�^NZ	RE�2����#ǹ�WІ�SŊ
� LB�S����I��g�b:����@jq��	'9I��})N� L�d���a��USY]#IS�۾�����[W���
+yײ��2��Y��Pk�F>�,�Z6kO�\��3CK�[c�ʯ�Bٽ��-���
�ti��b邛�6�����z	G��`Ǚ��v5 =�x\{��\�s�_/�����-.6*-��6��=:f�x� ���;D�����?`϶�iH��WJ"�MSV��ZQ���;|�-d�Jy�e�ȫ�:Y,dWoW�!|c�����|��`��)�j��GA}0H5�yfM�r[}^�D�����$�j(���Vj�W���r�.T���%�7�zx��q�m��� +��ӛa���ǐ��5�_�]�Q�ſ����~ZelVC�Ouw�K	у|� �m�N�\��ħζP��K S�nE�]$q�uy��/�{E��=�;�M�et��
��i$�^�+�Llž��	q��Gv���t��r�N���q�4���L�R��x�R~^|����l�ru,���Q�С���;������X�(�Z��;���+B/�J�{�7{�B�i8̧�s�xSw&nY��V��m5�Dhݴ��*�dW�-�_p농Q�O��b�O汲��'KdY+˛���[w�zh�8ȶ��fb�w[�w�b�.�8iA� 2�ǀ�f�N��Ki]�`iY���s���-m��L�`f���{��K�=b�������o]o�B,|��Xk;�;M�t�5��E_�0�3�P�����%%셾 �R
��(`&;�9?�Ùmoڑ�U�	+��~f� �M��14�+r�e��#+��I�愬��e'���q�.��4{oJ��W�]�޻(��a�I�]��$bT~�q��}�Z��D�^ݕԦ! {�ɞE��,.Vh�v��<Y����`�Ի	���r�wc���!�n�*"��S��k���^K- ���s�5��~�w��1���	��n>6Z��[#�"��n���V�;|�Rt�_2_��Z��[����Q�����n�Ұu�� �4��["�i("����!�D�ዖ\���#������A9@��B�f��}/�0m�W���z[U@����_7O�"�H�1b��y�l�'�.<���� �$�q�U�g��p������v��c �k�#����?�����f�K�m�f��*`�Fl�>9�5���H�N�����1/��ӹ|�*˥y&��@-%T��W�b������ ��m}%�N��wƭ3�A���+���أ�[�8��I@ؓ/~�~�Y��n�*y��{5������~0��؍7{*&`�'��2Ԛz��C ����S;s�c���Փ8�V�w���d�N"ߕ�%�<�y]��X���FJ�Kn�*�1
~zzJ9�x���)cЋ��Wm�Х� ]�x���]� �j���W���j0�+��7�Fm�׮���?��#w�~��ӑ���Vm!�T�4�LV0�ۤt�앯�t���f�M��z
�g�=ܚ�u�hGS�:�o�d��������"��NR��%�4�K��fh�� �o��`�����v��[7_^�0����9����K��"��/���B������$�51鷈��5ĭ����s��&P�MM�<����81��ue
�^��Evi���,q�f� /ro�������(�^8Q6���`4Y���Z�S�5��2@PY�v�8%��ie � I�3�h�qLA�� ��ϞbJ%Z[�~�[�,�կj�ſ�����XW%��_tn,{�t�D�'�fB�x�s,J<~��p%ʃ�/68��ՈԮ���d���|2��&twuֵ>�#���2pިJU���Ɉ��Ƹ�ԤFÀ�[���]�Fn���&�����s:�s��/���I��2O�v�Y]�Q[��������L2��^�a��m�؟����1�a���#�'���1��c!a�ƪו�(���NP�>4�d���v�{��%u^�~s֦0��CZ���{'�/�أH�9�Duc��Y�
� �QQָJ�C�ؕ<��̞�{�d�:�3��6Yjz%\���Q9�^<��W�I嗰�X�飚l��sieV�kZg)���m�{.��=s���<O��IR9d�Ӥ(gY�g�TZ�"���1��S�Xe;�Яlh�RH?����(,�Q���Bo��Ԥ`I�x%�#����U�U�
��	`�9"Bw�cj����&�<'N���8����̪�qy�c@���<Yb�30x�K�Hz�c 6�<zh�s�&9r��k�o���4"{��J�[�ʹC�P��l��L 3��3�vJ=��ww�_1�ɦKі���7j. �}ъ~#��%���c���#ɯ��҇;�40��B���K$D�^q.r�0�6���5N�ԓ���ykԙ"�-��DH�l_�	2om�?�� �{��&�h�a��&�
4O�\LmNJ�Eµ�\˗/�l}��e(�4K����M2"l�D�^L/�[�[@~��5�&{��re��8ꙓC)o�qUu���6�b��m�å)a"�j�'d�x�[�u�n�-� ��5%mj;Hq�r�o,$f��zcKf6��*P�yn��!΋�����Bw���L�0�����Jny��9�×��.�K#��W�2Yk�l�N����S�X�L�TTt+�S��cv��1��5��R�����»�x�M���T����r��(k���㹝S����,\��bcΗ�%����eQ)1ཚHq��1�#�P�ޥ��Q>	e�x�P�ч�[~�t�2K��I$�[đ�2��[�ܡx�/��C'� �@J#��|]6H�A|�m��̎�G#�^R]@�=�_�	�d�(;!�.$֝$�"ui)D?o��X� é=D{���S����d>[y٣�j#6"i�fBUo1�{�p�έ)�YX&��W�|�̵}��8�����ݮ�ط����ۖ?�C������ވ%��8Ό&[�(��蟎���9�������4Q&�k�l  �N���S 1W�M���%�u�J��	�3ә�E��:e`D�o2�yw�b��}'�6�͊�u�ŉ<-j:���l� v��o)|�����?[:���m;£[O�l���X��B��A����VWI������|�4��ǇF�͛�4B�e����R�Uoz�)���Z�Zhe����!��-���tH7!F1�2�o��l��}JtU?�DS\���q�	����&�e�����g�xqf��M����xl��e�D�'i���^)��/d��\���+�!YT�A%���&�I����c�v��/mOStV���9������կ��hg]fl�M�/׌� �|V]C���X���SE�߳e� 9I��U�y��>�Ǩss��|Z��噵3���Tʈ��߿ߣSj��A�B�z5��ؾ�/�~��"F�H}$<�T~Bt��N5���D�����ܟ��h�������8-TQ�ݏ-������7��WL+#�3�fM՚�(���uN�/D�H�loE��-q���?I;X���}����Y�a$�橔��%���3������%��W�w���[� ��V�L�-\�ѧ��]���,~��3T��޶�&�0r!�Qߗ-�<��W�iJ]���ҞG�h�^����EгL�) n3��Ձ-���,�ث9�Z+�S۷k�Q�M*\�5�z��$�yj>_����Y �Y����NT�g��8��}BL'��H���f��MviM��`��,��p7������Y^�ח��� �腽�v,��sYZ�(_����#~���V�aG���m�ʕwǋ'Y�*�U��:VO"�?G�����W>wdȽ����Jl��|&J��pR�X@���x//�>ƷN)�E_�)[���k)����<ȸ���|Nk{C3�����P��M���^yřN�l�V?�m�R��4k�&�����ٙ�q�R�I$9��,�7$��7�9���0�,z4��������7������P�f�����QC�Kgh�d�<)Q$�Hr�u�V"���&1zW�gE��Rtg����
S��aa0�Ԩu�%�KhqY�|�4$y���D� �i���{I�^�^�@[mfXDT��RN���(��[鱂<��KJzI�|��	����f�.<x�ĸ<3F�Ċ�X�N�6<�"L���<�aa�o$�mQI�U�R�21�*�U�Ζn		�Ň9~ɴ\�b�T������|L��@�7zJ���_��ѵ�}3��>{l�E�b$8z6��ܗ�B��Ԅi`p�[x�:��/O�6ƣ����	�&�cMf�eB�Tv����aVU�<ؐ�ʗr��@]�R�Ż�.Aԓ����$���/���s	W4;n�@V,�[�6Pڒ���t]��Ňdi�w̧��J)U���nXt��L��+�/~J!c!�� ����/���P	��Y�JI��#)l��zI�s>syT�̪a!;
U��ӛHj�B�ٷ(�A��.�b�4�� m���Q�������R����[�ow~k����>�W4�?84ʦ�85�FHH�>��S�EM%h����sU��9�M����gU�|[d$w,��V7�G��b(r��׆�}�T�rU\b�.�[��}��>ّA�/J��Qʸө���Z=�������"pO�jf46�E,W'�|e�����)�F`r�`#�^����3�|�E�B�}��]�Q���G͘g�~�o��h��0�'���x�((��eda3��D� ��(2v�o]��T�9 .�H�V����Ej��g�4��l!�;:P�3;������S�F4g��r��O����l�����ŻJ�󳃵�����f)��#{�?�����w��������
?G�۪�#��NZ�`-`��c�\�"L	����R]O@���6���,wL��,����FO��CO|�2����*
g�@����� 1�,�Hh��C,��!&�m͠�iR�]�C��l��.�7}JSU�8v��������&.�8�h=llB*�od�c��Y]���;��mwo>!��^�B�\�.TJ�5����I��s�/�y3�}�o�T�3єQU��5Tc�G)��K�^��s�H��C�Wd�?g�
x�v}8�G�������5����|p�`���.,���79��r���-W<F�HƝ��O�y�����8<�Kk��&��?�!у%1�z<x��eA�S��WXԸ�vo�0��3>+��d�h�(�Ŏ�)/f8�J8���"cҁ
{+�
%Y�`䤁�v�$���/s)xF�xՇ�K��p8�s/��{=g{!�4�Mx��+g�.۴h�h�̩J���S�m��Y��N�a=`t-dk���ܠ���'�>�t�����g��9jmmpɨ�_@�Ķq�
cH�}w؆����톉�S�ZdFh��7�ӡ+�:�F����z��rIiwIΑJ<'���l!�eS4f���\H1#pp+pXS���I?�%�3{C�q��foq�~qïx>����X^gI����2������!�m3�9��F����"��(Ds|d�c�.eP�2`�?|׍�4���;�Zp�ւ	]��`�g�]�$.ې樳ԆZ�l�_JA�p�ٞfz�ƿO��Ha-�~�����sQ�C�ms�/��.j����c�=I�[0O!���o�-th+��+�@�<Y�/�����;:h(�|��Y�!D�{��ؓ���%�Fǳ��=>�v
.^瑎��'ߝ����&�6����0!M\�f��3yڹ�o���F؂���MJ��4�|{��<:> �8<�M�V�#��=�����HiOW��t>wN�zr�h��,�ȵEO�@?Z�:f�~�^{/)�Ӥ����/Qy�b5q�K��V"s����tnf�uM1���h���K�����\�U��-��x=m�d�����"�D�Ĥ�e���d�at�*Y3���z��6ǡ{��׍�(�Z�/xE0<�\�r��՛/��c�#|���AltCc�w����ȄQT�ƺ|<̨_��J�y d�K�CE'�3�CÔgH��?U��pi�fK�޲W"��}��Cc�lM���2��fO'.�<�~��^ism»� �L*�s�2Q��u�0sgp��;t��(�Pr��ӻO+dJ~���ꁌ!�!k59�qv����)��e��}LTvEp�{�z���G���%��2q0��M2p}�����^�3fs�Z�2��19>�lb �hE���1�z�,_�yt:�lt��DL��[�C�*ʁ�|}�M��,y����=�)-�gD�J�7�j���0Bᓶ�Y�A�<؃,w�l�t�t�2�������P]��7�����]����;�n��7��;奁(n7�����߃��o�x���Or&O�4���ś�bǋʝ��a�pTi]�#{)�͟w�
g�����5��c8�.�T��V�����p+t���{���d8�@+�I�S	dV*nHtS�i�hOr�O�P
k.E����f�=��J��ͥl��Z�ũ#��s���ſ�G"��,b� ��AW@B��B��x�����]{aW���(�Y^K��'�$���|B�m�[ke�,�~�5Y�U����u8�߸\��#u�a�h�%-��N�ǧu)�0҅W�{�,@A${���ٴb	���T�b^�Y�k��������x�H~>��&@�����.2=����/��<6�/���_���x��ҧ�D�ƽ�9$��ƨdG�UQ�=Ԛ�Z��W�6�i�M"��ǻP��Җ���w4�n@Q�'M�� :ܑC�����1O��@�p�ڰ�\�d֗���ԛ����F/��=�+_/nBDO*e�6ྋ&�A�[���;Y/�{�r�Dݎ�Н%T�Z�~��(�^F�y^F�]�h��cG��C�i�:s45����|}@ũu��%wx���{qx{�0R.��A\\C��M�YVdW��#ƾ�K�%�V��K�F���{�Vv��a����� qQ�������Dʄ`6�3�-3쵢;r؄>c���9m���� A^�����&��y�Q���G��K7�e������qv�݌T�������v�h���<^#D$/#��Fw�`畺�So�8��!���7� 2��"I"�:�;^��"��,��N��o�2Ҧ�ĸ¹O7x��i]�#G��R��;Y�.�P�(��gÀO
�6~���Ɩ�F��B������L$hT;��X�P���ؑ4 8p(��1�c�/?�)��ʵ��K"�� F,�U.����r�Kp�Zl�`0�$|����fX�$�;�`�<?'��$W���i죐x����٤�o��B�Z;��k�(�Q�?N���cU���h)�1��r>I��A���{5���=�g�V-��w�B�T0 ����k�}}���1wP�4m��	����2��U +�|
��w� W�͇u4$�WM$эI�,X'�l�����X��fbA8��g�&���c�-b���J&�O�@�mli���3-3 ����e^�I�8޿3����f絪��c�!#^�wR�0!�l�j��B�t�󆡷��[��zp����/Q3���!�/��"I��Z�{H<�S�^Ln��e4�}bc���{�ߗ��c��V���x[�،� q̦��B�>կ2u6z�)�̜���`l|	��(*��?�{�~!;��H�.�Ʃf�ł��_2���Ȟl�n�G��3c6ylZZ��'J���Z?��d��d9�9P-0}�L��<:!��5-���蔦=�C�	�8?C8��`9r�6��ga1�� FYA �-�	���8�ѽa���cZ������ԩv}�9�j@~z���G�;���[�kPF���	S�D�Y\���=����x�р5�� z^�W^5�K�z ڡ㸗/�c,��!a�VU-�#/�W��^�͟T������1�]�h"0��+� ��W��K�X����$V�sY�׳�l��ѧ��W�'�R�o��gߦ�	LYJ@��$�ÒW�9�1qƬ�M��X�ƽ+�}�?Ҋ�`Y�o��j�Ï)BҞ{>_Q�o�V����5���3�!|ɠ�e�dՁ��\,���r��Q#�O���M�ƘZ�6�ϕg��=���P[~�r�p��&e񰾒�9u����~�a�V6<Qr�ZEܱ�������r��Ȝk�&Z�oR|N��`>0�,%��+��f��Ǩ�l�X�C7o(�,�0B#��Ǆ�F�q}�U����B]�>����P��"����o�-�<���jF"���D�u:5�U|�����G3j��
��WO�_����H��6]XM�?��[�[�V�]�����7۩�?
7H��D7a�P�f�/_���]�G%�8*��hU淎˗0�x���A��S�(��S���ԣ�c�+�$���G� �CN�xW�� �_n���\���:LJ��4f�/�
 � ".z6x��~x��_M��s�m�v tvB���bg�<1|U���>�R��pG��f����էa��%2
�
�J��b��=�Dԧ���dh^�������[�a�Z;Aj��\�F�=��� ��p\����N���4�m�:�1]����PK1k�%	P�i�Z�� ���[��Q+)m��\��g�m�;D�&Ķ?j Έ�Z��SWy*h�~K����9���2��:#�q�Y:��M�Z�	�{5��f"��]%�~��P?�2'��ϫ+��[L���=��T�
gQ�=a;�-Yz�����_ �G-�#�Oip#s	 '���b e�a;���=ht��I��h4���u��\p��b%aҌD~G��

�*�ʄ�QE�^l�ׄ���lE�,թ,Bx����ݪ{�Ȅ��wj�L�a��*���o�ݛ��ZN�3O�(�����J+C�	�c)�p{#�ٖ���n0K���w�6/Bs�nDD���e`�����$a���ozL�]��@�ѷ����y��������5��7>�Qk�B[G|�E*<�8�1��=�����*N8���[I��\Ԝu���HV!�:S�[m���9��V9}��G��[6!�d^n��y�4�R�H�TmO?P��x���g�eY�r�8���%H_�hi+���s�:%j -k*��L즫�x��և����)^ݾ�WJU��ƪ=� �zB܈J''hjj��O���0�m���U�~}�����_ش�:P��n*��^'&���1�!~�{/ۘ�"m
g�U�6|�m����¹�l��)�F�*�9������^���4u�V�H�A���씖fb�I��Z,�}�,�F��̙D�*_|��0g�Q���O2s�h�W�q����?Ps�ܾ�����7��� ]��A)ִNz��C>���E����i7J���ZD���N�5f�P�E{w��O&R��Ir���<#�L>��n*$ؘ?��W�!�tv�m]>�$�0O�AZ���@�Ȫނ7�� �ݾ�'FQ�_J:#��@� ���b-,N(�ݾ5��T�d�!��8�P�Qq.8�����v�o. '��Ijڊ<bm��wΚ�� ���{�<�u�ˢ<)�Q�zqxeZ�b�!�8��۰U�S��,���/�|�Dk��j�7K��La�����R��� �ߢ{ߺ�:�F�0��W�c���Л�J�w��Ƙ:��cF��}�r�ӕp�����А|9T�����Q��yҬ��Q7���v�!�z��s���;)���9y}��G:SNǠ"�l�[�B��s�l
�d��	�1i 6�i���D�3k��V�)]���:�տg�0�
"l�FP3|��|ܚ��M���<NP���J>ڤ�>\}8%:��҇��K,���Q��*��C?���~�ȹ�u2#��+W����w �mл�R��?��1�lh�Β�P���Rc����Պ��@�؀��dR�Bx��h��m�@H�k��0�zc�;/�� �Py_"�0�,p�v��ý��翖*P�#����e'��~NPb��vN��?e
������]�i��m[lN/X�dә1��U��}����T,�J���*�؅=�yW�F)��KTw�<�����[$N�����v�����:W���|�o�Y��7�D~}s31�Ե�dT]���j�A�*؁���E�y�4d� Î'��[@"VX�|y�>'����d#�j2��ٞ	��@���=�`M�ح���;��Et[-�\ħDG���.�$K~C���['�0<��ԌOmC���U�c�ʷ��k
��P��:��I��e�������%�]{^�0��teF:����*/�`��~��G���"H���ǈ�7h�$��E��G���2R����J��;� �<@+���
�kU��ȑ^:V�I�<���2`7,(tj�&J;#�/t����N�z溨[�)��)i
:��c���M�ܣ���@�66�B(��l��Z|@Ug/=Xn4�����v�KM��˘��
٧/qwC�ۏR���e��u�����x3[������M�D�M*�Zݥ�*6��7��� ����s&��1&�U����I���|����n������Bgذ/���ob�����T(�B���$K$��#ޯ���+�뫪t,3f�<�=��޷��F�$@t$����0�Sbkւ�����Ѭ�s�TP?����koe��Ɋ�t��K%e��j�*��?4-9Z"R� l5˰�>��8�;��!��/*/�Oc	rr��8���<�\e��ۅl�� >�ɉc9�t�{�������^y��l�H��Aw�a���
$_S��o|��7��x¢�Ϩ3W󐜪�	�(=��*�  ���D��0��[]Y�g���<Qo�a�^K���PĜ@��z[��Q��{����XD�n�G8��؋S�6��أ�ݼ,LD���lzY��b\<�Hr�>!!6wT%���l��U	Bh�	�x1��0f��z����t����'-2�I��@�䮧�Fe��Ha��V�FrJ�m���,V�\�F�<��ChO8��"k�!  \��U��R�Ka�0j\ �bi���n���QT$J�a���HU�=Z�H�V���r ,�ʻ�\����pj'6=��)���WR3����/�-� ���bm��j�DHz���a��k�iƲzx�P����o5�K����AU-oX���u����	�8��/�[����C�5�g�������0���ε�de�</k|rSWE ����� D|�'T���eB|��x�8��:�����<�*�c˰��+��8��/��q����tT��E7����0�rp�nΌ0k��CD:�'��o	�pj�>���R�%q6����}�����ꈂ�jd4љە~�r��1�#���[#��>^�#v�G���9WY
U<��p�?�)�Y�k2n���̥�]��&���<�]��̳ԗXeť����Y
X?�k�������R�#nq��LO�ξ�'-��j�]�H�'J�#P��:JI�2R�0~lǫ�:��n��}R�����.ۃX+ٮ;�.���S.����PY�i䘩:�*u��o�.�o��R���S��$*���>��UI�Mdںp,
}��1��@xc��+���e�7>�^vg�Y��%��&:V�x�&HʥhM�?��c�퓨�sx�A�������mB�O�P�{��EL����"X��u��ű�Z��yd���4y&�s,"�i=J����ɖ��՝4�}�\U�w����rяܪ�KoDa��ǟ�+�(&I("�N��<��ߏ�}�үj"j`ز�vD��Tл�@k�*դ1�1*ҟ���H�!'F�)	|��v�{+��hO�Hg4��(���;��UAĲ�;�/�gL2��:�T[X}$��9D{��J��jfz#K���c�|���h����-�Wd����Z�"��M����c%�*�M:7p�}�	+8�t�S5������'�&�Z�#��':��@�/�誢�Ȩ!��E�O���n�#0�ֱ���ѷYkQ�,eR�/��IǾ��#�dv��*WS��O!�US�g��t����z��K�4[�gix6��Q��e�۳��.	��V�L�/LI/Ng�H���Z��$�]�������״Ϻ�'aW3�u���hX��Gx4�yO��J	�;�tf������ps�!8h,L�V|i�|#�5 sZ�p�2綣߬u��D04#	d��l�p͚�xdW�a����?�	n�pY*`�t7��������J1�<�!�!fg{.�>�|��#ap����؊����:�!�(���=S�'~�(��åaΡ/%[�Pܐ7� T%�q�E �W@�w�I���
o)�t�Vy�V��.�̘�O"�!}_��W{��t�'���;Ù�u�K��H �B-���j"�څ�����sPv��{�����E��O:ᭅn�	Xt�cmoX�jQ��CK��;h95yO�qg����+w��2v�(|�������ߞ�P"Yr��:�Q��O�Z�L~kLQ��n)^*}���=�s��]����lQ$�İY�"�@,ۑ����}�`rĈ��t୆����L^�%��:`'�e������ �ڤ����F����I֚����eY�����1�Â��Ĳ�IC@e����4���� \���
Ku��P~���0��b����F�>/�=D��H"қAx΃�L�^bO�<e��I�l1�5#��'����'�P��j�j�l�}�$����h;W2Zª�?��w#[��/�-�~z��H��Z�����~�]������=�W������5�qk�8����8��6"��hr����^��8�����Q�5�H�JF�������]U��µp�ȫ� ;�PZݼ��VyF;�&O=��3���&��"�/����i;aC��f�+�J��c��5�s�5�q� )����k������g* ��_�,l+�D�E��ز�;"2�2�B��v��Kߢ�Y@��̕�Г�{��\���+A���{��ޡTK�J�/d�
'���!pU/(p����^�R6~���&��5�d���V ��C���!/���S�*�O7�[�΂�t8�P��3g���GE�4h l�%}��Sv�]�F��h�A���;,0;� \+]1
�lv7���+����8��q�Kt��I�|n�{�u�]>c;b�f�:�3��h/�[)U�!R�����;�t�q�7ƿ�\1s���6�,���o��v�1�횲�oݝE'd���G�ӱ�9����b�p͐h����P��Z������$}�d�����+�g�7c��zV�q���V�6�_�� �z	1	�ya��煷�C�G\[� �8��.^�a�w*Q�pF{f6V��D��@�J��i���t�G3� :��Ҵ�%�=�)���j��4������C
 8c�\H���3�<�Oؓ�R�SwrDÔ�S��I��#pA?���?����|�Q8�0h@C����Mue��o|8��L9����HW�	.�Pcݸ���O�����
�Z��a�sv�i�y��3�D��,+S(�G�vQ���g�6��~�ud6�BLa:cS.�i禃�r͟��|�pu9�+g��/m�X�g 焻	 E&:�����������<���0���+��I��6C��4k�I]���P�L޽���#��W�jaS:�Km�yp�Tnetu���Ʀ�t�W�4�*�M1��hNe>�v��ۀp��A,�3:
���i��J�ޒ� !�=
"G��������)�+��J�S�Q��?���V�J���{��ɖ�S���-��YP�h<�Df��zpdʂ)�����y@��=7W����d�,oAeįy!e��;��`�[*ֽ�u|�M�����1���ɭ��L��?\��j�z�ߡMW�:F��9�����n<e���|z��*�þ����9S5n��p��TE��!���0S��I�m�3ͤ���8����H�X�ıZa�é�qb��9 �Bb���C,�����u��E�ˌ��^z��B�I�����ο���	R�Gu��4Ԃ�����<��qrmܨ.m�9פ5;���)CqDd�~ot�Y~&xo@q)��� pb6����j6��4�sf��㚩�Y���	*�|j}]Bh���9�����G41��W�v�8"� <���;l���e�U~@#�1�S�Ӧ�8�m}ˮ:��_x8���͸,��O
��&�]�6��p�fk�g�ւS��xy�ۮC3Y�n�(��9�:6*�A?��%W��A�AJ)�3�k�<���o՘0(�V�-�ǜM��l�<�ʏ'�� -9�b�\˻ݳO���ο�ǭ�;�W�Q~�s�)���qI\{?����~	�� �y�;m��0�y��31���2�c�8f��\</���!��U��)�x�k�\�j���{�,H�ba$����	��h�� ��56hO�$���ҜԐ��ޣ�E� �崵5�{YW���lC`�E� HV�j�����������Q��Hl��1��n�4-��c9��I���m�\�ŮVO���V�o�s�Ws̙33ZBG^��x��K;@�*B�@U�E��;������{�ozh������~�ƕ
�g�:�4�$�?��fp3M�MxC�Q��̀�/��+�Z&dK�F1���c�BCA�7ݫO�w�b���]Ne���A!t��&ޗ��~�V��K��9S�;ϒg#ֹ	�e\v�l����+��up����}�j0n���9�B��-�yZ{�]'�l0|fiR�/��������z���l	�#Y��]fyR��z������9�!�Q��ʣJh�hȾ(K�D�_?���t,b�7[��~��IE�H��Lk�^���u�l��:~<15 ��}����4�� CSV�:����CaO>}>@B���jl�M��<ڳ�)Y[r���L�9v��&���0�+a�c�h���s؅����o�=�k>j4�"�|�u��i�/������"�jw�G,��*O�g�Y�5��j�HȰ���k��Tg����L�������I�a�>N,Q&D���n+;���#�L�Fu'}|6�p"[u�=-� �w�^l����:{�S���.@�2Yeò�
^�d��1�L�����U�}�I���������p����9�=���`�dS	{q�28��Y`�p�*wI�Q�����v�q2_��k�X��i�e)��l�a�{��k{e�2��! S�}�n`,Y5%�%�hGml����vǃ�"E��L����2LCc���Cʅ�})�t� ,{ZS��L'-3��{/ݛ�Y���w��7c$�#���y�fH��W��g(�,����~u���Z,��uq�W�J�p+O��F����s�{8N�w��~
��P��\>vA�[�]�ߗ[
��!�N1��^r�xX���r����j��4v�,��T	����}�3t��o0�ui��\�����y�d���J�sa�ȳ�m!�.U�ם��~�\�)��'ںe55�\>(Kd>��A:C՚���O�M+3qiY
G�Q3A�.+uӝW��
�2�^3���fs�<�(���D��	\`~m��/OJRgS�uw�V������֧/��+`�0������?IAY����s�"�0�oe�S�*�S��B-Z7%fL��?,4\L�"z�
�6x�������D|?%�Wx��f��p�^�A�po�3���0)�w>����W�v}�FX�)>��sN�743�EB~Z��~���4&q�B5�9��,��W"�[�=(��)��0f��f_�z`�o6҃8�x�������=C�Ⱥ�}��w�F��;4��3��r0��&�^�q_��#<V�K^ת��������d�<�S"|���H�}�L|r�D	����|B���!����ȃ����r}� �zm��7vmL�y��9��j�X[=��^ˑ� �� 4�%6��h��S��=i�+F����}�S��R�	8? g} ���a��2��T������.�JM���� ���zV�|SQ�R����>$�H���i%����C.�6�v����S�g�f� ?wx������Pm7� �v`�{Xeo1el4(��5��љip��V��$��y��%�����L�T8�i�����u�!X9{��J����'h�X��g��WW2�A�5P�ײ�U1����� ��l�*t���ڷ%�n��\�zH
�q�/@Ͽ�?�ZW�u&�dE��mټ��yY�6�#��<K_��?�]bC'��A��F���ıo_�`Y���d�Y��O�d	i�3�{&0rw�ޥb��KbQ��XeƂ��ב��09�o�22���[�U5��]	��ns��[:zm�+��@E�7��*���G��.K%����m�ѭ�j�&�P�j�1�Od/P�S#~���zvIj��l�;?#�z�o$ Ꮳ=PԀ�krG�������=GS��y��a�du�g���	DF �����)�;�=��02+!��
d�|��"�-���D?�]�p4���g�h -ᅮ�kp53�ES��+�
�lY���m��e���6��z�)9�c�[�go���}���a[�I�$�`�5'ی<�f#%����u��(CW�5Sk�J���`���#��%l|�����E�ӚdUc`�	Q�
�8mX1�:�j#��%Q�����Р��%�֪�y�p��Y�'�}H�E��7�ei%��<���;NmXa�s9_lb��1�C�ĳʷ�ƽ�%��$�͢�Ƨ�k\=�(Y�@%���B����\W�$Y����M-�A�W�k�M$��%��������{��;�^�0���	nr�Pg�o*��N�v�тc(H=�1-��I� ���z�S@u����(�3�7���fim�0v,�9gF%�?0Ѡl��vJ��~����S@#����x�漙��TZ�[�.I'{�~���2h2�q�3�ޯ\�C�c!����m�N���G�	�����(�����^�!&!����/k���ɲ��. �m���=� /�2��U)�� �!X'���c���Wb�;�������X�ڞb�>��o�r;D�3���*J��4������p���r ���pg�d���<Y��D��PT�h���'�gC�(�YFg<��7���"RE�42:��f�H�F"�|L�����n3��$�"6�N/o�+;++x�����iɭF_��̅`���P~���3n��o����]Mŝn�N�p�5�E�ak��@��>�O�!��+�d��U��q[�U�,�Z��3�2�����NU��`����)����&9%<�t9Z�s�xc7!Rʝ�t��4A�ـ��vV�K-s�X'�"�8��x˫�7A\�ޑ��&w�9��d~K;�0h�?Pr�0��2�����X9v�!GnZ��������P�NU���ėg)0
�Ze}وw���6z~�yo�����5��#�����J����2��qte�
����l4�	˱o ��cۃ׃d���L0iO�#�n2AKȠ����q��hd�C���U!�ۥ@F��B_���w�l���D�B��_x(�5���~dJPI c��D���? �:��E S�I����1c�w~$�G����P	�sw��X�u�[��Xg$���|��w�����+y��-Ŭ����]��	�`4 c�3g$�z%PB�\�z�=߅��ySa�2�拥�5.�����!O15�	�I���N�O�y�]*vgNh��r�f�C*bE�X�0�������������ZM&@?�`���c$J�%�<�h�\�Ȧef�؏w�c��9
k�0���1�9��g�	��0=W�-��{��A�$Ƃ��T���?2�Nk!W�WN��F#�Qa�뼭����/��S�%�K�M��%�_���Ez$�,&���P/(	
&x��Ǩ���Y�MX��n��]=CZ�t��Oz�0�+���	�F�F�'�����"y~�Br�;<˝K���S^�1+�zh�7��P$�>�Ғ�hS��=Q�4>��%�sQh���	x:<�(�^�	������}��(b�B�%3_34jĴ<]?u/{�4aI���u�t g9Խ���\����ZK)y c��F��&���3��S�[psi4�8q��{�k�3�g���2�O��W�¢[��M��h��?�F����vC	�م��hyf���TE�Y7��i�Q��
�	�m�����K�<�z�_4����)20��~%ʤT��AHy��o�n�}�2�.|qZE���8���D��7�≧C�I�����E��HK $̈��dS0�2�ҺL4)��,�_�Bs���D�i���k��i-S�����v���8�b79����ysCCb��RQxͤF
#GH�h^2��)=��o\�r��*!P�����<�GVt�Y�����{J�t�霁H�Ⱥ"7�݅W5�n`NQc�:�+z�h������6
1,����Gn亦� }s� R���%�/��R�>���vUP_�C��"��n�e�FR�M3t���*��j53�km��vC>PKs��a����b�����$	/�]�$%-M9T"_��������V5d�c�KB���,������ec�Ds'B���p����g��Е[O4Q�F_���E~;�܊�ЌQR�ʖebb�ϧ�WG�͝/�"I7g ���p�T>;!�.5��y�%�E�>o��a�S�Ll� ������~W�o<iG	xa�|��f)ؚ��U/����$AE-��Iz�=�rki���z�&s�f[��xf'S쪁���.�����{�(��V~<�N��(Y�kz�O���pqmc-�%��cl�]����b�?�k��KFb�)$��.d��$A<�#1��<�&�J:�.��P�+��HV�vg�ir���yk���`���$���҅0^�C��e�+p�۱�+{4�	8*�-Ov��(T�,m�P�#�&���Ǧ���9�&�r��?ړ�q��ry:H���"z�� ��I�H��0H+;ˆx�;�䞁�����W�X�4�=�b�)�u-G�n����,A�0Lv�14�o鼵��,�� ���n�K�ĝ��X~��l�o�=╻��ϡ����dSt�G7��KF�i��S����I�͝1X�x\��$���FPf�����v��D�/�KD�w�#�7�����!������lr��g�t��M���[%8L��?�q�-i"ל��k6m�j��Vy���T�9q������c�d������
�5�"�+�Ca��+k��1Y]�"�t,m�@��s/��rj>*���-3�d�}���� t�qf���oHC����|&��a7�%��}�8(�Q��\���2�z����idMU�yF��2Do�Mj����rV�-�{��:�^g����P���@7�v6u��:��~�����[OM�=&ä�l��}71�;��S��fN(\=�:�V3�f;�wB��ڌ�9���.o��E�>m5k���gm�*�(X�hHva�*/���h!�Kʱ޺΃���P�b�p�v)y�x�QÈG�Ϻ���WW���g���A��Rx��8X�/�ݾ����b0YjnJ���a���k�?OW����]&}�gi�>�j8�J=��O�Y0������'���z�=1���/�6� �O N���1+AO[β�6�����+��X���-&{8UY�c��3{���G9b/��U-�>H�/���&`�AH�P=�XD��Я���s�켎HJ:��X�2����+ళڝ,��n"A�'��$ǈ�9��x@ݦZ� 	S�[��X��JyU��*t=jt��IfT 8v .�hr$L�����((���Hƍ���~�3�*�����˸Z@���q�3�T$M�}�}��wU�qÌ/!�t���\�Q���?`��%a��e�X�EG�9��0�*78�9,X�SpG���t����Y���Y*���|�B!,���L�� ��p>�1h�6���^��Q�������I�)�V<w�1�~�U͉���Af�����U6�	��>�g1�&�=XP�_���Al"'٘�ݺ
zO0��.`�4t`��"��6��_N�O����Ր��/\�	.u�o`/t�y�����fP���ie�D'pdp\n	v��S�ζ�1��_�,�m4o2;�zE��=|��hjoƣw���G�ֻ�f҃ɿd��*
��o���;5��\���!I�8�:r�2�]�v��H�[��^��:u9�:�!ۙ�0��|S��y!���f��+�ےR��UQU~��� �q4[cD����g���tu#�����O�+4s�r���J٤����5REWJ8��O��N�e�g�d�x��"�I�rͺ7g��}2�)��V��t�G��}d2)&k��驰~}�]%�F�j,���e�'�2��	q>���W_�*'a��(�WV��j.��u���I�"8��<ع�=����v�Z�����gd��*�_�%�7��� �|���;�a+]�x��{�O���MT�B�"S��j. ��/��#���Y(�w/�HGeǣݙ�(?�_-��f�e%r��$�=T|]&�M��_�����3Jh� م�g�UZ<~�UP���+�Ĵ��2Qp������{K�/�8�|��$��k�޽�'3�7�o�Q��;��KXN�S�D�H��)0��:�#�Mu�m��l :pC�D���\�7`jS���:��Z�ʟ`3	|�t���8�8���C�:|��g���nw�).���#jX��v�A����_	 ��p�c�ӄT7�t��n@B8�/���AJ�<?�@qa�QQi]��R,W��Yt+�����.Kqͫ$�	�5�y T<|D�i��.��v$y��P��#	��$�#>��!fy������j���/�ꍧNr49B,���Qa���-o�c:�!��j]�Z't*�;~R�V����`�Ty݊{�ܩ:ZK�<J}S�NO�j�U&*E�����7I�-Ka3�,�>}��	�o{�["�I�0���U���D�RF2�^���J�}#(揠���-Ih��W����M_(',ҭ�nԭ�n�����v�������AeH:J��д�
�XމX�
��������y�m9��;G�G�5A>
f�-Lo�9�-��lb��Y�7eS��V��4�o���Լě-8.B?��i=ϗ�$��]��������i��r2N���Ӗ?�7Ԟ���'�%ǅ/x�|����;��
Fu5��)`xu��Nmj%��ě	�ZZ:X�ۙ�|��yג�S-��Z]J�w5��4ؐ�;��	�	� Ů	��Gp�O�:�2p|�nSy��݇JX<�����4�P� ��&lH
+Ib�Ľ�:�@]�,���ڪ��r!ZN��Ѫ�*���m�W��<��	 @�<�T%��h,�j�>��W|o&[��{�᪳�����j�<̯b]H����]�r�T�K�G53�����CI������!��������_��i��c��������ͫ"��nP����8�U/V�3�'���	3}�����4"���N��LT-lRc��jqy�a{�m��E�~���*��H��A,ST�`���}���k
NZ�0��'cTj����x�{]O�D��3/+�^��Q�[�![���^�c�F��/%.���,����9#������Q����RҸ����(��.I��u�S�4a�78^� iۚYWO~�|�r�|�΍`�����G8Zx�x��bRd���`���30H�N��q+�'b҉�O��E�;1����J��/up��|"O
�r@��	��`ѫ�q�i����=u�H�{�v*����� ��^�����ڄ�X�Z�	I<�N���=�W�5�c"�������%�*��_�b̎�ƃ=�K��L<#�ɖTAF�u�,�"�>2��Y~|�-�i3T� �އ���h������h��	���)��'�#B/]�~��B`{Kh{/�L��	��o��C���!�N�����L"b�fkI�$(d]8_����_��h��6�`�B�=��T�w&�6%�F߸i'6���ğ�A����W�sq;]��c�lП*������=�YΎl�U� �C��ʡ��ݙJ�p�6��ܚ	���ŸA� �|�����̩2:���jt� 
��g�rQ���B	�%�#�L���
�?c+��f�!o[k�}�KJlӹk��.���0���� -���G6����*Bh��>�0�q�2H�;��>e94T�>a�!�������䱜n�4A"|--d���<c[6`T���L�����T��S��\f<@Dp�5��~4�.5r��S�KJ��+��"�"���^��ޠo"�%G�x��祙`1���,����y�P�4�\��|�Ɯ6���B���O ��b_��1`��d����'��{��y&X�]���NZ?�g� KlP~�MнH�l/]����c���|������;D��ˀ�o��{z��*��Y�v4_y��{�ku,º"4D$K�����2�ZQ����;�[$ߍ����������G´��lϊ��C��OO{���=����X��lT�6^UO�rc%�.��w��8�/��g�{6>B����9�|��OorE5��#�� L��+���r�^���N�Kz�z�?[R(АWux$1���d�;��!>��t]�M�����䦐�ꭉ�y�;��A�-�&�)\n�`=�Q�u��A�]��I�@�h��su9���]ͫD,ܑ�JM~�e�f�٨�z��ڱ�#�GE�^A�7+���K��.W���G{���CK����wV�k���M��`�O��O���o�D�'!��Z򉕫���A����S�!�Wq�4A��K���ڭȗ�Z�f�:���;\'u��ϱF�iW��&Ro/�1_N�wx_uJA����%݈��*T)�:���=!!�&a�,d�p0�9��$*Ã��MVxQ�*��7Z��D�V�~���R�9f�a��t���@8��9eNVP�J�jeZ�V�3�f`�2z�飪/]cu���H��+.���"�>W��j�m����x�3W m�'�r��8��GJ��?��2�`y���ڀ+e�s����<B�, ���L�Du����De��y��ͯ��OO5��D�JtaWA�F�9��RF`��܊������c�G�Y���	ȦyL�xZΧ��ߨ�CK���mW�2���h��۪����1���0��� �\d�����'  �{'^�P9�hNp��v|�7��8�h��S:?)�K[2�٠z�����/��]��JA����ZFr��N��b����Q���j+ؙ�v�Pn��]�~�.b3ua���Fpݣ�Ҩ�y�	���I�#X�Prer���ۢ��U@ma�NS2MR��=��>�G�cƠ�~n��=�9#��O��h��Oi]������ĺ��8��u�:���i�hCx,����Z�NMi5���&��u�if�R��\qŹ���>Y�z����yI�{:���@��"t��	��N�/��Z������Ժ���ϊvs	��?���L��le�3�3�*d����%U_nT]u�}p�,7��I���jzP�p"ilJ��Go�k�W��]��ҪE�>9��lt�#���w�����!������l��-W�a���<PWe:_y��������r��fY��G]�~��H���gU`j����]n�2ѵn٥�3F�#�φ����i�ӄ��ܗO6�zK�u��J�G�0~g��Y�m�n��rW�|r�A��A(#����#Tccs̑�x�/��wG�P&�pјLBiJ���)������1�jEg@�vӂ}�/�/��m6�K��y��6�C��jo��F7Bg�?9�%Z���M��^B:�5
E��z�q� 6��ѽE�T�YWiЁ��p�������7��Cj �Kc�;R��|3fH�k.iƏԷu�#|�X+�h�?şr"�ūȥK�V�v���g����9i�r�w�VQ0lN��xͥAߺ��C���hM5m�ك��u
~���X߈�G���E���[r�Ego�O��@����Jy{�Sny`���n�\�,Ѭ�!�$�Lc\�G﫣R��/�`&���U+��TKt&�`�J*��7|Q9ڔ�2b�fm��|X��|���UR�,��0n�j$���$�j���L	tf4���"6�rRa��mI��>8�3������RS�Kɨb!FS!�A|�Ј�#�z0ͯ&g_�e�(�U}if@��D����ߧ�R~]�Weǡ�j������3�ѥ�,��\�������*��/D����C�ɓd�5Жy��H�D�}u=���[�j`y%|Ɩ��"���C�&.�,2�m�������CY5Fu��Z�������d1O�=�!�o#MȺB�.�Tb�U��eU#��:f9=u=�}�
{[5Ų�x3 �W�:m5�%k���_k���-�ji�T�q�qȽ����Z�� =�u���Z�~��I#������ґ�e���-.��B���B���,��������
	����n�c"����Ы/�M-�� �tvBS�IER2�F�6��hi@$=�V7�>:!K����Ь�w]�G�Py�"���I������"��Zs���$�f�[S�*q�Q�Ж������
��Fxu �Q�S��f�/Ί}�����`EH���ʠ倲�(Ws��v~.�gN}�Jv� ����Z�
V��;����]-�-X�*��-���!2� �7,��q��٢R�����y�r��B4`F-����Ϊ=H��9
�.�	��Ū
'Qʕ?�=�A��R\9��'�I�Kax{��0LϠ^֣ٗ\l!�[���W3��c�"R�@���L�r�;����9�/�g�C�9�CcL"��C(l��dg��U�;%R�k����^д�.K�F�ǹ�2�WǺ!�2лn'��Sr�L��Fj�D�Y�}�{����2�f"C�ʺI �S1��Z��V��1��ǈ������M��@ӧ�)��Z����dV ��ⓠ����DX�o�ܴ�̟�ib��W�Q�V ���Ӷ�沤�Ҹ�h��H�����'�����Wi��9�g�"�r�_%�L����F�W�`M4�f��/��q*�Z����1G�7پ\�В�����=Id�
w�62����w`6�^iM0f���X�A4�u�
�.��K1����TU�A7����Vؾ�{���9$���hS I��n6z�� ���O��ws��<�7�3��@�A����+Zڋ�9�j�!b�%�u��.gIh{��TH���a+����p��-p�
��H�~�fi�|z�p1)���&���D��4�[A��|��f!-l�+l^���_lz�>��x�F�Y��7]����7�~��a��?��iq�����Oig	E��:�݋Td%>.�����Q���{�\�b<�+�"���Q@�#h�����C�މe��&M��D�d��U41"Q-�y�8�Q(y�C�3Y�6cƈ�!x��!�Lpm� �n{����׈[ ��V����e�>����_��zĄo%��]�}|��/aX��؞&���N�2�\��������jn��"���z���+U�]a��!a��T��.p����ʓf<�\+:�WT�x��tT,ы88C��xO)q*���E-_8,y�YW!���KOQ�������A7�6v��]Z�k��	�W��'t�ޣ��2��FW�|n�����M<�k-���*�i����a}�H�%�)�(\��2p-�pZ1��x�m-�}���~ ,���b5*.q=^�:-��į%�������4����I�t�R�l%�����XR�?ګ��{9��W܌Lgƥ(;�r='��X[��B�s�����̐���������
v��6`�Q����ӣb�gb�Q�@����.�'��D���0G�Ȏ�GJծ�	�5
����[l ������c�۩���ө��ƻ�>I?I�U����f�'����V�3�����+�Հ���8��.@�l!mq?�ݑ�k14��d��!��"9�t5���1rn4�|��>����6E�����7Ȣ��E�Om}ˉ|{�"*+���|W�p��Ħ���i����y5�ĩ���%�����v1�Z34l8�����C�ݗ�͘.�u���]���w^�$�">*$�-[���#�����h�w-�΂GL��g: ��2~/��,]`U��8\X��J	��p ��6ͷ{�dM�wa�	,A�����Q�w� v7/�Bu��Mk8V^�z�1��wg��ʴ�%�d�x	ح0��{�84t�.s=�%G�+$�a��R���(�9��$zH�#�R��L\��w~}�VbuH���-�s���x�Qc��F��FgSA���I ,8g�Mpx�	���"=aj�.���N;� �<���}!P�h���3�%�Bu�|��U
_�ały^�L���J�`9�`j��>sH�M��5�0Ҹ[3tɃe�R-=N׼����+�J��[�L�wg#t��G�JBԕ�c.we }_&F2�W*�櫣�{�e�|:�xk��WԹ�GS���W�+���u�AۈΪ�����qK�Z�ùN�lX��ǝ�)A�q�ܥL�i�C�V#�ȃ���q��}�8���*r���o��v�\����� �t^�Tfn{���n��Q����F˳�	T��E�`�Q���ũ!S)�U�Vr	�P�\D�zǄ|���C\Q�Pj�~3�O�;�����O.D�?�,�%����/�#�Z��NZ�gu�W�5$0c��T�X�����j�L�u��0���C�˙V)9�)�E���4����b�����u{ս�,���lg^c*�$+UE�"}�DCg�B� �ԫ��8���..T؊*�T������/V�ݐQ�:��/��(�����׶������[�=[���8��Lդ��`�,�ȍ�n��H��;�7<AP�۱�Y\�D}+o��#�;?6� �e��]�jb5խM�n�֪��R��(��q������)�+���F�׊����fC)ф�m+�غ�3������D{(�'���~H��g�XԨv�ի�\R��e�pq���^���NyJ$?�#���xIfBTr��u�k�V�Z�M�_�f`?����\k�}|)9��!����Dǘ�"�hc�>����-cSH���W���H��
rY���׺���A��m= ��YS�\ک�JH	��0�&��!�S��b� i�RY��.�����T��]������Y�VI��d��\?�nG���btV-�Ԃ� �Y�.�Ch2�/��L�[��]���@���۟�S�.�`$9?3�;�A	%�����oMj�mJ�@L�2���s=��QS���Z�툣W�K4��/Gx�da?��w���f�,������IP@���oTS��(�i�G���H�4 2�=���\?~P�;�qxH=��qZ&� ̧i���JRt��s����P��=EM�4��|�e$f*��"�|vX#�*��v~I(�)��~oh���S$%3 ,U|/3��� �d_$x���n��������5��%~��]�����-���S�ʷ��X��.�ǃwJG�]O�o�M:��$!�֤g�c�=��S<u*֏�_�8�}\�;����f�'G�S[򩄹�z�\g!���`��4���tqt��<2[���Ϟ�D4�;4�R0�?f�c+��)>��Q�����$W�o��T˙����]����1�&���M/��@�W5�) m�ױ��`E�Ư�.Po:�͆Z��,�������?�j�v��*)������־��KRV�fV۩�	<��{3��,��32�9�ʂ�wT�|����P-f�R��5!8WWe����ZNy�H�C��@�k8�����{�L���L�A<aN���3�#�}tnNE���6�a}6ΕR�n8 ���-�q{[�щZhծ�v�;I�0O��B2����P��y�}�@�j]x���5�i��ۨ�7Q��e���5�P�<a����Nhb��-�AP�}:�j�@�e rN�Vs�'��V[,R)l�����u��5Y�S��г6���)��~c��:��Cl4� H��������# 4I��]7����:�%g�A��>>cy]?�P�(�>�>��=|E]n���9�p�q��c_��Y�_!v�k��4��lr�(�K=-�'�L�<7��Ŧ��'u�$)�J�3:��lW�����jLo-#]�[b6�\__��)��Cq�Lj�N4��*��s�=ᙇ2�y�о�^�ڌT�V�/��W�ȣ�.����'�!b�#'�)�k�K�N1�e��%����5��I=�����U;n��V��uS8v�_�)�ĭ�.� ��#>��`�d`�O:��'�S����B���kG̣����i�2 Y�q���� ���K��:o���t�^�����­�| ��u�<*'���&m��s����9-�K��Ef���*���L�'�Ɂ����5�7���◳
��k�এRO�!�/� P���%�EX�jr<�z<0]�J��z��^.����3l��3�k)b���hCO��氅D����E�jI��K�%�z�&�f��'�~���p�R�جn�����H��ah����'wj�Ӗ����텦����(�|�(��qTj:f�� �#�S�H�&+�e�j��4"2V��E�b�:�U�3��ܖՂ���헅�q��XV�yI�K�ږ⠨Z�D��覝D�h�Ui'9z�V�#� }�����?�Ǔ��#="3^����J/�$���աɫ��s�:'��J8`��[оRJ����)��m�pYW��3�O���w�����*�"�B��n�&vuf*��^���g��$��7(�T�UZ�F)�:ɻ�|n�$6s �{�̙����s\T�j+����y����� ���yC�r^Z$ݱ]�e����_@HUʢf3#�'�T�M��ㆿуpJ����NP�_-&��x:b��s����ͩ�/��Ṽ�Xꣳ않����h�w�zۆ�2����BV���ET���5�t_�9��x2:f��,�]�6�Ͱj��^��n��V���o�(n�}%����%k3�^� ���{��_}}z��� �8�0�q��K�QN�o�_W�z����j��/�m��g� �3�y���͜:L�g7SB���2x䁋O�h��m���a�*7���9G�DG&�")B-*�w���w��w��^�~�R���5���s2�N1�j�����h��߆�ѵ�iz5_,i~Ѹ$�E�񜔰��>�n:}:@���G��9���f���h9�'!�k�4LԈ���:��v	���4����NPn��^�9�� bx#QiQY,C>�?ư�ͤǯ <d7A�&��!�����i������Fǆa!��|����Ļ�U�+7Ֆ~�>�N�$�S�#ߐo7`G'��F�k1���p�h4��.�R�ᰴ�H#�>����*~�9��Xf�:�s%�$�ye�}Á��Џ�i�<�Ů���AΔ��)X������Pp1Ig�9�q�6h��!!"�7yAb�I���Y6B���a�C�a��RS�X.  �Y�۶����
G��lۧ��h@|�,7�6>Դ���8<��^�nNɋ"o��3p5�A��\��G�'0>uza=�<� ��ջ?���}����P��'p[/}���U�.�
��Z� �R��k=���`t_�5�ǥp��ua�"1���Zij���C���s.L�,��"�T y��|�۠��G�g�y� ��({<��m��-��'��fo�hEWl����+����=���:��Y���*Ŕ'���Ğ?�? ~)�r"G
ð�,�kV���{.��|藳em4�,�2��h��&w����F��7+�W7��s�w�a{�*}���X
+<���5��Sq���!-��r����[�)�����xg���߶��}��lZ�'aWn����.�n���i8}=�r���ෟ����y��o����r����2%bj��D1c�@��^�f��)XB��>F�CE�f^��^*J���Jg{P-!��ZJ4皉�`��֤�;�D�茉��g �'��]����m��N�kLW�YD�\�̩ �‘�GZ0$�a#n�]��G���HY U��&�C���.��>J��FׇR㾚�jP�~�8�����X �U#�d5�*QY��G�ĺ	R�`�xJJ��<���&C�&�̹!z�Yp��� fR>4�8�[��^d� ����s�I���}o��2�t�F���ճ�Y��Ŧ��������.����z���j3�Qo�%��!��S�������~ϖj,pjz_�2OC���nj`OW������O�m�~���|\�&��O���~�5u�I<�(�?k��I�Vy�H�f�L)#-.)�����x�1"��"X�� �O��˝<�ȂZ��{�<�N�(UEP��(s��1�%xF&��ĈHψ��Q�ѓ�-�h9�wr;A]_8�m�hfyG��,Ij���gG^�8�k��i��Z� <V�F�m��";Iί���|��w{�*�,�E㓾�u];#�md`�:T�!Vh>�����2Ok�Ԥ��e؞%��F��*���^9E~����mg�Y����)����E<�D$����k����Zڥ��q���l�｡y�/j�y��e�B��R;7���O����.����a���<Cn�jJZ�o;���8��O+�}q>�Rt���J���A���e7�Ko�tc¥"}̧��}_�������F#�sDSu����������mM�д�?6��ӷΗ��F����X��T���]�����k�c��t�D�uz�X�L(\wOB�
�=������Ŧe��(8�8����.+�`>��6{�.����$��0t��N�Uq#:g���[�b=C�)B�@��B���;X(1]��yO%�
�[hKS,�����s�|����A�����v�:	�͙d�����
����\����3z��[��� �������m5�y��!3.��s�O��ۤ�q����k ��/nң���o��{�r[��k4i]�o�q�����*�0~8�Bu��ǖ2��L���p��1���yx�����o���W�WV6ƅ�&�[���\0���w#:�~IeF�&�<�E���/H�*�/:�/��Y�jE�l���ĉW?ʏ$͜��*�S���+e�����ҋ�!͝��I%n$+֍��L��G�p����:���^���^(���%^��Qp�ϬZy���qm0��Ϗ��N����:A�@w����]����S?N<����}:�Q�+Kz,���!��pEp���ݦ�_�d+9vDs��9��#c>��r��1вA-J��r
���!-·����tT��O=d|fPe��%~ cğ��r��-s.2�]A𤧟���=xwY �&�+ͤ�Ǔ�ɲ�ku�J��M�ąsM��+j�U�A����:A�"�n(W2���N�������SU�@N�U�~z�Ʈ+sS�o�� �F�@�r�U���JN��H��{��׀�巄��]ju�n��2߃q+W\6V3�q�3��U����l����Û0K��/󦞿��无[�_��6���fx�*����$���/̷=��܀��g��F-1[w�D��^!��*��:��g����_#�A���j�7��Vw�ìr���̐���b����)�!A9�	!;��c���%�⽑u�����f�Ô��4�e/�{���|E�2����(�L��� ������'�gK�ڏ,V[��!G��$j�z��ƺ���,��S���o�����]���A��E�J��"OR2���]O�/ڥt��u�r�J�QN3!�/��T������\p��!@�t*Xxq�����8�n�f�ɠt�X�b�sq���o9���-���"8Q	�y(:���a�/���{[&�������]�����ܱ�8B��Z\MKގ�fۧ�r����.��#�K8kxޤlI,4'?��Uq���wf=��^�X�Yq!wو���K�#ݻ%F���K�LĚY	N��T3la��M*��a}`7F4� ����y�5�
OIԢ��c�u:��_YJ�0�S��-��5�ma��A��i����%�纖q��A)���
�0�˃,�s#��(
t+[}L9nѥ6N���ɗ��˳�����ֲJ�W[�.��7��ukd��$K�|�ȱ@&k�e:�R�i&��ƪ�<�}0E�⋢�� �{L������GH�YBY�0-S44�dSfO;YK��v���iv|�<�]� ��-�d��������>�?}�v-�iUb'���F+�d�bT���1�����a6����_-����A a���"�Vْb#��'"ydC$�<��+��-�V���J�O��hxGV�6�ޤ������^�*ѝ?ae����b���9�A��]:w�,2��~;E��-��c�c��Wa}�$��(Y��0�v��bd��d�qdGM�P�����('8�X�y�ϲ�2?)nߥ�LY2�$=A$6��F!��@���<S���D��.^�C�������Ww���� �C�V]UjB/�[zc'� �J��o0o�r�v�$�D,EU�� `�X��W��3�y	m&���6��@��j ͭ|��
�S9��
����!�+�+���v�Q���?д����d�7z�wQa�k֢�^��q�0��OO���j F5Х��󃶹�W� �c���W�'i1O���y4]q�k���!e��X���	��r�f�ъ�ϒ��6���vLm*�'Ku.��,�&���ڳ�j>}I����X5�-	B�Ѣ�i��N�-�q�'K!D�U��$h�E��M'�,�6��QK���is �T�vu
Y����K�Ur�ڼ�/��c�J��_��u�e�ܴ�8��P�}�7�˃S��R[�Q�cт��Ϥ�X9qNe��&�d���^>	PNz�_��L_k-��A�Z#�~�I��֛j���Ř���R��"6���I���ɳ��r֩�[� .�_r����H�����Z|ٯ���2��	�6]\l�)�9\_h缠4�)�s5�>T=Q���3��1�XW�sc��W`v���뀭�SWՉ=����u�����
߮ˠ�ty=4��m#�`�{���q�e����0X�R��"J>: ?|�.'��LE$���P�j��;���P�g�D�*7�k �C,X��!�w�9��]�r�m�
����ƞ�7uꍘ^lx�JI9�?�^�����<��)Δ����@�~��\_�#��!���?��ߗ�Lsq_f\-�-#;�1]�/�w�H���{�T<1��b�W����K<+��`!�pא�	V���>{bB䛥C[�ʻȺ;��s��ͳ|�f&��O��%��x����L�V}z�r otֲeʞ��D�����Ŷ4�������3����u�@��X��w��V><��9/��q�Bf�}�ƫb��O�G�Rds����P�_qP��u#��g]���>0b�x�ɗ�~�Ú���m��r6�S�B���b���0˼�5�>���M������J}T��t�<p>!=�����pC�������aiy`�㩱և�1I�#��B�sJ'5��g�v%;��*qk��,!YJ��hez��:���kU��F �	����	���Fz�s�"S��
M������[�{�����3@j�<�s��c[�l?;�����M�����1����M!8�rb���ǔ�k����E�K�w]nk�垵e��SN '3:��As�^,[��H�&����gqLM2�Z\�V�3�3~uq���1�J�;鼜c�H�I�ͭ~���Ź�O�4wa�_z���Jr-��$��#����c�PUzA���.�1�~�q+c���:�|,�uSfF��96�Y�'%�����%J&�XI>AVK����+�($���Xv5�>#h��ʥ���Qeu(�9s�1���FK��~�=�ʓ=��>�w���/�5�2f�d��!~�AI����_�#�d��V��A�
3�2Mg���@�D��DQޏ���y\�N��TB>��֟>�{�?�����Y�a��D��=��U��W$���V֚L0|�5��L-�q��y4)�@�
��F�D� ~�K���PĻC��%%]�!Z��9��c[�w:�"�4���GH ���h8�5c�����$�睃Ȯ���[f�]!��7>�����_�e��7���XJ2��F��<�j�&�n�n/��5Ğ�H�����	�F��"x��{�'��p7������ը�VÙ�]��~f�}~�5��!��T��A�A� W�AK9+���P������9�9���u.�m��|���Cs���[Q66m�r�o;5=�/e�����F��R#�H�椝���E-{��2f�aE_4���g˖�\��fj%�po1�ZDi��kQ �@*�1�&_2�
=ߛ����C��^���ۭ��/�,3t(zӄ�N���t{��`��p���HV�!v�lFi Q
�g�Z���L&s��C���(k�T��Y�i���hƄ��xы����ff=������'4lN�EB��	���6�bAt��O��������9�a���Y��q�4���*��#��賬#������������2otĻ�<Tu�P��i,�~��\Þ��x��{d�г<�C���Lt���J�)�=��f1�݊�D�:��_%�8��ȶi�:��+uk{�i�ޠ����G3!�^-�{Pb^az=����}��\�:r�U&�/�U �	�X�a �\��8u�^D�����(������q�!*^A"�u~{���k�69�9F�Z�����b+�,�̷�i�k:a�m�.��fe�[1SR�_����V*�����5ͷ��A��]'<"�M�h������f�������i5q��Ȕf�4���>IkGN�i0����N;�����D��:��XK�ﳮw�
��;�����2�4�Lڥ�WD��RhAY�N�!m�+3«�&�Jc���u�k��2�F��
��r-]v��~�c��Q�s~�:����N�0��6'P��cD��=���A���Q�?�N�&d��6���V�
~P�U�d;&�2�;��Ĉ�-2��L#M��*�G�)�Ēòç��mve��1 ��q�h�zH�n����39��l�F��c��['b����P���`��q`�9�B+�fY�y�h�;���|7���z��I��Ȑ��uZ��Û�>�x&��k� ��M"��M�	<z���cG�v�����i6���n���٫O�sD1v
a�u�^��!!�"94�g^2d�dդ|��߹p��dijnT s�F��������4?m�����=
O:-�CN���@ \5��RF{Ԙ<6�\����(1�:
F�*Ƽk�P�-LC�D�L#U�٧��@����  �͉��z��Rv�#MyK���1���/8+!f�>��wV_�s���0�8��@��������-dER���%�X�3�P�]�1�1��`���9��"�2��H�c34�బ����0.J������v��|tߧvOK��FZ�-op���E���. A��OTCH�4�����E�����x�4��,�J䦝�'/˿X��a2C�&�8X�TX�y�����>���}�w�t�2��5'��jVͲȥY׺�G�ju�S2*0��!����\*���rO+5�����
�m���	�3G)���"uf��w �s�������
'��M�����3b�& ����'�#�F��"q���e�򫱹Z���-ڬi���pV�,\��A���+�R�u؂|h��]I�V�e�k�W�������D|��O"�Uʄ���ܯ�rv}�����6Q�o����RnIf�o�������#@ˋ��b���U�l&��T���	�8����Ӥo�m#D�
KB���u;~j��xszi�&��D8�mv��yc6�
�G�u�U���'�1Bv�� [��8�f��%3**ࣷ�8��5���涧���ot��/k�ɍiy@^�A;2R	`Ӳ��m91�R��Z~�� N!����!�cQR)8g���⭏(����-��)L����c������H{�+�d���
R�5f��cq�>"/��qIN�}�
�79Z�<�K�8�Z,k�͘Ŭ�]��JK�*���Ӌ.��ڜ�x�#�{�*��H���-������ ʩ9'6] �('�4�}�X�|��K��ז�5�R�.7�U7l� �f�o�@Mwo8�a�er��MyrB����Q��L�>���dDv^1`r����%�20��@z_�e��*�>o����ͽ�!`B��g��a���(�!A�GZ�r$�ԃ�ȣg�Eo���#s���s=�Z��t�a��kʾ�qv��ND�j5T���u��*�;�Q
�{��\Xkξe2���z���w^�i9�X���N��1�v�֙h��o�m���{ė�4>X��vZ��3N�aU�@�J�c�iZ�IG`��>3��.#��xC��K7Z�SFqĞF��t���y�������ca��n�*��]Ӫ�%�yz;�Q����c!�l�����o����-��'_���G������x���4�{��G�q�&UABQ3*�g�{る4�j2<�G⑳���?`	'����"�XеE�}�Sg ?t��H�x�[]��<�+��zF�mԳ��a	�a��Z�o�S1r�
�&�xT�~�����=^�bx�<��=�y�IK|A'|��i����J�Tfw6���D�0m� 3kva�maQ^�Y�$�|,�V�D?[�� !B7`R�`�$��(r�ѫ��u~sF30Ṫ�?K�o���dHf4�i���a�n��:��/q�ƚQ��T�u��c��'pd�`���=5]mU�1fs�T�n��tz �>N[�v�wRsn�p�����Ed�(��hm� ;��v����يv��"X-�D���ӂZ�K�P���nк���9HQJ±��ʅ���ϻ`�(��m Y�$9�ֵZD���%��]���ݧ�a�R�?L�*���s�@��W���Vx�	�J;���}.�芅G�6PLjb"����~�I5/��M�m��}fk�#f{��A,��\Ly�zg��C@Auo���n$P�U�zat�<T�R"�������S�c�wc\x���:|9s=�s�.�Μob�7-YJ����i�g������Ej�ت"A�P����,g��c��IײV6���F�M~(����$KT `��I�h�/f��.#+s:Teԏ�`�����D-�й'���f��	��1�1�#N6�S�J���s��M��))�л1b�<T���8'=��	!��Z���?��-��q�C�5	n9�0��gϱ�\ 4%�Hv8\4r-��	,��E��=k�_���x�U3daV^��6k�H}v����S�*4$et١�97��@�k+I�\�t�t8���ҳ�i���8�V�j�FֈFDڵX�]>c#�	q#>�J�m�GV�3R���]$��	xk��j�X��.L��w'؂V���������!	�pk���ө�S��0�88tͮBVc7����t��(zFbk!�IԄ8#��������
÷(�X�5��3<b�U[�X
�&-�'�|%9�tU��o�CܺY{k��Ɋ�r���2���]�p���f�F�MN����\�G���x=��+΀?��c�c�Y�u-�����xc�D�
VB�'o"g0-��80��[+v��ҩ�M�o�Y���;Z���@���X��}W]z� ;*�b���Uw�6�5��F{������ߢ�|��D]S�5�gB�O��	��U��yi=�3m�~EI}~�S_L�ֹ��������pOA�M�8��!`u�Q�v���Z���s[I�;�Ƅ!>)i���l�*&}�<0�k�TP	ކ��J�˶�p��/� ��J�� ��^e0Iw&P0�J9�Y����w��d8f)��7�?��7eNd6�|�J@�����	/Xd�@j�ߝw��������*�I⬈	\�e ���S]o�X��z`�!�,}w��n�G����la[6qO�R�Xl���t�뫦É��Ց�����A�!2�b\fR��I�i����j�x������`A�=�Kmq�S�^	
|s8�]���Lr$�"9�)�_�q�v_VE�|����ga��g��c�$(���M�!KD�kW�za��.s���H���X�b�i.w �I(��R,_�3\;q�L��|Y�J��
��1�Y�J�9<\�(F��O4�����÷}B
�[&Q��t��$%��M��ȝ��lD�-�lG��(E�c�q���G
`�a0b�����D{T$ף^�q]��p5�]E?�U�Θ�����oԙJ*k*�-�OuY��~�Z��*4�pa�������eZ�a�h�H������6O�'�!��n#��!�)�]V�t?��r�y�4��������h�t�۷F����[:�p�IZ���T����4�'�`O�/K�����̙}j]�6{�֡�p�;.C��r�S���<ݦ�,'#wVhB�����F-���BF���s�/À�p�k�[�U�O\L��^=��J�t��j�A����)�W|w�m����ROH�nHk2�{a�t]j'��H��0��ی��b��Y���Ͽ�+�~���D��(+�i�����Y�s�����hy� �W03a��(�γ���Zl�'�<y�Kf�<�z4��ޛ[B�0Y��0�K��@P'�j���w��?~�/���{�a�İG��e�B�^jĐ��$�ݐ#r�}��Mb���	A��Ȥ���,B�b�x����%4�N��'�����LT�6!��/������V1t���g n�,�z]��	��� S|�W�D��ȅ*�E��D=3�{�۹F..��đ�'*t�5�&t�]�}8���~�ʏx!����ȈY�L��V 2�s�Co�u ݠ�uĮ������X��@r�YB&�\���?4V�tS���i���ݜ��U�hk�&7���+�%���D+�v�f ���	���9�\���eoΘ���t�����H�W��H���x�=��ˋ:���_�[&)���Z�&� n����A�fJ���ys��v�H]��a&U�E����T���	��" = Ev[/���=�>��!�Yl���{��n 5O�p���F�!�� ��󜗷X>ïY�]��X��7�Cg3��� XU��Oo�oDh �K�"�7�R�)i�q����\[\�YNd��v�Uщ�7��"R�m���d��q���O�e&�v��;:��ԫ�(6H�׆��#v:�)�R
��$����Cro�,CT���>��,�W0�ע<�D�C�TW�i��Lq(m�tD~�|a���j�=�)���>ket�
{=Z��;<]:P
�:�O5�����O!p��8^K_[��P�ĄB�"K��u0�t��A��� G��15A��GCK$���1��v�x=�OFX]h_Z�#�;s��,��ȹ��c�AGpSR�hW������A}�1t7G�'�Ec��і�s����,�	*��Dy�[zvӯ�2/h=�B�X�D�yDA�����Y5�V�@���It:! cA��H)�X�ӛ7���羂b��dJ(!bWAgbUf�.O�Q~���^���W6�!�D��Bх��'��R��j���;�$��d�аu>MC���eJ�V�w��μ��*�{���9�\{vv���e�g��b���M`l&*�C�X�����V��wM�
����H�%�����[1��%���+L?δ!L6�m<�P�q�NX��B���s��^tQ��[��k.�nlE�k�/�k���'W`^ɒIЍ��\�h�#��Xkd�EM�o�0/��GՅ�Ȅ��nX�7#DG�}�eb���"ךz��&��&s��m^Y�^ə�Q�hP�J͘.��8s���}[��(�m�5�o11�D��M��T�QG��y�<��K��)�19��?�c`_Bex rv(+�즎YGk�E�N_Y1����9��t,� �ɒ��qƊ�i"|"|�nrӘ���kx9��%�z-e�1w$�^.�rB�H?B|X�q$���P�͊�J����a������_�2�E��B�)�Hw*zه0c%�
���4��Lb\�GW�oᣘ�9�8L��c%�&����P1׆c}G�I',Z$vd~�E�~0fjF�Sa��$%=e1���*裈1��V���?�)c�J�S�B>��\)�p�� ��џ1Y3F��9�5-����[�=I��+YRE8�ag]l�M�8�&w}�.�n�Jz˖��\l��L�2��$��?�}ʖL� �չ�|�87ܣ�-���J$Ӱ_`���>����-f�[y��Kl�L��f�:�ߺh������yd�4MN =�ݜ[��)�׿tw�¬Z.�+�vX��X��
��~��5$N�4��E�˷K-�Y�l�9�Q��Z�
=�5F � H�\l5&oy�D9��w�|����*�8*N�EwI��iG���<l;]1��x���%�w1�^Ή`��K�S˝�,��2�����u-Oܙ��� ʐɜ���[bh��Y�^c��eX�2�,��R��AM8�ň}rF�y+����k�Zv�3/�|}r��PQƈ�j���oZۦ�[�����1��ɔ�,Op��ǳ���;��HE�����?�Lu�5��CO�X�b���Ů�D�7�Z�gy������ߠpUI��&�Q���µ^���� ���T�>\����vZk~����Uml&�E&��E@���|J�ۇ0�p"��çH�9'4���[)'�]�LH�zq��a���@��&B��!��������Zx��H�Ia<�ْ��;�J�gG5(��:b�Sۘ�
�oS���A�H�����/@ip�Ť8Ġ{�ّ�/$zT��{�9����~�d_H��� oG�E�b�M��B eaT}:r�b�y�۔_D��%��7B���P��$Z�ѯ��a�������r
ɧ6?L���:�"w�Y��C�(�������V5]��$�g�@lm��x�Cj^�.ecNBB�Q�=M��e���I�;��"�-�B���6\�}���5x��Z��;�����rgY񈹉��uG���wr�V ���
�"��P��wBU���fU���mn�h�3ɑK`>0��(�TJ�)��h=��]��\v7�#��}���>���Knd\�;�����5��;=hK�Ȓ�
�8���
�=���U�k�ى",�r��X�pd���)�^A�}��������'�N��B=b�����f	9'�_��n�>eʗu4=�Dg�"z�k����FJ�г�\pX�ۥ����t�L� �O������CΡ�׾٬�� LL�&4��\Lf�C��rKoM��]M뒫���N�o�����O��G��1�3�}Un�p�"�����9*I<'���}���9l�NW	<e��u-���-�������W���taَ�*F��X���������N�f��[v#N��q���AT�D	��xy�ؼ!>�c5|�&�/�Z�h5�^'*-��J�����?�9���S��|���R�[�x�g3�)<�f�_�d��@�&�������U`�s�7b�xO�`�}��M5�83V6q^�ɷ�¬�Z�C�F5y6�a���V
�S�����(������mQ	>"���0���<�&1�Y4\lؙ�"E���G��0�m��F���S�z+Wו��L~'��nk�o����Z?��>N���ǉJ%�OG<��{xeA�9�J�YnB^�5��J�6�TK�W�U�ϰ�8癢d�ln����n���2��CR_���=LDr�--����r�3πt�w�5ޗ�~�B���y<�R��斟��r_4�ʛ�a5�Y3�%��.�a��ѳ�3����gq���xq�9��5'�&`��Vb^	�~��-OT�6X��]���ur�s[����s�+�>�^�J!h��ؔ��؄��wl��΂��q���fN)h۠,��n��iG�O+4��l��S�7h<%Y���Z��
��5,�������Ʌ@%G��0�K�������{o~��:�s�8�:/�G�ٵ�o�yc���;f}72ճ����)�G����}�u��WX���vdF����z4�{@D��.J��>�zk�G������G}�8C�b�`q���F�X���=ng���1^-���On�
 ��~��?x#?;�Y�M�]�1o`�y$����A�ߦl�>>w���#8��,r�-�k�%/7�a"��_���i�*>�αJ�3��
��E��9/��TN�B���0�`�~2��RW����ѧ2��$��J|PSC4�a�4��s�.���b{%�w �>��o�]�F�p��$C��hS��U]��K�;4����f+֛^
�R���}�k�^��(�m��t�3l��{q��cjS��O�I\w�c�:<4��8�6����:i+����}k�c�9��k�ׯ�������ͭ|:� ��w�D��]Z2�kFEk��t�_�z�5o>�z٭_ �(��'&[w���Ϳ�)���G�(;\'��ْ��3Ȍ;X㪚.D��
�_��b�+�����g��v��
-��A�(�d���_�59�0W��h�n��t����>�/�b:�3Kbz�5J�Ĵ����٘#����̮�jϵHyc�k�6�	�3d9��	k�0'1L^�����y���^�/e:=MD�c���a�M��2�	�|X���A}��Tڽ	���P|dg�����nX�D�]ʌk0$�:xcS����V���3��s��)O1��&v9"�p2�=k�p5�P��g&��r5$y��Pqcj������^>�T�L]�PA7�੕��`�M6RPm����eC!u���)�d� �2��+�P ��)�f�q�k¤5��EjT5"I�I�!	a�ם�҈�A{�܌�<�G�\A#�P�er�L�s�S��l6�S���g:�/>�]?/۰�G��/��VBrމ5����5�l�=zU���	���xj)��E�;-�:%��ZD��'��@L�i��
��KS�s��$���r�6vY-r��?,���,7~a�_e[t���͑#� Ag�-�� BYK% ��`Ÿ��wan{���HrY�mֽ]'��|%ړs����
xI��iG8�Ϸ--���ZH�>V=0ʣ�&Xʕ/i�uz�i�v�&��ry`�(V��#X��)�OM�t��=��q��Gx�#F��b�v��5D.R~�5l�U�L������n��w�JʃMk��ձ�� ���x��2�v��
��G���p7H��?�/u����o�f:(�7�����8�EL����>]��ߘ�I��Y��-]�'�����f��mY��'g��j���d��޹����{����H����뤹�|� 1��9}do��)D�%���w悽�Sd��Џ���J.Z��7����Ͼ�((���?c��Pw3��ZܞxJ�� �U~)۬,Y���s�������o	7�J��v����t?+������k��[J@Ϸh�����F�CX��*�f��=Q�α=sG��YW��]�ז�>˖n��/�.3&Ƶ�"G�lA�F�)��Tw*R����+��&�\��k��?0�7�O0������	���'�����{H��[�<G.^b�a$荅%SvD�n�DY��M�8���)�~�Q��䢇�㲨�Bp2Z�\�@9��n<�BB�-�����|O�ô���f��1��
j�t�������zN�s|���}��[�hq=����itsU9vZ�T�*ǻW��ٝl�Ow�yp�X>.�)�f3�X��od�+�
�V�k����j2LsK�ⶆ�cQ�S�K��3QK�n���w���s{+�hݰSǝ���m�K��C���T@6\�d�3�*�b@L�^E�0�_�o�Gd�J�+0'�좝x�7M~ -�~�j0���.�����S��F>D褩\�]�,�f���(a���P����[�����'d�Q���\�)Z`����O�t��?��;-ƣY'�|�)�kb��yLo(�	L���������)��6�݌4s�r�}����2XI_(�����_�ԥ<�$T5!ǽ��:a6[�#z��G<Q)���l9cM���K�-��/#�.q������D��0�t����`ɜu05??���]��"1z $xP�{L�[\�Hi>�=��̖��=(����	w�~����(>�FB.B�� �J�X<r�n�L��EP\�+�qO
оri}�0+7^����g�i�J�BR��
��j��YU�Y��L�a3VC��G!�U�:��΀�G������ř9��>.I�|d$�h�(t����v@m�m]S��[���li'ᮂ�(ҭv$cZ���eZ/"=݀��L�S�·hl�����5g�n!�0-��1.��Zu'�T�928;d����z)8i=�v9��^��RF�h�#�.�pՔ T��r�V��O�-C\K��;�T��r�5�{�mc.*�
�i������
&x�Ӕd�Z��"�����H�
��!Μ1�����&�|�*
svA2�r��<x?�0T������8K �Ps��QP��<Eݵ}�Bb��?��;�s�&�XA�!�7%$��MȮ]�
�p6l�s`w� Eɑt��G�~uH�.T���8{܇{mW�&[ 3z�K"���)��q���2!�;ʰv���q�2!�a�li�j_c�z4���2tQ1=���M���ׅ[�����&CX���0�I�1�J����iԜ��/K��oSє2�U8K9�� �l�z��*�뤉�&9���=�@
HVW�4 *�2	y6�G��S%.}��	�$��E�>/|��4x_b@V`u����Ӊ���R㸕4|�U�K��`�m�5~m��|�8B[������t4�
�^���=bg�@)���W��������Y+<:=o�]�㓂��޵�k}��G���Ϝ�(�eC�	��_�9`z�Xl�� |Ъ��Ų(D��'ᄼHi2�)�	,��j�Z?��s�:�
Fj��������cWj�]��P��X�eq�����y�-V��k/��g���Z�_}-����q* %�j�DD֦�l	�^}Y�UUَU$�E7�� `�W�p��T�3�R�7��ќ�ȅe e��5Ⱥm��7�T�op�� �P4o֓�U/�mBnQ��W:3���*���ӽ�	�`�*	�]Z8�~�;�ٙo�Z��3�<�$%���{�jw�(� �t���GF�S3���������!�*�򺃎<��r��z�2����V���O"N6�A�P��w����g�F��=5.�
�#��E��	_�&����I0ӒFp�i��5چ�i"��=�A�n���am��7O!������M4���+e{@x���� �VX�Y��g�Ɏ��d�C(�2\B�-z^�d�@����n;�t�\�-�����|�Ԧ�B$���	e$��/m4�BC�/!�慎A�3��+}����/�{� ��)d�!��|[�����n٩�/}�2\&$ݖA+����s;�ٲ��}�F��ZD���$��vs10|�w����J8�Ki�7���_��} �֌�e��#����q?]�4h�_�l�,��2��Gޘ�6_11��d5A&�bF�Ӽds�S<�ņ�M�? ��=���pI ��sŁ�t�:iP02��L6��)qcj�Tq9C�V��e)��K8ƀm���4� �������5��P^7���x���A�<�6򥯔lt�;~Tv@V�@7\F�?ݼ!
��A�~��6���w���9�����H�����ar��=�f����W�p
To��u":{8��)�~��0��3rB�6�����A�ס�~�<+j��M����H��P�7��4�u���Aqs�1lR��i�}B�sl��F�$S�]%a�Z�x3�Q��$8��`v���*����Hc�X�<��^�ǳJwբ1KO�%bGd�A��¤M��|�!��F~d�E�����еP�yĪ�����/�ޤ�ݺ-���D�+�+r5v����el��U�#��^��7~�xq�A�yh��5�&�#R�q�	�f��rqK��V6�Ԃ��c�&����Jėo��iX��ʠ5��&WvFW��Mi,,��t��+.e���x'���/�J��B��o\|�K���^�h��)q��m�m��8;8�����܋}r�,����E��qh�� ��I�/:
d��Q��
2�Q3w�C�j-�C����ƇS%��Iz��;����Cu��^G�
Ik����gCc��V�A0���_VW+��$��L����,�������K���'��OQ��؇d�n�ng�½������������ȇ�n�G�<N�r]D8`�O�K�:,�;��ɀ���e�!���5�L�D����"���h��t�X[���x��W���7z���J�{Q��3�ߠ�a������de-o��v�����
eP�l�0ǻP�[��~�ڛyP1&���>��z �R�b�/���V�K ���H�?f�����;���V��! �:��������?�xU�f>G�V��w 1���8n���#^���A*M] "l��ㄤ:���gs��]�HL�?֤n���K� ��6��y��k�50���+�l���J��7<���=�ҢQ�7��ҏ�
5t�@�
�%:�w�Ӳ��(km"�n����|b��i��Аu"H��Iy϶��KE��T�Kn����r�f[�7� `�q�9��X��/�F]�X^y��v�ڿH��;j�P�,L�9(�5Wk�sx:��5��SEa2"8����>��fN�����Y!�&��&[%��kf�Q�~��۫��m������K4$л�����_V.�p�Q����]:��;�	�T��T�ɾ3@#x�m����E�<��I8"Q֎+0���nݏ�U+t�?:�����_@��9zx�E-������hl�:'�4K�p��M�n��Hô�D�8
��^>��W"��T� �O�HfH��6�9�>��SOJN���	��} ~��cbV
��#�+yZ�gQ9'�[Y����}:!d=p~C��7JŢ/��`����DV!��ݙ�̙�����@���Zد8u�)��Q�3�^�BZ�>��וּ�'���c�����n"l:�Z�����>�^cUD�@0���Pѥp���fЙ"��I)������9���p3B���
�*���0>��P��",�F���$ LH���)�JhT��I��ݸ/�n�$A$������yrU}F���8���� �+��8�jh�m��晁r-`1}ߤ���$�6��-����󉾔䑪_P�I�J��S��	����[=�(���;���QƘ�{)M�T�5葻�m�=h</m+p��������-1�Ia�j�d��1�B�Tq�i��LNuL��b ��X�_h)��e+#��zD �B�BTU�賻�1��77=W��A���%�8��J����\�S�T�� QPBR�(�sTR�M��̪�K����Bz��1���Q����鲛��6��R~�!�?�/��/�	�Zw�61UH�֋�_!���fSmh�C.k�=��9#h��r1���]s'�OlgK�b�� !�?�,�'�?j*BkCxUb?u�\���.�B�����z��R�Ȗp���aB@j�X��jB���������@�WY3�d��4lQ'�-�{���X7/�9P:��9�]�2�	��L��a)1�U#�9T�U��Pcb��<��O��HKM�J��G*97�h6����~�	�6Q՚2y�w��q�f�3g�	��wA�"�彽���Y���e1��۩� ��b��cɴ�if�r���Ep�w�G_�%�8S���k^��++R>�KXtv�+��k[S��!ٝ3��=���hL8��1���:		`wd���eu*��6|.ٯAm���x6������kQ�b���2�\�9c����p���	sE;���B~�<��:�0�/nfz�V���'�x(ye�	�����&i�M)qg�7H�{�����,D)���K���
���z��	�޳��s�;�b!�>qV��KwԸ>���=���/�C>��`� ��<X7@�E�3~3��7��_1:��c�<0���eܴ]�?��|
W�n%N�V�K��؜&FW��:�W$�փ�����3:V�(@�����s�8l���V�c�T/�Q5��eBKќ����}� �AK�H��A���;�GF��r�`��������;��p3�D���|:Dr��v�V|V4�����
�L;�JsHmp�	G[^9s�/Tn���0)#P�Q7L��g�k��pq��dV��8G�����R#���y��w��?��T��P��Ͱ ������������S��? z�j�2�^؜�
}�����z��m�ҀH����4�l̩�Q�C��5�޹6w�@��ӑv��w��ۊ���lL/�1۾2�J:�ղs�v�ѳ�l�0��X����c��9�.j"'"&�~*{�"sS0�|�1yw�s2\�ڡ0��FL���G�?|�X	� 'j4L�5Зu��o��N���P(GH�_��RW~��w.L�)��ܑz��/�J䛯�&ƨ��(
%�e�n�=f�%=�`��&��޽�4=�yz>��N���3{V4$� �-"�~. P��^��Q�^K�P���m	c�R�/��|QX���B2ۋU��.�'������ρ��|�M�[v	S�]Mt�ެVs ����Ӣ�{�d7�	��4�n@�pw;@=׼/��ٙ#}��z�].��vh�5�)7�q��MM�FݟE5��.Ho�5�1T�g����2����[b;]�La��8�Amv��R�#�ƲR�}��:�qY��F6�\S�L�Q��������٢jؓ�B����� ��[M�[����-5�4�9M�*��W��a*6�K���87�JX�.�J��Į:"4���L�M�\�w���R�!��-V����5�W.��i�������!�E�B*-���Ο%�~Q�K�~φ���z{&K�ܟ�k�2�d��27l&lA]kޱ]��q_<s'�.!IL��窒Om"�qv����ӂ���	aUq	/�W��3��>W�E|�w����o��b�ZZ��Y�5�#!o?Ge %���z��QDHܙρ�YPV�h�?�/��:~����eEĶz��.Y4�}R�-&bE������{��E��@���Q(kvN�̼�����d�,S�29�M��гJ܍��Kʬ�x,�-��>���7\��[���p�*�X23��������\��9I���qAey�IE��>�����	�J__��#$���j]n,tͿ[�n� ��K'�@{D�)LU3�����6��RsAM>g�͌���}5�6<z�x������.��R�v�[z�o�	K� |՚q�k��&[V�-4�0먟2%P�nY�Ҵ%Y2�$�m���Z<�^T�v�HF7l{���|�EC-��Dӵ��<a��Vz�:]G�5�P��Ʈ�0*w���c� X櫅�Kߴ8>!�7G_�8;�M8�z�	{y��M�db]۝��:�V��pB����>�X��w��+����ՙ?h�|n�6�Tz�{������òWjE���[Q�Ϯ�yS���%�̠��A��J!�6$;;��o��$���Y�Jj5�xf=gsD�K���;�C �@'k �]d���y�l�%p���t��Co^���:�	hYX�m�@m�>�y'����@W��1`T��M���q�t>EЌt�!߮�7�f:gu���s�|�ˈ֤��$)3P�����ܤK�h�uN%g�g=`�R3�3���4C�A����^� 7��)�?�]�^U��DE��X��N3ĜC���x
G���L�67"h�i��b���r���Oڊ�u���ۛ���.K;�ڃ�T��ȫ��w�Ć�|�ߦ�hUL�j�ڷ��m�u��	_>bc!]Wk�2����嵹t�,�BI���Fֹ��Dn��'��Va�%��
4�K� ~�'���,}�W��|��ĝѥ�k�� �z�7���&�]���=�$�=
	�Z�^n+���-�q��R���k?�����PabL4fT��>�����+� l=Y���r��I��N�������߶��BU�E}�-�	T&@o��r[y��n QǨ����ב�3^\��左-��M���`s������ò��;{}�vc2(X= �e��r�[���!������<Z�KӮ����Yq6';�	�� T�«��]���B|�3����5�h��P.�eD�u�u�bHV}�����wT�J�Z	�I����?���T��r�z�T���i�R�%==�|Y,nKi�A"p�4�d���B���scv1�q�\�D��?=RVש>y��ȿ����2'�go/AL��࿀e:�(v���K���{�%�J�̔	\���U��W�MM��Q�WT�<����QL�|v�6n�zV��
�oꓩ"u�������}#^"��aC�9�F�u�8m4�#�&�Q?\��ř4�Pe�*}�ѿ�������b�t�. ���e6
����u%[�����Lw4�δ���h[����ɏ�VR��f)�n"�F#�Mp���$�'�۹�{�_�<Lj�tpOE��|�[�'"p�y�i3r-]�D�G��;���D/S���4!`�Ћژy�5��9��2��9BꞱJ��Y���dD�@�
0��_H{�v�MSyˌ�S޹w���k��N��0�ukќ��8<1^����[���2��-x��o�,�d:+���?�w&WK�$�r�l��F�ۻ��Ѫ(M���Y{p�����M�z!QA�	{s��yaÈ$A�pQ#?�@)f��:Q�0��U�if[�s�s&�F ��3��jF��?��Ȇ0����
��Ψ�*������p�"��F��jfѮ�#�����'�U��s��yTQ%f��Ľ�����B@��`tQ�O�3��U�LI�t�'���]��
��^L��^����yc-z��f���ĻoK��|8�l�<��*�����}Q��MF���C�ft1q�
B��~UQ���*U\�6  �DNT> �2�:��O�mW|Z�1�1S���ҹ�.k-��`}Et�$͇�Y+2�Zո�F+��3���Sx��>�� Hֻ�ج�����%�I�e��+�,�A�NG{��+��^*Vpx��T��g�22G�ʕ4�K}�^oI׌�e�i��:�a���B��G�(���TD�u�<����7����g=��đ?J ��Q��b�-2BC瓕ھ�/x�/�O�1��`n�eH����	j?!�5���v�kӲ�Z'F	���$ub�s���l?��RD��hyyg�b0�`>�a-p5-m���?���M;I9�L�%w�)w^����֛�p/� �P<�_���3F�>������G�	�Tn,����5)�Ln?�qɊ;����7��������6L�D�z5$���J$�P�Q����U��Ğ���@2�*���c�*�=�:�"���yo�pêYH�KK�n²<�_b��?a���+�u��5�a6�
�P=�1(�zCuz��B��X�Oq��/Fi�T$�{��0��ԡ�c]��N|iО_����R���4j�b����~i�L�b����P�|�,�ū���k/�H�ր��{4��P�,���t�:��Ɲ��`bF��(bgy��d$��UH��\���Hr����e}�����ɞ�w�5�s7� N���) �빂
��Ә�A���d�V$j�ĭV.��Y"I��=��T_mg(B�Q2�Yk��9Ϳ�e��ĞJ_ԧ�Z�Y@R~�*�:��O�����_��zH�v\�%8��� ���r�y:���ڵ�!l�99S!��v���y��j�J�QE������O�
�]s]D�R�I�<�ۚ����Uc�p�irM�`��-��"v�h��z��zRo��T�ۣ�`�G1�JJ�:�f3sS���y�T)j���>�	��/�%O�|\�O�B����|���Ue������2���>L�Ԗ��l�;�[VAJ�1�>gZ_W��i�z�Z��Wg�/9��+�V�}/�UQ�IvR�l���?�>�7�?^�9E3��M�'��R@�����\�x���m�6x��	��`�8sΓ��ÕNBZ ����)�$�N�i��Uj7n}A+�/�k�E�6f�7��R|^�M�2��<��N�ۡ�v�N �*\TM,���<E�����h78�-��/Њ̔8$�[ք���	�\�_����{;��R�+�pC���e�Gn�^��1���=tLܨ(�6�SCd��1���Ȁ�2�������<h �9�_�O*�B��!�~�;�G��y3�a_x=���t@v�q����*�I�(�I��;������u#@�Z����T
h��C#U1�C#ɚ#�T>;!$a�Aێ�9�J�4�*�߄&����h�ߌ<D5؈�#"��5��~d�l�9�[�YT��F,	���
y���G�t��7� �(�g�v#�:��nT /Z^6�gZ/�g�g`z`n F��:�=�!�>!�q,���}f{o�r���6�^���y5'�����nj1��z�˵:x�Eք�r��
�2}��`ɲdW�X��#��s��v����:����y�HLT�o�v���b�Dtt����S������|>Iio�F��E��X"��c�da)~���N9h=u�� ���Y��:� z��f� ��{r�a��B�(@4t��=/�Є��hw�=���db�����71��L�`��.b
r� 6����rP�>�pQ �K��)��:���YX*�^�Z�x����B�iʚ�P��f�Y:��--�,?ܸ"N_a_az���Ҟco�������Qt����Eș�	7v�mpij��Z._��Ig`����.hu��&rC{��j�p͗��dG��0�j��v���z�ū�l踔�t����9�tA���aCٜ��^�֨^<�r�	�O�M��Izfm�p���5���������(3+B	�X��P����@P��Ր; _��݉�pϕ*�d��C������MZ��	ȴ���q�u_�ffd]��^� �э�O��L�Ԇ�f�j2�fRpȆ��@��3�W�RQ�,bY��lp�fܼw�!R(I�F��O_�t
g���y��]��Z$����J��z�:s��I܄��|ϧ���>(h���|�k'2�t/���&�j�v�����®y����sf�)��*�Wn�A�9&�dw�oA�F����o�l�ؗ��_�5��0�m��K~�.�K�r�
�y0}D�!7����y��A��,Ξ�,����'(o��߶���8
F^^hC��lv���,zժ��uS�<��~=#��}Q���@����҂���zS�-|�	8��ڿ�s�8_Ԇ��Eu��U��<�e*A�� Q�{���ב#}=ӛ��[wu���S�����Ϻ�	V�n�}��`0���!yt��P�X>��jƐz�'�0���d�oU#�*C���R�.�����dY$Aodv��i�g`�(DU;ɻȌLFQ���Bq�\'�L_��Ha�o1�9�.2�����������f�����F�y樧�hU6U���l+�/9����s7cr�B�{&VO�9��g���������E���e�����Q���}'cvY�I�4�]��:�0U.M��I�mH4�S��q�:TQ}P�����!x�w'�u�˜QV�C_d[fX�3�k�Q�#ӑvd�E�"���Ԉ}�iE��C��:4�w�h�Y����v�~)���u|��϶,�M#�P�P��o� �:�ne$��H�%;t5��{���Ti���bL���*�{�}��>�)M!�*���������p����_ U%���@6�,�+����D[s!�
�+2�z6�.0���Qz���
tH�hC�1%w�QS_��M¦ Q8��%��pހ7G��9N��誅�[ڣ{k#դ]�Z�f��[Xw�/�4�p��6����dcƷ��m�=�������Q��.�����P������3��L��y��s7EA��Xmw[ͯ�/K0��.�t%����M��+��2N��\����1�-r1�j�*���i��x����n0'T2A(���u��έ��3�ӜA~����2۝���.���7ˁ\�̌�wd G�BS(���1p�����Nү�~[B���+s�)���j��������qo������I:`�����E��Rk)�ײ$��r��V#,6;���;tr��%��`ǽ�='��W�n�m���rM��!I)�KK��5��Z�q|�*�cW��p����B����>�V6ږu)�ל���h`P�:D��N��V����>V7?!H�j�"���07�^��-��������$[
�����<��aʻ$��P�g!T 9��x��h7���{�T<���:G�<$�9���s�<ЉZ*�Uz��3ɬd��wi�,��Qb�;Gۛ��$��єT���"����w9�Ԯ�0j�좮�H��[�6�(�~U/Rׯ��� -��ʶ*P��Iw�͟>�b�hhط=�j)�g��#"��_�0����R=�L��/�a	$c�+�O�4��0�/���>Pi�Z.�::�8�Q2y�i������3<Vb'���Ʉ��a[��0-�[R]��Y�c.�[�X6;�V���M��cW�>�_{�`�E�A�Eqq$�9����[J&(j>�K����]D�l�o���@��@B	��$��&sD�q �1�ll~�ķEI��)C���mA�>�\�j
�
>pX�Ǽ��I�q(���^��X�Z�j�&cZ��~��t5��j���u&�F����x�Izw�]ts�.��!�h�{�R��%N;�C.��@��)[������$�o=�ㅪ��ճ�=��x���y:����I�@�������Y��/��b$���z$l�啵�:��������,Z
���(���I]�R��ܖ���'
��>NC����9�����t *�����x�4͚�p�z���L?1��Tu�F�3���s�������m��!��"�T�����&�u<N 2g��\`����{+m�L��br��\�t}�(E����u�u���BG}�H�ܭ�2��Nh�hFk5ZT6��3M.��h
��G�>Bw���z�'E]�Z3�dt<|GO#|ɝ�v
@���|�}��+n��3������>vL�$��(�\j46���vŲ��4"��z|-3w�p$���
YcM��o�=g����6G��s����`�:�P<�*?��������0v�s��b>K���WR�r��2��XCQq�@�gs\9��jĿ�8�ۼIxҒH6Z_:B�"���ʾtgg�u�RMJ�� ���9��!Q���}eݑn��Ϯ���1t����hk��q����Ae���v�rL��K��j*��"`_��H�SZ�gX��2�.p��ĜT,��K�w��:��������J�G[�����4R���7�\�\N�a����7����V#�YK�p-�$+�M"C⊗~v�(��"��p�*���c���٬U1�g�Hq"��<���)�8���]�'�;RS�	�nS�r���DF�BB��7���_j��fYz��:fd���o�.����E
����DE�[ɱ�b��0�~�CZ���-�B̂3��h=bM��U$�g��t�zD�oG�&�k�{��q�w����l[�g��t�X$��x���6���*�vXK;_1
��н���"�!j��\x�\*P��aA$֨���@MmO֡����z��]�e�!�Fw��!��i�ΑW�O��7bsH:�Y�|�}����{>��x�AL��DUn"�K�Y�L�,�NvA�Vn��d'�e��n^Z�헂#z���-�mB�@L.n�ͺ������Lr�|FX[�f���f�0�UU� �5�!,�UI��uE��x1�"��쿐)M����d��ͅ�%(N0�j+��Y	�*�v��11��<�0�y�D��{!��(2��ھyzl���%��/e��f����|�TN'N�mHYHu��k�qQ�zy�؏�˿�;x���mly�t��%���R�T�B�!ͫ����C�$�?��ˬ{Ry��+2\�<B��;v��,e%n���o��꙲/fD���z*�wuuݣ�t��2b}P���M�7ca	T��K���fCZl-2�FmD񵟿�bĦ7��"�i���85�
"8Žm���B2 2?_�ɉp��T�!��BO���3��7�X<C�b@��^VTL�QX���B}��$�+9v�m\ �4�*S����t������ӆ����Z�/�t���r_$f�!�S:@���I�T�G4
t�1���udfg���! ]|��h�,���X��ħ�{��X��g@n��OѢ�$x#����K��p#�R$�Z5��Z����rB0����ttU�ؕ���X˼��j�\�� �iTu�OY��[�ڣ<�#�*�}����k��<f仒7��S���Q��l�����e쾨��X����pBo��BNDA� �_�a+�p�|r+�ʖ">ʹ����%�7�'�Pzx��Ü�87)3�we~���sN�٩=���������5:B��p�'o�hcP��a�)L٪3e������K?��yP�j��u�SC�qRD�a��nM�2V7%Ǵ���@C��֦�=�v��$�g,�¤&!P�p��O��n�\�Za�E���ˤ�+�g�M���&�;�u����ev�S�AC�������{���BNxמEvgq��/��r%��/������t٨���3�R��Sh� W�)��_�aJ�7᲋Y@�Z�w+nDx_����"�ӻ�;4S�)[��)�";7��̙�U��0�AS �_�Qz栄�!e�٫4�%@�)���+�Ǡ3�H�pD�~-��ݔ$��t%`ZX�������"��|'�\J㉫�[�g�����D�[��"p�F�@�V�9-�MD2�.��2���j�锤�4y��I`o�ܰZ%L�ß�U�8�օ4]U$h,E�	EE}x�~�� �e�u���j� {��|�4A����e	Ɗ!�ȝ�8��w�%�rJ�p2G��oҊGA1�η��m�~�7�s����ς��1P�t��t��ڽ��᡹�D��b!��
^^Dp�2_^V�#� i��L��Y�d�X\ݗ�e6X�o�"�/osepH�^r��DO�t@�C>L�ƴ����_���{�Ŭ�j[��n|��y�ޫ��6�L��7��Tqz����4��2��[33H4��e�d`�P��=��dA���Қ�z�8�E%��1y�M��wJ;��r+����}����*L�wKJ��9�yq�kq<h��Z;�Ȓ��`�/�x�����H�ꤔx�%��9"��d?�~���Nز��jm;��
2 �To�Ҍ�;�hn˓ʟ�V�`hL���P���i���zk��$���r�x�'��˼]��|,��y>������ڀ���B,�!굷�ڣ'u��h��o@3�(T�6v�Px'��J�ռh�u,�VsVa8
=�����q�3�Pt(��<��g��n�9���\j�!�9˩�.��0�<Y��W<�8��Dw�k�c=إ$��BP5o��`n��9��.��(�4f~�z�[>DJ��_Td��Yh���������427��*��t�_�w<��Ԙ���(Q-WՏ���بp���I����ULH�[[��ќ��{�2-�����4T��`*d�u�����a���]���)����4 C+���%�|�u�Y����ԈP��"�e���S;�ZQ�� ����n][kp�������P+&=nv��0����=�_]�s:�7iH�H�+ �m����I!�|�v�+�-��j�W$#�/gKMfmh6B�КS"�`+(̆7�8�#�t�L��x,|�lq�9t��PE�Vb2��1��}X��Ub�������K΁��͇N��c{zv�r/&�s��)p4?=�˲�[�?��>���x���C��s�GR�sB��,��Fk�Q��16�ST��W3D�� !�X� =�<%�,-�q�ե�h�C��W��쯇4���KTD��p�?��������_WK��W'�!���8�s)f��m�3m�y0$��F��h���L�Vr�����bN�iNc��r4� &V��Ij_��\6��7�����TH�wJu���f�[!��m�M�􁘭�j�LQ5f.��=��+X�Ï���p��>}���V����N��Էɿ�mw�Kq�}�{�x��гX�˶�)��+��p ߾=L��Whb�&� ��[�|�+�lpf�o��oC�����`�[G�| .bE�~G4�R��$�b��Vs�'��/�����ڜ8�C�v�z�y����$�.R OO\�����9�~]>�����U3�I�w�U�f�^7��՗�����ئc�~{�N�j��0�� !a)�F!�M C�783�FU]�O_�h����&�����:����J�)"�n͈"]{=����R���F�%����]~`(|$��y�d0߫�?�K�1A�WĘ�W��^h��5 �d���[�D�,k�9���)����*�(�~*��&�����{��+�.�,.�@�ưu��Wm�p��Ha�[*;z�T5��d��/-����P��\*��5t(�I�>Pi��5U_5��՝��9[�0�� |�b���'}m��A�x�d
b�CC���K9y����@e9'#<c|�,��6��4򞬻���E��� Rr����.
�F3�S�\"��w���xB�k��/����&����?����V2��-�����#�b7:��QQ�;���dX�1_����������C��Ɨ�$�7���y�`:��4v��_+ݳ��@6�xA�@^�k���i�	�*_����I�+�����Wt>��{�H ƻ�d�H_�<�����;��~u��Ld��5��*��V�F�t�A������;����٬�����3t BM%y���J��xC2g�E%��cb:}\�����aL��NEW*0j��>X!)5�5k?��/��+�o��b��cƐ��<��V����PA�{��|Q>���̀¸�M�dc�Ϧ�0 �	�+�y��W�%�>�<�#�0�d={HܚɡV�C������IASU���ۖ 7��Yh��n����Q���4��m�l?��Ц7n?#���L:� ���aÜ��p���gJ���	��S	~����EO/}r`a�}���Ґ�Ʒ�׹*h��kt�]dߓ`�N*��Ɣe��Lֆi��ɳ�o��_�2'��z�T���2Y� ԫ����]�l^u��[,2��۔#��ͨg�r�3�7]��s�����E���' �[��j7>I|ys�k��A�Il"n��)��`�Ƞ�ˢFԅ��;�dY�^5hn[�7�#s��W_�IC�֮ka�Fn�&�1F�Fͧ�N}O�����4�OL�-}���Ŝ�@��Y��	���{1�0<eG� u@#p��c8��[���:'��
p��Q�QRAaa�Ղ6(��<�։!���½��YX��0ld��ȏB#����(t���酆Z�۶	�S���4��P�0��
� ��&��1�MY��$���W�������0��UM����t� Dq�GF�r
Ծ��Yu�H�k^�>^+TL\�v@��G���:�p��P��VD���1�eC\@M�G�M8�����c�w��<�;�j�C��!��-Ρˣ_�ɵ|�N����fG����1��	��C� �@H�^`�LӚ��u!j*j:k�6�A�ȼ*��8O���2�m��� ��?�z}�)���� PM� J ��.��u�ܺ�tψ�� qH�V�ls0�P�2VQ�y.;�_�J>�m7�2�G} B�0�4W�ta��G��P͒�an��+&A[����ץt����c(]hp ��IN�>��?�l)_Ag��oP$cx�)<JK��m��ex�.�P&ŗF�4�z���Q!�mt{�P k��7��BG�1׽4���8��r�$���؎�+�b���?z�9��T�RWA�C�t�xY��4y?|�چ^Tؒg��:���OG�Xr[�9��W.��n�l�\:�BFN����;�Ɵۚ@�%,��ζ^���4���[I}H� �4�D��p����m��{���=��J�C�gŐ�1|W�U�>�Rc� e{"ě��ބ��y��@m�/�\��Nk�<��%�u��x���.a
3��_��Dt�3[�{]�+�9���{����
�jïA�V(�y�rλN�g8W�ٔ�:V5�Lu7Y�0��|����Bm�|��}��{���7�B����
׍�F�h��)�I8�޲3n$� �f�z3ՠ��=r���s����Ȥ�Zu����֭��R�Rx^�9o���e�Ր�f�Y嵛1H�]jH;]A�
?/M�H��������<�<�|�"�D��9������P�\*�-�^@_P^%�}כ8E�cM�k�o��^���"�
;7��������gͫ�L����Ϳ|�a�SH㒅�M��ge�Ⲅ5-ߌ+t�Յ���Y(ʉ/K�H�����"�'��Ғ���*��gN�S�h�)��8h"H'Bgl)iL�
�=�����V����鎲��(\�5�'o�%
f�S�7bԷ%��!e�h8�`1�d�ľe���,Y����b^i͏�:���D�P�W]���ٚ!�"�7�
�~�E��ԟ�3�ƚ��k.t���J�;g�����ϮjO���_ >Jqθ��e�П?�ِv�6�+���9��S������ż-z�p��Tx��E��`�� �up���\�(�t�L�Z��^���+�d�3A)��0��#�_��ܼ8i�F�����':9���\9k@���ƂڞϦ��$a?�YרF��@p����v4#�1YQ7Q�*`61�p���M��(�+�i5P��E�R<�u���b��UTtW..�U%��'Άh�tr�^E�6�}�_�KÜ��B��q�X�ϋ���_ʰ�צ������J՞�:�J���dS-�d@bd�d�S���?����G��%l�����:S���mUn��A�w��И�0K�l:D�`%f��Dc{��u ��/����a�y-�z%����\ ^x�f���_�1�=I�G��ztK�����4NgN:�U������K*�p�~��SYY���$��?����è�6Q����C9��c�;KէX��Q�^ݑ���f�����zyd�^R6E$/��{@!&�xx���v���f�Ty�3���K��~+;K�3��~�I�W�B��3*�U�dP2,,�� 
ߺ�y_��7vh}"��K�1������W�z�P�#Z)/؇i{�aS�n�T�;�av4�Tq~��%�T������ݮ���mO2��ݠ�	y^���_��ɔ�-*���?"R�;8a��mu��4g;#05髿�"�?}���w�}����K�/g"�S��c"~��p����s� ���2&�Oc��TdptΓ�u3�����.�����f��[��X��s�R��]P����߰<c��샆��^E؃����A]�M�-��_-N�'R�̪B�̖j����$�v#G��.��0]s��!W�cT����=���sK�������.���X����&������)�8e���VB�T��
�,G��(F��I�#Qѻ7{]�2%S�5�L��iU�ٚ([�0�*��"�D���K$q\�ҢZA�૰��^*7�����]�~�8X7׺'��x����= R�E��!�h��)�~I�%�Fg�\2�s�Q)��������TZ��(1����y 
��^�Vݹݾu�rY\�f���tk<���A�	iΑ��Cf��kj�o��g���"6I��r�RMCn��\�ں���cC����2����(n�4�Ce~YH�*�ĳ �޳��TN��Q���Vn�,8d�{Cѿ�i��o�D�p_�?Yd
�uEph�����#a����{"ѹ[�XEe�H�q���;����筬^ky��DHq ��X���*�7����ǘ��se>���m  
L�1R-Q"hW�+Y��L��Y�f��#+	$:���By�U�Ϯfn�1�
���i�'*������Nn��-��e�䄙I_-��������ԡ��.�/�%g����,"�Ӹsg�/'3�H��W�|�.Ti��(j�I��k�����#�
� A��	����С���,�l����+%b
�գ��܍5��;��4�s��9mx��E5�5��Yp����(Q�"ˢ~ݑ.ӇW�ez T��v�������ܲ����ldN�h��_sf�.dy�#��`�9�y��uU1���}+�8�]�+H��>���3[��g?�����Y�7?FAQ1�����E��3N���E�q������km;�4���t���������2�o��)�=�7`͘]y�2L|�5��"E�I��hh��f��2��a����:9Zɩ8�Nē�iP� b�m�if�u�R���kƼ�N@���uȂ�0*��ez�n�77L�����z��o��r���}�پ��)Mt_�Y�ory��m�
�\�9j� ��z2�e��$���Н��gϓ�ć�p\C��t�����Cdԓ�h8��\���D��=�6J��ʥ�q5���f��������@j� �5{&(t k(l�%�s,4�����$�6�c��KO�{J{CK�^��9�<��޳�.:Z3��ў�),2���%��x�-����	J�!��͞^���Nr�����Gq���o�O�ar��ke�H�f7���=pZ�a�r ���`���I�8���/�V���Ikb=K��n}3��^sÜ6|M����`�rv1X�!����؍��
��0&�0�C�қ�1ºWj�R���sX�B�!�o	5]�b�UN^�N���Z	�h��<E�@�Җ�:r1�s"~D�w�rU�99������,�&E��Ddf"5���0POV���Ze���#ǀ�i	of��2(�;"a;۱�ޏ�
c�1�"'h J﹌L�Y)���+1�K�02�^��4�d5�a��H�S*="����� ��$��/�.a��.6����9e%o���WN,%��J���fX�av�~� gh�8ºŻ�{���x��Ǝ�'篴ou�@|�0_�(f��?��"��4�B�2��so=��JJDP������p>��`���c�ކ�zI�-V�UUn�O왇߾�$�Z���cmo��,�eM�X�.��D\�>� caI2�'vGnQ�NS�XB�}�r�9Ր��@Ä�֥k�0��s��|��a�=>*��	j�4 �h|(�#�@¤ �DLK^x���+vE�G$qWf��� ���2D��7����hث�����s���2���8�Bm�+�X��Gʽ��&*�z���)��G����þ���5�\�&'�K�%i%#L��o�n棷�ꎤ�3q`����bT%�)��9�h�{6M:���ǦoN��y�,i��� ���=�0k��ԟ���'��G=C��_�<M&QQ�ł^�-b�OX���=�B���#�F�3P�`?n,_U���>�XW?]�#��W+�bK��1�r�9�(6�8�*�S%w/��[}?������.�(h33��8ϯ3!�g��믡�� 4�z�!⊵R�/U~�q6&\�����O��`��C:3d�Ġ���y;�L.��U[�N"�?󖴶1�{��Ċ,��י��pB����t^"a�M�dհ�f��Y��%+H��b�J�U2.��Ȭ�_B�p�7�I�"ü��s���y���� ��,4����8�$3�6X�I�<F�ʹ��z�g	P[TcgJ[�9j6�߹�Tu�Њ�>�d�^��ŚF�#��H�Þ�VH�o��e5/�"�#�F��:�����.ZN��^aU��@$V��㨬I�\L~K�Rp������b�[h-C�#���wV�8Y�uG|`mcC"���������r���!x�FR���fr�+v�ׯ����V��