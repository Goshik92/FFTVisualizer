��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��@<4�*H�	��4����b�7p �S��o\�Q��������T�K�U��
�"g��yJp��Z-���?ꍙ�Q�_5o��ԇw9K5��[a���4�+z𙣁B:��D���H�~a��g��
��YIo���1�.4$�jck+�{_uP�m|8SԱ�n�� ��s[^��]k�2��C�Gc	ćH�͐V	Ry�`�����n��|L}����Z~}�r`�n���f���3�ڝ�g8o3"i�-�tX��z��$��귎�"���k��P۞���mqhQk+=�+x[O��&|
G&��?Pm��r�3 ]j��̪�)mµ�[d���+��&D�C�F�2�!�ޏ�y����χe2���ܪu���?^�`m�fg_P���<��x:� Ɏ_ 7��;)%�(�@_Օ�Oh���A4�`���M�-l=+[Ʃ6�(SA��)C��4��"Z+�c���G�����Z���u�uA����*�dQ<Y���8���6r������&-��!1b�_-�|�z�N|V�Y�����?��|U��2{	�jX�"�L�)N��Z��_����0~j�+F�)�`�ڐ����LM�͓����J�;RT �9h��fON������K��փ�0��[7H2����-6I&o%.RGIʇ���ZH�iU�#͋�V� Z|vg�Q��j_��Æ�'������ܻ�B0���Sq{:P6�e�o#���L{�/������T�8 sDD*z��5�ô��p�/d%���ЀM�7`*b��6�B��]� {E��
e��/O���,A�أ~ou��!��oqH���#�]���܌��	+п_\���r�n��_yHg�zp�d�z㻋��?N��&��ي�����z�຦�&�D��&�2'�/#1U�;�~d��{Pn��)E�*��&��f�c�Q)�R
HO@��UD:�M�<u/o��M5�G��9Ua|�V4�׾�3  ��P;��D'�+��Yң��{�64�y&qK�2��|���k4uF�Ώ�ޚ�n���-��'��_�k�;&�J�iU���^�����g��p󓬾Ҫ��T@���،��=/��J�G"��5��R�a�%�F3W�w�0i�Ӻ��r�$����V��R���<����Q=�`r�ݕG�$M��$:�B*d�G�n��c��6�>�#q��8���x��/l�����PIU1�y��
���a��B^
���'��6.6bc���ؾ���Ց���	�<�4��л��2
�ڏ�8$���������F>�X�4$��yJ|)�5W���4�ў'VBBoTԿH��ZOoyK��a�4���O����tAjG�(�"-"�i}�+xUF)"ں�� ���x:N����_d�>R����.+���{�1{��^��	�]I��gÖ$K�|�]W�b�Ьl�@^1��du-�F6�m͹�ݿ#�Gz�~�Fˤ$���T�r�`���ov��d��}��q[�%]{m�}�<<�9-E8��2����X/X��g�Y����QM2�)��O��o�Aփ%��#�q�f4C������?]D���j�^C=)�?�Cr�Jo���H��������.���=N����g(漪���b�'�P	�fV����1pwI�����yT�"���9  �d{7;_���H_m0�?�U���m픱��o�
6�OC�TSn��V=7�C�;�YB����wʍ.	$�CQ��ӝSض�V��R�'kvqdU}p�{C��d��/��M( �����,���h�����rs�`dvF���B��i��������T�c=�@����8N<�{*<nG$v!�	4��ow�_���9�s������&[�BK0����y%Dr%��ץ�q��D��Ċ+����$�Ue��r���d}:�E T�ceq����W�,���� QA��I�V�҃���`�Zp���,�.���c��$�TȀ[�k�}���DW���������&�p�)�mڕ����[U�ݲ��b�~3��@��?;�Q?� �Bg��D�T�_���d�isKڳ	q؉a����chPA�S9�],\�d��Ț��zT<6�:L����rW�Vm�	q�o�̺v(#�1��>!�Ƚz�C��ʉ�h��0��ԙO��
a>�$�`���doK2���M��Cl]��}0�~ ���su�e��9�R���HmY��6]�:�ļ����U�e"���?,�d䅻���/�r�}NP2`:o}�B<��ݓ�^���䒚���͊�-��z\�6=����p��!)�����0�AŴ��/Gߗt��6�RϨ|CO ��H#�AP?�����E�J�b����س�܃#º�����, GXJ�ϱ��"���x��68I���,����5��rW/����KF��h�F�h�qn��E� �>��🞔Q��E�K�n���� m/��Ϻ���/cri:�̤��X�=֠v�y����������B���[���dyOw���/ ���� ��Фv����;a�"T�&�M��
'�`����xA�n��%�U��V�-�"�'��^�G"J��
j*ߣ�(EuR��K��j-[��u�{f����I,0�^1ߜ=�$��f����c	+���̋��[��|V���
�af���u�0��DN��<���X ��{��P����>��1�x��ݾW��yHP����¢v�ۥ���q���N�pm�rnȠ�~%<�owu|���ȿ��k���F��Ad�AHC��=�1lR��eG#϶t��ԙ��O\�e��Z�����P}�l���4uQś=W*���Ë��jZ�h�5�tF'@S��7�;h�+� �o%�@i ��GF���Eb�l��y����VEr����koᢞ��e�	 rjH�����8aW=$��r��n��̞�s87��R=u^�CV1��#xeK��*|&�=�`s-���"Qs(h�Nh+�Ԁ�w�$��L`��¢� -ǿ*��v��j�Y������;�:$���a�T�1��ϫ�7>�27��Q�K�W��"�����{��������*�
�����v�s�1)�jȌG��%�@Z|��m���i�٤� �
~`dD �$�]霎���U�N�:Ոq<��E�uѨ�Hm�e��*;e�����5���w븮�{���n�ӲI06� <�_�p'웃�OPS�ĚX��7������5�i��~}��x���u}���OU�Ƴ���T�yx��{z��,Zi���]J��6��|C��9����"-���>c��T������Yނ#�+P7���:1E�,n�*��3���񔂤�w;&�BS%Ͻld�<�}�`5���ap�b�4<�us��'�����>���Jw.�A'���f����xC�G�[�1�BX�!��S�]=��~>�n�3�2M�v�q�T���ο���4�4�<4��IH�E2�TD��`�	_�c���R�3x��#c:x���K|wO����{���L;���Kv��5���c��v��x P��R�ؑ�6�8	�ȫ�@pz�r
�U�ӒjQ"�:���"�ȗv��qB�\����y0Œ9��G�Kc�����\k�*V�N�!��#��YJ��ލ�e��A,�:����貟= $��o�y���0�a`1p{ �6a��K�t#{6̏�FqJں)p���O�m"vK���{(���K�>�ޔ������=��A�q�`��\aWi4w���l�k0�\����0����yC"�������=Գ�׫�w �R��B�x�n���� ����!�7n�y���h���%����v�dFVߗ*�'3�&L�Ɓ�EY�;v� 5��|
�����{�����<���$�=p�`@۴�R�E�b씖Ɣ
|m��(�0�k(�Ker��^��#�r��������*a��F��=�������c��䔡#��lgK�{�Ő�B*���햣���t���2GHS1���׀<��7L��jf:�m\���Y�hIgK�~<O$�x�����N���!��J�%���"����l���:ER��f	{��}�~�M"�^�� 8��[^�l:�(	Z�Nd���
��3�OU{��ᔙP�zR�o���bbh�(�rF�ٿ3�PuM��$fh�-�ϯ�Ӹ2\���f��C4��ʲ�����s\�ᗓ?Y�b2����d�l���Q\��򇌴�����{GM��T
u����z �..���W��}�͑k�X>P��8]���3��G�� o�3�Ľ���� &�;�nʗ�6e�?���MGY��/��MFo�1��{@6�32��Ňy�7����C��Z�r�֌�4���6K�����-;���X�'^R���Q�ϝ!+G��_܄B��1S���c�[_��j���۸������G�?�~�J����
w�	eU���%�E�S0��ػbW�k�aNS�;H9p��
�!'a�K�r�]��JىQ���d�S��k~���W	��<����6dhq�ܗ�nZ?ؤ%��'�Y�}8z3뿾�0��o����ue��'�]Q��%穦��'�YYԟ��Ф���������:�5	`P�֦S4��D�/��<`��do�:�l�^M��q�g��������f{p4��g"1��@W=W�T��L��8��	L*���>Z\�?�4 qU|�jZRs ���6�Dv�������e��>���=]��
���-ñǥ�,�,�F}hc��L]܉Uw{xEmv������Zfʁ��b�#C:��l�w����f+��Y�8ntt8�2r4u�te���",SJ��6��=�apIQ��xO0�]y�_����3�����p��>�;��C��<��R{玮f��9B����O�B�ꀭT]��S����]}�ќ`���B����y���K)��f���[��`@��&�9le�)�팸}���g����$-Ͼ�^B�-�	 *55�1�r�_���u��?C%�J&�pM��e���K�������m1���{�&�|�#	�R�s�0{���), ��������wϫ����$��d)�\�!�ȋ���]>��v8���W�| �jrm�6�x�� w��7���$C���b!��2�-��0�#?�}o�2)V!��vE��������Ӎ3^���{�1&h_V4�06�x�� c�ֹܦRO��~u��L�|�P�4޵�(?\�8�Y��/���rg�.	;�i���Tl�����Z�G��Q��4��0ϰ*����.k1�ǏoI��8[�%���d��k:����)���B:gݴ�r"�L�䬆��.�?a?f��Z���PR��}m�-Cl$�sn�볤-ح���J��^�da]�=п�f�~y4�C��?Di&�r�~̏E6֖ma�%��
�"�'�B� �����
��"�㓲c�\c��s狂.��_�X@�vf��m@��ٱ��:�dV
��#�V{�>��F�E�oo�������|m�@�8���Q}�&2/e��Ԡ�p)x��$0�TF�BM"ԵQ+n�2���������)�O���Iۏ�u�Ū!".2��H��I��)�Y��mlT�6�E��Oc��7|��%�N��z��9�>*��WjP�G60��ޢ����0��EL"�� ��?z{
sv`Ѹ����)���:ſ���D�bB��K�������B�*cY��!�3��9P]6�|��%b�:�2+Bd��C��F��'�}�j����žSu;���(	.���w��e�b��xL�����B��Q�&�9K��� �@�HG��<�hd؃���]M��TƢU�1{�W��I�xL~��_��t�f՛����8� �������z=�2
y�'\ �:5U��M�����~ץ�����0�r?��b�����9�u��7�h�ݢ����}jc��'���D!�Ɋ�͚�h���!�Rj��1��@|�q�VѼ ���b�c<y��B�qå����*�Gˍ}Aq=�A�yʚQh�!\�@���Ӹ{Ĺ(�ǌQ�
�o�K�z�{e�&�<�UC�s���c(&�W0~QI��M��^> ��d0����2�W�!��)����wF�H�4Us��v�Xk	�勷P�u�
ȿ���*�<r���I�dZr׭���u�p���ާ.�;Q��yuu"O�������0�-�@�N����R��;���Rq���us(>���������(�-��n2x�*ف�)C�'1�M�P]ϡ��1G5,�Mj�N�������tP��y�`!�Ĺ)�b�M�{��R��� �a����(e��z$�:���p��֠%���M{�;{!����g�K�/�����}X���yxs��Ƚ�ek�1�? M��?�`��$4,��|v��+�̱NU�9��X
�@����͂n��;�D�h*Ĳp��~R�L�߱��.��)��~�g$�䝛�~��fI�7����^$Xa-�I��NO��&��<2(E�hV�:^�ڰ����Cg4V�thv7�tn܀�}���]aM���ZX)�Z��ci#�<3��u���t�b]������;]�<<�2�R[{'S"~����z����"F$�9�TU.޲]�ȍ�� 0k,`a6���0A��'��f4?�b��j�;d �xq�x�e�a���� ���$6Fط]�㐮�Q=]�x�=I��Pn��G��Q�F��a����N��bh 7i��BP��Y�o�s/`p�.�������Jw��F+U�n������d.lԘ	���p�9[!v0�c�4`�����Se�%�ڻ܉�ĘI����'RiG�����T�r��'x�Ղ���?gs�u�x
��7*�R��,��[
]T^vE����|d �,��(ٖu=�*Z3�J{� �n{S���z+�a���N�k,�+��ƷuE(]�$����ma��h���i�=#�Q���ܛ#<d�7��'4�&W�,�v�%f+�k�#`����\�������@�-�	�M�w9�0���G�������w��9c��k�U�-fxҲ��׺M�!��I��`ti���V��ܕTfV�?L�����Y�Y/�P��H �����Q6(�d
�ŵ��ri���[�Z��ll�w�5�9���B=�K�c��͏x��
��.'�rn������<o6"`~���F��j����A�-.�:q�q�qkCd2�*R6��ԇ8�m+W#�vx�U�E�ʛ��������K��A�K3�G]�,m��9���B�Y`/�G�)rf(0?p1�Ӕ,m� *ւ�+'y�
> �$���sfݻ�$(�?�Fjf z8G�I��g=PSP�':������="Y!��d�~=xT�p�L6i�qFMDH�!K(��*�b�fեR�^�cۺt w��Xe\M�q�]��Z%�㫋47|&h��\+����e+��y���c�W$�"��4���j��l��P����D���X���(�2�@ֺ�{!�V��5�Cs��P=�~l��JtopS�E{�3u��M�������a��b#�I�`�J�'j%u��.�e?y��4���*;��/���f�+��쭞���P?VQ�E����C�g�4��{���,�t�ܱ�����q����cu;�<@���ËB�kw(�Q)9\z�Y2xo.#��7�6��L���K�(2f���*�@�?�� T9�y^�_i@A뿢�t�����6��$ٵ�-ǿǛ�Aպ��� �,�;��,׺�U����8�O�D�Q��n��h�? ��	+p��&��(ڡ9�6)���1�#�݌��Q��{ 2+�Ý�S��g���D�?7�!i�H6Ǹ�����=H��s�S���4R��y+MZ�4�V�)B�u�ݐY���[@�����Ӛ-w���l�cˁ���F���L�W�е�F2�i�{Ș�GY�ͬ N�L���!Pp��&�C��`
�'�˧�[���gʬ����8���Jf��~�M�7~R��Dyk�(E{P�S` ��dL��ɾ��S�2�u��P"[g���݋���A�NX�iZ0��Do��$Df|.�caY}D=g��{{	���}���NIF�i�3,V�"$�3�����lK%n)��z4�W&Y<u�*�i����_�<ƿO���yS����$�H@��j�gXk����2�+�n��|��������!m��G�mg�W��%��T��x��pݲE��z��WQ�fׁHpe��͏my^�E���C�`gs�!>�
��^Jl�R7=|]�(��*��4deix�-��d��L,�͍��fFq�OB!ðsH2�W,� }?���=�o���'�O//�=w�	����́<Y%�.>?� ��Yo�ow�YqX0)p(�if�BO	���o� C`���qo��s�y�q�0-�ˢ���f��A?����ƥ'�FRf��ă��S�P�&�sӴ���@���#��:T(jh���t橜Y�����41o��&�RDD\r���m4���Ԟ/Q�["E}lZ����c�l�Z=����n��ɲP�<���l�i2��ÿ��z&3�7ɽ[�3�b��#�dO�|[R����Z<i���JbRSV�R9�ap�^��_d|G(�Ҳ��跱TJ�������$��|D����Qxjc*e���d�xTkP48(��� kZ]؇�lM	���Ax���~��JMIF��xD�:��&?��ćf+�I����#�Z�Kq��d�8)_ϱ1P��.E+m�i��6�b����QD����l���+7�NX�#�s-HE)�ɜ(�3:3���H�����^mv>{���;&���{+*	~ءuHDt�EAf�"�T�ר��-[�m�.�����4�����SK�Ӛ�wV#[�gr�5o/Srx�Ћt^�'|� ���U��ƹ4o�%�^�z_�[;,ڞ����8 ��v�^���Q�O�I=��]8�|�L��Q���v"d�_��u�a` %�Jd�&��c����i{o���I��7�d:�\ @$��_o}�q�8��Ѡhq&�s�.äM/~�^�~�yH���Nu��$���>͝����s�_ˎ��ɛ�o��ںkF"yH��!v�U��F{yf�::��hV^xF���gjxq������+Ȥ*�Ԭ�hm������m�׾LS.�hX�V���m5(��Wl�p�G�x�yw
�{��	����0�^�``�=�I��������MȆ�d��X�w��;�P�I9O!'�f=!��.z�H���k,�����&v�0�������S_�O�,i��,*�m/+�Wь���Mīt�H�\�&h&����!��'#ڱ�~���-*����b
d�*��0v{W�ģv J�2���aXȝ�2�:z3���ms�J�t���J.Qs�,a� a�����GmsG5/�{��3��Y�3�u��9p��l@tp�:�Nn��3�6��Z�6�@��>2o�J�^ѨU���aV��r�93���c��f�bR�����Z�A{�6���*��; ���B���$��g�Sm�]���R$
V�ǡ1�D�2���K�A{��UW��.݀��j�Z�j$|�e8�n�z������]�Y�ہa�c����l�I<�[l6]��T={<f��)�B�\�K�.��a��jp��z!�Hvt���\,?�ѩ%��y������itK`T�������Y<�7 �z*,�@�����q��0�ɚ;{cs���`��a��Z�}�lK�:A1���x�,ڇU>@!�-�qec�H��_��tO��������d��7��u*'!��~�S��V�� ����tO�R��v��Mo����x��e$�:���� qz��x�������� ���T以P����o���/+�1��?*���D&`om��:X�h�\��HҴ�:VY���
TO�;k��7�bf�I�8O��@�e<1����6��^����B�>ε���:���r`��"�kE�<K�4�����~����(�p<Nn��B��龲0us~G���\����Um
�&�)��c�ʮ�k�9�T!o߲���!��6�Qh�?��|"2R��bܧ�WP�/lIׇx���+%:�<��N4�u��>CȲ_>�a`�ٷ���z"AQ��������k�/`B 9L�|s����ʍ���sň�����V�`�mJ��a�VZڤs~:x�M��#��"�j���o�U�[n�Ou��1Ģ�0;����6"���tqͰvu�'NC�k�con�D{P��r�[W~��b���QC����lO�@�{)2��K[�D��2$�C�	���Oʀ�Q�݄�Γ��p��#��x>I��jh�PT�ڠ+K��C��G����%s��Yސܫ"��������[�C�`��r=��ns�q��"s�����q�I���f��2(���K�R0[6��;M����������J=@Z�O���Pѝ:�k���zGLQ������������� WrbZ���P�츐x ��<�7�3�*Mw5Qwj'�z�D<� �c���9%�(��8l��}�����?ȑɇi���t�~uJ���^6>�|��j�:��IqԃFfa7�@��{�\߯�d�kɐ\ÿϙ����D9c��/KD��T̵U�(�;T	��s�t�_���R����J4�Xq?-���%I���l� �.2V���������!$��q�ʲ�;��3��m�?M�@�u�%��D�)���<�:�%���c��n�n>*�5߹�_�4�dK�J��X^������kŲ�>Y*��+���Mҧ'�aa���8�I��ܑ���z����яbϭvDLBu��hF�-�cKޥ�# ����sn2�"�Ňyo1����{���hK��v�%Ƶ�	�Nxƕ�]te݆鿠����fhu��z�
��璏PX� �,>�%����a�d���c:>����yV�\������0�.�{;�b�c:���,��\f���t�T���"6�9�2���::ܡ�b�!�� D�Q0���!g��wZh��zebˉ���m@og3	�~+�)K!|���zUC��:U
q���Z�X���&�T)T�Fp�����_7տl�z��p��'�/��`�_��L���+�6�VQ��?�to��FPD<F_�i�B/�?FfS��J�\͇9�%�U��wMV�x�.˘/�ha,>H70�%Ϻ��}t���=L�����GXm<H�H�8c��y?2'�N�L��/.P�͘ʜ��8�O_ ��ȍ��
�5�/�l}�/EӺi�M,�4���Ow�h��sܱI��S�y��|��l��[ՠ���w��F�MFǅ�n~A�9O����3���Ф&Ya��-$�N*\�H`�	»������`14ٮF�[��o�楙��Ƭ������2c;�'�*����	z>l����)5��4�K6��!%5t7U�x<��F>�v 6K��QA�>~'�g�wH1���^��7��=�B�� �7�N����'�M���>�4�r=��΁�Ny�1z��\�f�Q�^�Ms9�=Ie^B���(Y��h�X'H�w���'*Y�+6�j$G�#Jr.�Ʒե3��{5��}�Q^#>�ٴQ"�G��*q�}�N�� +��]	���Kg&l�W	�H4���[頟;�ê֪o����:��Xm�W��
����1���~�^M<T�v�W�7�#�%���3���X�2xu6���W�N0��Ę��I�T�_�f�B@��%�J�7'��*:���ѕ�<��^.^Ǚ����C�� ،9i�v��o�+�,dd\�:����Lv8~�w�'u�UK��CH9��2hX����-��W@�7�Pǵ�%mSA�	�g�7]���{׃/��/�5��zB\���{������ށ��Z�Ig��Ê`�)帒+�E�x�������"Ջ���i�����8 �.bGw�L����s�Ԍ[����᧞�y;�����Ϩ+C/�v�Nޢ��U1��`�6`�UyD����z�C��(=�`\V�Qi��a�/Ȣ0��XPI��������K�DT�Qa�˿g��a�%Dɚ)��$>\u�^�Z��#�J��J����Y�SE�M�c�����a�ΣV�=/�N��{�Hr&����U��]Ě����Gn���@5�k����JO�qٿ���K�ys�|;�_+�)�q[r�[���0+4'�n��,�Fh	�6�.4/�=t�0P����'��2`�X���5��G��HL����O���Ī��@�렗Ӟ��{�Z�w!�8c���\�y�o<p"
i���&-fjF�7�Y)�D|�K
Bv�t�Z:� ��e��W-�<p�˓���=+�-��&���/������a����ɰ3V���M�\i=Ϣ�[��frR����F���o�� Ϯ��"�`���۶�LoP�ā��������n��
��O�鮝::!�Y!��WR����cI���������S}~
Ξ/h7-m�x����eG���Z�I17�X���#��`���-Ʈ��K�h�R����t�	q �;�/A�fG�É&�X�Ѥh��X3�uוj)¼��[SSfc@ٳG� 9K�>g� �Դ:x�E�W	�K��Q��_�d�vĢu���K��dy��:һ���X�Y�2f�.���������S�����ҳ��MER��{�5
�)=	<� �����t�U�e<Z/F��~T�}�}vX���z��3%���=�ɢMIkɼs鈫�l�,�uk���̜H������4�ta���V�Q��၅�f0�//�c9���H�>&t�^�����ˌ{ta��_B�-��T��B�y��征=�[ч!Oaۅ���>����p���k�EJ<o�vn,����D��$#���h�v���^����`�!����R����U�zP�o�T9|�;) ��
.�8\�PB_م�U�g��-s	����D9���W�HL��Q�k��+3A~��ư*[&�'�/� y�m���3��V��(]�����;.E��9&HqL��lP~�GF`�]c�:)(~L#p��䎡9�O�N��`Y�ی�N������'��Bb+,��D-IY�ߔvo�K�:�@N@tɦ��t�]w�-K�fU��H���H]t#z�x)	�
Q>����3оlUX�آ���&�*q��\9ZstW%Yᜉ��0�jmNJ�eJ$�M/P�
+�<�#.�I���ʠ�ƨn�����J}{��Ž�\�D@����C̃�E��D�\o$�|q��4ۚ���b�8�U#��0:���v�Ed����7<w8!A�e�怜L~ ��J�Z�/���hr�l81���I�ᡩ�XB��:R��Y�oT闰N��K�2B��|;XI�L�,*B�BB~]�Q�?�NbvT��P��2ٝ�����{�N�j_ΉD�,�!CA�!j�?�@�ǲ���L�	���T��+�=n�"��@�񣁷���Z�ȉ�\և^fz~��4175���Ezl��-/�Z�N�gP$��cB���)b�-} 9a�N?ږ=��`DA�A��D�@?���D��g�q�:7�ԀI+͡��T�O15Z߿	l���_������O1����+�rPv���.�ܓ�x��G�U�ﬂo���a��G�<e?Wyi�s�h�8�+
�et���hmԳ���X*���Va��=���]f��A���B����+�l_I�E��,�](���o�g�I�N ��f�lClu�,�M
%��J�[���:�h1��R�ל*�I@w��.0<wO�����jo������C~��$|��t���$qK�QE�CPqC�6Lj��E�,�>�[�������;��W�9�.�ɭ��L����}q �i��tNE��s�x�#5��,�K��}�c���m���z�G�|j�g���l����n���C����
/�b2�z���Cc�j��t�0���K(�l���ťEW>�)s����5r��&���!�ȓ_�a5P���R����r��XI:�o�Ub/7U�i(�s�����r�j�u/�����6���f��5���,C�EDՑ۩ևz���hi������m��\�!UT��}H��R�����y�k5'�9�����n�����9�!�P1ǲ���z��>UYA,_mF�y�&�x�z���(/�\g-����f�hc{���'n��g'���~��퉪1����I�qa��������P��������=
ߑ�nA���.qpwsUضd�p����egȕ�1�����w��sD�>��o6E�Ps����掅D�&9d�ȭ֘��l������5���R?�4�+x9��]@DXj�!��k�^�J_O]�����U�G��&mU֖��D�b�t3LG2�O�;&��Q�0/B3�����ٜ��h*�ɯ;��P�bp
ח*���zV�����8�x\��9J��tԲ <�*�*�$^3m�k�����`H��!	���Ea���z�1 y/ŧ�8Sݛ����^r��GM��M�J�0o����[��7���w{��7���K��,M�8����R�yv�atg��J`NbG��b�����Pk*CZ����,��� J�I���$����w��c,���c�/jQy��s5���!��*ptۏ0�|"Ӛ+'�B�aG��]{���tjwٛ<��8��f'SL���&�wn
7���C!�,P�J�~�{(p:���0Z�����(n6�X�!G/����E:/#����+	���eG�rz���M('y=��'o~,.�|���齅5Q�˓�a�(�Cc�_��v�F��;oH�)�W�z��B�5]�O����aԤ��ΨyD��N�s�K'-�o�
��0-c-�Îؼ���5B>.�2�:�Y�2N��ŷ�A3qg~	!2�3�h�:�$�&s��zkӿ���"�D�`Bz��$�L�ڶ����=��d�V�n�J���L��Kb��2Ѭ��T��/���UL<SʽX�����Ab�y�ɨm1le��S]�$��&�ZW�7����V���;�%�:E�Ȫ曦?����;��y�_�Ì|\�ȊI��mBk9[��.�� �F9E�RR�~ˉ�E�T�vCbm�$g�PjMz�.�ZJ�"�^��1fg ��l�������VI�Z����P9�9�|��.e�5���a�y�|����l��e1Inqm��I��1<� �Fv��ΖY�b�-`��e&���cJ&��[tǧ �=�6$	b�����|/h�Rr��3U.A��y.��p�)�����V����T���( <��� ޅ-�^Y���24o��F���>�(�?<�Ũvk؎��:�Qb�Vn����	!��җ������t��8Vng�3}T��j�@G�ऻCx�>Z�s��V�{�L�(I��#�M�ʓ���N۷H^��q��BYk4�;�y���pi�k�H�9;A�5 �cz h��h����h>�S���	��� �l�I�����I�z�i|Uu��.����FX?��R�\(�5��Gr�g���7��{���@A0��E��JÇ�F���&J��W� *��	���2��yE���6F�g����z�!`������p���E��Y��1�Y����D��G\����]1�ao��"T4��ocZ"���)��%���������� �{U2�WH�;.�&R���:�,���b�;�sT��Ge��7�@�"<�8aE�T���7�`��I��/S�_��=�h�&aY����tח�I��>�b�ޤ^��O�����X,��5��9�Q�� ~�R\ß�x"���P��&"^:#��w�	�/#��]��@4#n��>�MC�R�m�<��:H�T��^��2�$�k�X.�|���G<Z�*�\h���i�ΛО)���(ܩ�@q�h�FY�q"��1b�*�Y}A��ɋ�p��I�R�� �����0���C࿽��$���ZRh�<�ǆE�5�y��@'�P��
Bj����/`pn���{	���O⯄3#��Sks{~	M/�M8n���:����'x�N�G��21���PӪH3���3Tm�)%����s���PL_w�{��������2�k�#?���A���ɖCQ�L��B��hAwn�#/'F�J�G��o;.5\ySАy�V��恽�+ჟ^�|1ф�;!l����(5��2�#��
9!oAUܬ�9{C����N�<�3	[������v'����_Sﲕ�$%r���_��b��d�u;��AKQbWDu��B �t0 Ū��<,��n��a߰���׽v�
�Oxb���kCf!�����X�t�����fLzl��v Y,���V��N��#�>u�عG4T|`x�	K��l��vWu���fs��BWk��y�<�G,+��i�P�xG≻��y��Jq�%l7��`���B����;S��r��-��t;0� T*K��4��3�3(�lc>w��X�&��}�~;�#X+�u�L�N�I�d���$/a:9���'�s��	V�yZ�x��Jo���/$u���
������|��p������ 
�*a�H0���w�r��伳�j���hąv J-��+@=-����r�,<_�� �����g��/����(l�"�=H��9���h�=N���Mq-�Z�Q{O���u�G���׭M,n�o�rߟ2A�[�{�G6�L] ��SRl ���?{X�tTXP�pϧ�VZ��08w�B�ʹ-�������ĖOى�^�3h�H�)1��K&P�4��.T�@����_�l:��q��d'ɻ�|���b�V��,�*���+3� ,�M| �un3ɐE��B�v&Q�?v��ښ%�#�̬ډZ�r<#�>�YpC��O!��Am|��R^H���}�_N�����'f�t��Sh���$�v`eb��2*�3Ĩ�� ~Z8"ZQC��r�0!����L��o��;�w��J�)�1Z�����x��X�`�Ebl&�Р�wzh�7��,�#+��r��K�U:w���=���<D==��`W]���-�����?��i�׌ZR�4M�Fy:�e�J��a��E0|��i�H�-�)��͌���@�v)k�.AQ�gS9�Hؼc�����!��K�i��G1Y�����n�(h�,��|�Ƹ�ac ��F�nO��=Y* �	8�waŭ�	贒?�	hU�ڷ����*�Fne�	r���h��~s}KWk���Ҙ��Gw&W��8o�f�Z�A�L.N��n�A1����\)����Ȅ�8�<7�&P�p��D�	��Pfx����J�yS#�����PvnFG#oܶQ]�ʃ��˝�3�_.�F�J���HY�����ްgq�|�;�����o�#��\���n��nb��Z}-d��X��L����ɠ��FЈ&�'˩ۗ#��
X������8�4��p�_����c�a��F	� Said�9���W-i��M�-K�>1C�ae:AnV#�&��/rBq�B�h����h�,��e�e$S 6X��������=�g
�����<�yO��쵙�R芬.T�CĤ��Zy�4za�h4{*K���_�U�x��0�h��c�G*�Q�ώ��+>N�|���>�t�j�/�B����G��ľM��C�r�Q�f������1��xK��c��`�Gd���q� "$m�Ҳ�.T���q��܎ⱎh�l5�ߏ����0(f�mZ��o���37����s�r#�N���˼�Ҋ+��w��T�R��Z�����k��Lՙby��Ql�"usn�0����)��F���leXxGָ�� �mM�f���V����͢���lSaGP�g_~A&c vX�ܯY���`��4@���'���C�^+(������!�1)�S�B0l��ܨ]��A͍��'dG	�踈��ue���nj�?��zN#�1r/ �` G���TH�h/����D�����ZF�U��u���>JF-y*~!��X��8��}�b����6�^&���84���O�^��IQ<��o%zֶ���T3�l������z4B^`�"�.E��|�:z6. ��dӑ`y��ja�4}_��)O�G)[:�oΈ5���W"���{���U��H����|@��A��e������h��m��K[�Q���Iս�A;�1�O��r�0�ܗI�B�>�^\%7W3�U�\�G�����T�.��ļ�2�ׇ¢2�fe<��"��)BCތ������k�ķ{7��E$��x��l�m�N�m	�B�+��п#�F�9��7�^��/�O�ú�$�v�`b���d2�Ä� �t���[�B�����x�SSg�9݃�ϟ'�Є����}�]�-��I�mѝ�Ƶ�:&��S��=,�ݳ�؏��1��o�_�Wސ#�P�o���̞�\�+�as�L�6o�%�`�>//�8�9���U�U��S*�8��6h�i��/�5t-��n�M�lq��'"�T&�AjS�:{DY>ݘ�ڇ�Q�t]��>
�X��7(��Xu��%��v,�Vo�0�c�W���5�r��A�u�k@�lP��)-4����]G��߀��X�S�H�����j�d߁����ut�6��oH��7������J�pO��ʛ���^z�d$2&scM��4���toG��s��"T4��T &Ɋ�T������Բ���09Tx�����Qu[!̔���s<U�ѣ���@�5���ڥ�R�b�bʘ<]b�0��u�Ԇ�\#��H����8����&��<��+�*�*���ф�E��͕�#�A[P��!����î
�[^Y�A��+�b*�g�V&��h�+d��b�l���O��eWf_�Eh��Ȕ�Wd����I��u|�Y��0��ڽ�����g�`�]��g%��U"��{�$xUK����iS�m׭����Eec��<���[�|���Q�hr9�A������w�	)�26H`*�{�>����1��O����͹h�I$�P��D_�_h�ʤ�'l��D>��|E5lF�	6��9���fr:�$�|�2�������3A&ks�za��"���K5l��Y�+nrׇ��g���QW�y���?Ǐ�8Y�0�R[7u�VBxb$!U#6	'���zGG5�+v=}��(���������^�S�R;�#�v��I��=��Q���4M�0����� ��������>�����R�6��N�Q*]�j;UF�2�oS���z�>;φRYu��p�w�5E�ߝ��n~�<8%�=i�y���:�v�?D����Ё޷��?F��"��-�LX"���gq���ŨAX$��VH#��y�z���7��o��$�L�A�a�2�:�'�E=f���YS�Ү���$��Y��iZ�Ew���uqm4�9t����:��}�k6�X�&���Ч����n�B�\94SlD)�Q
oo+;�Y��� �H���5�v��'Kt�D�V3� �~�k�y��|~˱��3/؇V(`}d�0�[��S����=ӈ�����!0���,���5`����Z�3:�v���rJXͺ0��Ͻ�[��|�~թ��5����+��6rK\!�g�����*�yz�]���~\�:�J�f���v4��p�.�\B  ;?TK�udK+���j��E�O���~B��zE�D��u :��u�α5(���-��Ȼ�3JZ�S&7Q��
Li݅�����9��O�U���ڪ�c� ��}�mwrp�s�"���rFT�&�c��������J
�|sߟ�(�����4�IuqZ:W���NO#�V��G)�b�Cq|PS�^Jv�C�,��f��L�`�$z.�w*��~�	6'��</ׂMj	3>��H���
�j��}��@?����.��tp��>p* s<R\�n{�Xew�7{﶑�j�yG�"�Z�\iA f�')&Q��C�y�CW���ۥXy�)�Rw}���?h�Mhq�U�08	$puy��k؅���tbU��o�B�o���@�N�]j��}��ΐE%mG��uȣLĝ�-Jۿ�ۂ��a]7��%B�/1Q�)S��:;Wa�*�<��Gw�+�2�Q�d�x�p:Y=-�0�gjs��'O���)��:Y��5����{2F�G&���{�)�$�1��Q�fyybkFnm����&V�˱u���I���n�|I�+a4C(-���^0(rɲ�T;��1zgf̸�8�J�T�����IO���oS�)��>J(N�����w��@%���/Z�hb���8I���,��0k(�e�;�"�2�t�df�}�[R�3�����M�-iк&��I�P��{�`�/�,\^�p���/"�:��S�{�=7�nu�61I���v��T�{eo���&K�6���[��E��Iܜ���)-�R���A���_�<��Yw϶1���3e�����ӫ��Q��W���-z��=n�G�.�u�	Jӯc���+T� �פ|��dI���e�EA)��qT4]�C�P5���6PTm%~�v��uȅ�7p�7Ku7��]h^�8����mR�s�2G���v�<���m�]�;{�m�o����N�C:�oT�nܸd�z*}�5~ Sh�����(ޜ�~��O�P�³��/��l��Id�
<�܇�au�/�-ị�/�3;��g�����X���!8��񢘥>�X�oJ%���+�J�� ���ɕ��"�֦�6_25�YΨ��C���b+;r����d����^�c`㥁��~S+d�0bf�¹�_�R��c�n�Ph"�{R��L�|�[OsJԠ�[��m�bj�Ń�s�V��\�e˫&�LX�2W�\�}�<Ť)
� 5�9�wF�4��mw$M1�<�֊�Q3�E[����b�:�."�Ԉj��ҭ�U��OT����������8�4���xG� �1���6ڞ�0l0�rO�pr<aLc��%Wփ�9g~Z�J:��c���e汎��c�l����i��_=k�g=G?0J-.�������-�
Þ��5�p$C�*�����c{ҧ�z_=U�'��|�x��-�~�y�<g&|�F�V?&�e��P�a�]���-�Ocɏ�qʦ��lzv����Utg7J�X+ v��<��F%r��/�n������&��f,w��d^�+K�]��m[���u���(��ҖyEӷ�x���=�̹�P��k��#�.�!�Ů�^��)��y�i�\�8�"I�Ax��⑞����F�����㊩TҦhR7��o����R���S���J�����P�w� yW>�}+(:ɴD0�6��}���PK�Y����l��D2k?��%֝�K�����}��̨��8Q�
w��H��?�{%?�{� ����+=����	M���׼6�՜;=��+-���@z�Y��2w�R��LcTB�H���5��̫5��%3�k�w��WM�c��;�Q�	�@��;A�N�I�g�=��09��c�VOK#U��d��ׂ���ѓ�>D�[6��~px�N�/cJ�����Lg�#7��[e<~��'�A�Euq#ui��xq��{6D���7��t�'���|��f�<�j�?-`�"3; ��ԯ�]h�cmH}�/���1��h|�"��sP�G�Œ2�Ӗ�[�CLAI��؞�d hjee�ǥGr2�$��1���MV`�-�L�t�}O��4�������������te�����e�~@n��6�����i܋�i��*�!a�{�0�7�M�<��#��ٱ^����x���m��f[����%���Y�0���oS^n%��$);ڕ����r}|���rb�\�@�C�TT6��%s�}��ta2T�3�Մ
�����,na")�1�8��5��lC��<��}' ���}�.�^viB�{NfC
/�Og�ŕX|�_;�b]\ǣ����&���>�Uv�>��6�����h�,�5+˹�E�e3����e�u9��Fzڪo��=hW�X�TL���ᐂ���&\P~@�8� 	�~�K�y|~�H*�f��A4��H2�����ye�~��۫�ϳ���0�K[f��ª	Ғ��K�e���iB��t4����.��h��U�o�R 9��yb,�����ɿ��"�Aۂ�d�9E>	^��i��
 ��� �qP����~e�R����u�cr���x�Y�WVlB$�vo�gj=Drj�A�#s�����S��s0������TrzˢQ��z0xC+4N��R��E��)G����۰�|F�ݠV�ԍuEw�����O[���!�d�
 d��z�r��r�E>&(;2Wɇʹ��K�������i� R|k�*�s�Ov����6FW;iꘔF�J'�3���~*��#��`�&��/�>�G��K�����_(*���Am��Tw���.P>;���G�W�v��2kY�u�6�cC�j��e9��x<>(cnC�M;�9t���S	[J�j*b/�	
�M�~ʪ=Z�N���c���1���p"�s8J����$�D�-|����rV���
���wF�Xi~0��=C�˽t�o�aM%�I�uw
x���Y�T����Q���98�=E��}�Y��*=leH�;����i��u�x�o?	�mJ|�Y�2%S_@ b������6�,��w����e:��L�%Q�����k,��q��������Ԗ�)%;
��9��_�/�P9i�Ew٣^�Z���������}�T���{�z����C�.%~��V�2�OD�7���<���6k,$��x�5�	���]���¯� ��-�I�],,�J��^�9�8Ad�-b\�� 4�-|#�~��6��q_E1�սnঃ@ea�,�W0s���u�/L��p+5�y�q�2�8ϑ�*��bG R�y2S�_�T�-09�Q��n�ǅ��M��H+������Sw�ag.u���_��A��\�&RrJO�=��q-�TN��a��Y��ӎ�Ar7��W��ȋ��R�@m�H����pYS�훽��R�\�%/%�a���ް��fJF��1�+f���Xe����Y�.���K��R��f*f/���۬x���V�&5��-�60�%���vZ�;�K���m9�ǖ��D�*�2I� ��(v܏�؈W�ª�`��	=T5)����g��8��1P8Q�u傘����L�.5�6��$����={����[�"5���g>�G�؊�.��l�g��0���:6��N���)��,��9$5�EyD$г���h|������9�?C����4J�`���2wr��g���r���"nOp��#8/��ϡ����oc�TvBmZݡ��+0��s�e�v�u#:�qi�,��Z���u����uTA�ӂ�!�\]�-�9��Z�+C��ϑ��Ǹx���fW��m�,&Q��PޢJ�B?�6�?�A`�Mw�|<BÍ�+H������I:���k�U4�]Q����C��W��Z���s�[,�B�[mz��Z�K=���"��>��0�l??=	I$��h	n��s(���&���ħN�'���~y�B�a1���rݜ��}�0��B�@��Eu����2K�o;��ç�k=di�j\c枀b"a����b�wܒx0r_K �v�[H�1���]^��	"S�.I`���	s���|��K	?=h�1,�M�F�6��&c���&�����a�{�5�|�íTAp�%��P^����)��.�651C��P����h^h.���c��{�=<��'#��1 xO��i���y�Z�&�Jg*S�V���K�I�q�,�� ���;�5��o�Pb|>XE��ct�[̰Ƚ����!�N��Ac^��V=�x��/�+뫙Olg�����h�x��U�d���h�:��t���<�E�����1N�]�~돧%����Wa�17�-5��i
��˝J��ϑW��!&�[8a#`��0�>�~RT�Q���u�莄,�{�s�p��b
��e�`j��������ĝ&��OFP���qh�X�WXT��11f����h��w��+�'v�-�/�&Hc3��ڐ��R���|M٥\��`��7��%{�ܠa�"	KLB�#7%�<L��<l��/؜�t/O���VW�o�l8��z��۩���a�Uyٽ��.Զn��-CL����F uà�Sj�MgvV�I�}��V�<��sq�O�3�.Q��v�����I���-G�*�S��I�D|�1�gܧaz�i�����s��S~�Y�⯦�Z$�h��J�6�$��SB���d����S�
���s�K�SA#�9߀�.�	�Ͼڥ�GM��d�<haN,���b�����D���ޒ�Y:�$ ͔G�����Ũ��֓�Ι ��d�S��T��y��h��3���7�r��(0�c���
�ll(�?V�I��M�Ӂ�j8��$t@��]��!~�����q��3�_�� '��<g%�_S����+3�.-\��s�<����qȲ#�T@�U IӀ��z���_aX��+�X�(s�W��aʛ�i�Ź8bA��z��p�����6F���\����G�|�S�s�?��`m�us-&�Z��M��8�6X�4�yv���)4��.�V�9����9�Z��q�䞺�sR[[�n��U���	�0��0�R��^1�$��+���M8�!�;���_�Z�4>�.�c�J�,8�Ԡ����5+���L�����%ݏ���w}�����<���1����������k��s׌���[��m&��$����Cm�BG[Y	iy��Zֵo��D"O�tNV�F�]^��s�Q���� ����&5>k�_�IY�v����CJ��e�HU���_�H#�D�A׹��ƻ�[�X�z�A�U[l�P#�|AC�`K���[E���v�+S�B~��T �	��c��)	S�E��*f�f}��ZyQnT��z}9����'u!
d�5|���VN�X��0�er������qe�$c��6�v5�
¸��E���,tߨY������H4I�(�2j�ΐ�!����0%E�����J�y�-3�Wv�PaZkRߕ�,�ܕ�B�Ba��cR�|���|;�6��ݐn��NrVQ����A�߸�{'�펣�DC�ՎJ���CA���:$2t�x���[
b�!	�Kw��ƭ�&׀���d3���WV?�#�ܢ���WJa�6��y6A4uwρ�No���'�[���[XH/i	D"�����4[����C����^`��,��
�'����xdj2��C�9!?��nuFS�d��a5�|7ׅ�脰��\��p[�n�|��ǬV���߱�%>����3��(�;���F�ܼ|5��k:n"�� U9}Ww�4xO����6L�d�=��|lg�,<ĚS��y��)���o���}��F�.��^p?���^�x��!CcaX�59�}d�5�Fa��Z��r<1#3b~�V���$��yL��B;uHܛȇ���r���⩁�qH�����b�ﮝ6z�z�"���bF�>�S�ab%�:�P�|B�gi�-�������Nǯ��Pi�j�3��.�:V�G�z����5�u��Q4�;Z�`�T&)6������Pt8��(�e�JW�v����1�w>*�.hk�x�0�A+s5�,cR����fNխ�,�)@������r�v���,�����Ygrh7��60�4�@{����}�e���Hk�
�\Y��(|�i_�@�y���&�&l�X�x[�����4	�f5��E��Pn��|�+<$��X5��P���������<��Ƕnf���ߚ���m�E,�X����)���,&���[�=B����t��x�K.�Lx�������)5|ʗq6L���w M�_���X[�YB_�n�R�K=�nG���ɪ9��Ba�2�d��b1�٣|Ї�`g���3E3�*���3f'�n��:�IV)H<X�[	JZjTP�0 �M�Iƙ����-�{d-z�n/K"��3xϦ ��l_�1�\=ʒMw�7ߥ��r�%S$�I�W�J�=~.͌-Ŕ����~�{�^�.�X���-�<Ȓj}�[+	#��j�J��&����A�J�^;�8Mzހ���n%M��a�:&��1u[
ۣ��0��6V��&W@��cK^n�F�����֢
.簿���(�c7Tff��
i���Ĳ�
�]
�5�]���~�"|������%Fi0d�%��2���mֵ����$�H�l�so�;�>6��>�8�h�S/�"+kˋ��c��.c<B4e�!統���pJ?�5�J��Y�ob����Y�����aj���0i�����i��_�`��	�)�_Q����\�I����q�	7��V��sV3�$(D*��ڔ��Hh)Q:v����k�ݓ �a��fܿ���A/b��5F8M\����7�8٧�=�T��!iR�?P\��㙚E9�+��M�QV(j���k���^ Vo��uM[q�FQ��	���/\&4pخ!�WG�fұF���|w�`}���di{p���#�"��A1�$��\U55����(�f�#{lޚ� ����(g��	D3�O�t�=ǣ0���޽�W99á[�4��%`
������IuEy�����ב�.M��F�-ȱd�{�څ���2Joe��8m�� ƙ�T�Ӻ�a��#��2J�鄼��I"n�`�@ly����v5/�&2�[�q����#�ߏO1�Z[��#}8�a����8S�e���)q�Q���Va��+�;/ekO���m{G�s)>F+��N�T���˱��w	��~d��9� k�S�y#�u_p��?���х.��DG���������1�����n�j�<�f�;�Ⱦ���-�u,��<�ᦦ/�/������r�!mY݄�t����l�3󏮴��$�L��l�.����'�J�lSm�l�3�MX�d؁/�ڒ�=X��ML������Ӎ�N벣J^�G2 Z{�w�j�M%�@�6��>�8�15������5�I���i�\��-�\>��Yc�$,]�q��88�t���Gί�O�e[>g�rZG��p8�I�}�d@�֕�-�,�<���sk��c��ׂ���E�,9ڡH~����>��0Ck���^0�{&O�9�3D���n~dz���8j�C1C��[�_R�'F :2D>��^3���vU���`$�l���KB�uF$��A%e�? ���n��`��+?թh��χnsu�H�4�� c��&�$��³��je����(
N���3b3���ZĒ�D��`紙�T�6�P�����Τ�/i����u�q���y��_;�F�?��� �Me�_bzh
��Ø�����b�f[1�o}�tmH&@��CE����Ss@T^k%L��U����OM�[$�:���Ml,�o1'����5d�⦨�H{BYl6Ӝ����ʅ��ѠDah7��F�6đ`.���G�l�YwLBZ5�2�d���>��WZ�7���/��df��8����L3^���9z��W�G9[������Ϫ���h4Lr��r�d����{�Iϻ��.�}x����V�|��,�w�-�K@$+ъ��=#t�J±��"�.�8A������<�o�)��O滀��,��C��-�Z��DXVo�x��s!0M��&��o�C����~�7������Xv���(|R�b����f'�E/�RQL� k%O[A��D�4�@�ǧ�T����+��2-�\�~o����gl�>=�(G'��O�nV�p��2�{s�����A_�7�$ewD���=�h�Q�3�ں���_ǌ����,�#Sl竄�*�O��������\��|1�k$�<��|�p��L

e<�h�O��ٻd��E���t�w#�i�bЫ�t�ՃL�>!8�y(�״fo|�j*-6�s��rY2��4b߇��A�����;� ���#*����ҽ�#�+	�Z����j�}e��#�_&�'�m3X�(�9��B2���jҽq��n2�+K��˲�E��H��j��5�`��AM�,O���{�{���Y>d�U��Z]7�zb�5�V��+�j�>Bv���AE3��M��6�(�7��o؍'
ߜ�>����W���H�jg�3��B\%��������bmh��abv{W��X�bHa�s����ʭ��?��NL����f�CW��^al"Q��?75��! @˩3��!�OV�C�9�d��T'Bu���_�ܛi�7�G�m��G���J�ԅG���{�h元ؤ+f��K*�������3��|�~��er�/�V4����o$)�K���7y��I�=?0���ҀKJ�wA�o����>咥��&x��V��p��0�.��}��ٿ2u|�H�ྚ畘؞��s��i���fv�P���i��SPَ`l-�K����I<��n�|��:D1���6�j�5 �	�zjP}ru�d��{B�k�j��rm]�6=#����%pB�ڸ�W��t|J=�^ߐ(Q�b>��ֿ6Xc:���D� Z�R���`8�����xT�[c���W��}����/��MU8��4��\N�i uqaAנ8έ�]��xS�$��h(���˿����vD� ���~�Al��G:6�*
� ��EKj
����������\���$H0�h�̆i���厚���8�d�v�Q4\���S\]f��`T�����~���g*��j�>�ҹ�"���d�bٞ|^r�O���
�%f�Ms�~#s��j)��v��:E���m:aE�|�.�i�h��k���x"�rK
KC��&�cKI^��( J�q�Ԥ�ɣ��.D�뭖�C�v�>�=3̪���,p�Y�s�Z�sk�F�ؽ�4d��F��Z�����=M��FA�q��!�(rO�R"�<r�"����n��4_�tx��GUB2/<-5��{�غ��A�ʚ�ߩ.���E��}�y#D�{;�h�p˨՗� �)1erUB>�V	��C���s;����Qp��n������d�ba	m����\4`�^�-��#�D�]v��m��8��g�����"�
�����S��*�W6ӽ7f"��4���v��Z��8��Cd����v��\ ��~t�<��f�r�`S�� �騰Ao���]e��"�w�Դ[����e,��쑱� =Y� gɈsE;/Cȇ��O}b=C�1�����C-��,2���T��f���������Q��B]�����|�Ŝ�;5)��@��8�#��,Ӝ���ƤNZԚω�"��*;_Ŝl��ӊ�f�=�i�Ej��	ķl���	:�xpb�'���Y�ȉF�)/�.<��ti3��1P�ϝ�9�U0�ޮJRE�������<h����vi������ie�1�M�PWbf���W�vs�h�5OWڐwF��5 ���^�MOs�t��'9��3�?�/�e7���+8���#��Fk�XQ�M�@Q|��vSL����vZדȷe����=�)u�^�.u�3�[��\��m*��;o��{��<��/:���H�����F����dO��܎�� �Mjq�4'�,�9��Q�B;l����ZuĲ�M>��/Z��U���˽��Kcb�-: �ɫH�z��g*@9$�a[�Z��c��0�{MZ45��Sp�9І�0�4ʟ ��M�˪�zZ��Vr��C^�?��cԁ���`�� �I�"�#��嶷�n��A���6<���Ym��e�ךyƕ�ZѢ��!��$�Hf���H�=�!��{|4�����Ǣ���hF��)�*�A7�^΢4ޑ�\1>F��� �2��o5��~�b@>�@QB|����y�:���6�sAbbt=�oz�G(�0U���]7��`������g�>�����ҽ���;
��*W����P�&�|�����1?���o�	;�i<&$���D���g�B1��\����E�A\�dl�r�b��x*��?���B�f�39�8�<�ͽH��LpYXH�c��LN��p6r��Jlѱ��'�E�0\�M�����.H���
!���36���f�𷀠m�-ve8�T�Ǐ��dA��NQ�"�"��D�*�rW� ��Ѹx�F\ $_�І٩��6/��u�w�Or�É���_�1Y������N��ѕ`�WQRws�޶��tPӌ��0� �T�|�؊&.����ߗ�iXk�y��t��e�M`˱6Z�Z��1�d��J|P���}D�T�\��&zd�(��TQ.�1���q�±פ��[w�3@J�.RFʭ@�]��a����f�!�鏐C�u��ҫ��s^�\�aB�!���>�Q&��3F�����7gć��R�����r�0�Yzѫ'��҅�I[���;��v]� ���~���[F�E����2�����4}��H�v���o�>��Ѽ
��'�`HuA�rea�i�^��c,�Ϡ��,�g�������oJ^����8D�Ϋi �B��}�N�Z��!pe��lcv� ���_|K��.�E�?���t�d��|qp�J�s`��7�t��QN��D�kX��'[��T'{%�����j��/O�s����hd�;�G{���E5I�xi8��Y;)4�_��*�ۣ�59�6>Ջ���D�����	r`>1������n@�97�*�٥/�s P�zSZEWmq�0HoʭJTG��,9�^�^�}���a���^)�F��RӚ)��3�_�Ui�]��&�l4{�ܐ�v{��˕�e%\� H����'2�/Q��h�`�cmAF_��h����iw�h��4@�Jށ,�cA�6X�j����aaq@H)F4���6�Q�" ��Mؕq�c-��;Bޅ�#W��)�N�!��_AD�X��}� ��kys\�C�8rF�Mv��Z^�̙	 $hY4>�u�h��@:���=��k��K���ʹ�=4M*�Wd��ʀh� ���e�W��b��|X��jA$��Z�T�ɪ7�&�L���_��.�]�����@2��%^uˆM�y5�g�QwqT���a��}��|J�F�X�MH,4�g���������'�[Fc?H�HB��T�5�E��?~��Q��,7I&�l'���)�r1�ln:���K6髬,1�y������8�i�����tZ���*��R $"(ρu +��/�*��1�AP�N݁����E8d� ����&.a�0B�j���3����E_�}��@�#��%�5�bW88F��q�ik_��x�Z��}l�>@���"��`��;w� �U[�
��4\.h�������H�[Ic	�ˆ��{��aP��ce��7�,׸�<E��g]��y���S����<�`;�C#H0��<�hA�U+��TM�!�B��'5�M��\�
�n��+*3tB\%��IQs1ڇ����dݹ�}�c���"��oTh�Wjk���5������{ T_�=�ʎ�;j�p�b�
�?|ǀu���₧1�蹝���2l�x%����	J����>$sDҽ�������B��Z���,'X�/���f#blR��T>@L�+���sb��s$q�	?��c7c�r��������tX�%���l��3��$d'�e������5Z)q��p��b��(V0Ǥ�kR�HQ=y�Z/����{3�<I!���R_�[����� Ip'#1�o�h���QO8?� ��!2E�����}!���|b5��VZCWA��S5+V=�[rv �b�X�j�f�7�(˓EW�����/�Q�-N�>��ݽhjh�^c�т����;"��g���"�p�$ƭ�4��&o>~^
�Z2�˔.�`ǃ��?�8r������Zof��)c��p��-�<�0��������/_ѫ��h�� s�)�<�N�yd���J��>_��q����g�n��δ�E'7<���g���泦�6�c�,�{��U
�bFz$���_�8�zL�9a����ԣ�������v*3�'Y�pdT�ϱ�� *�� �#ju��+p������ճi#�/vfr�6�D��	M��݅�t����g�S���� _1	���b̜�nP��hg�F�v�����x��E��mwo�J$(>��~g��C�oa}��蹪�T�u��jfW*D�2�i�ڏ����A�z�G���l��5���+r�c�o�_.4���������s�����TGM�g�`U8��CH?wX^�D*��4�0]�����+��;��J+' [j�#���(���*�sƂSaU0w�0�?��L�E,F[�gZ�(���Oi�SQvЭ�q�~:Fg���+�c� AKc��0 ӗWp���8�6A�M�"Օ���}[�������a�BɯPOP0,��n�2�!��Z+�pz��D�ti���¯���\
��Ң���lA4�+�}(K�F�o˃���HI.�b�>O1|�e�3��w*��n�����`�P?Qv�k��<���!�h���� ����eN�h]�騢���,%>m���nqy;J�G]�D�����xb/L��麖����~Bȧ�C ���"0��h*��*}�ԛ;���a�Ev�c@�Y]�����s,D)e�P�랧bX[��f����pv��8O�u����c|�'8���=gF���S�9L�KW0�6kw���B�g��5�%&?�~�].A��r������f�Wt�}0�RT�|t�����J���+V��9�a���z{�p6m\����G��T�f~���q���3�Q���8��?=�*�k9SZ�"؝��6�7��եi�5��͡���� ������E��F.��$��s��,���[��[��P��%M\هX�����]l>�� �NzM�J�"a|��{��貈�M��1N=3U����f&��SQ^��Z-LɌ 2{�Ѭ��.+�Q�����-���A������ �pF����S�َ0�W��vB�%%�jp�g�񭺇`d�6T�B=���3�u��&SU���7`p � ���֮��$7�X��Ҿ�q�}^�6���+a	�M��:QD�?b.R��jXF������%���!K-2�>�ZA��ܓuD�\��]�����W��@���'��2�.jf���2�15�|�ٿHN��>��܊�4i��?��E�ZWdfQLY(e�!V����nn����������#e�n�k4��p.���6�^���O`�]����D�a��ٳ�:�\^[b���$����U��]�B����9�Q��8M&���39�;	j �jPc��쭢xS%*M���˓B֗A[�I`�]�[8�h��Y��O>쯔A�z�uk{Wō�],����|�U&�?�6�\Y���"{q�������0�a�fW㫧mmᕖ��k�I��6�BA~W��%�R�o-w�@팱��۩��I����]��=D�ja�a��H��,�`N�p��,��)r�Wo]������12�
u=⼣N�|������A�b͆sE�_g6��T�g�)*]�����{����D��|��)pǯ�^:+h$���E�R7�G�h�;k)ۛ��O��K����I��eq�#��˄��R���� �)�ZE?-A��şY�q��*GNL�d��A�|Od=(Ko�Ý�Pl��g6y��eRy�;l��������(���V�q��d������o�V�����h�֏�^ǎ�-Z��`�^��MZ��Ҋfy�A�D#n�����+�ؽ�� 7��ٜ���,�̽"����-�vv�^R͎�$6Ӥ2K�n �����0/v���{V� s�"��
�� ֵG�[��'�U���@��\8j�ϴ�b�r��#�x�O������~{�X4p�%0��N7��%ǁ�օN�؝l �$:�����g�m� �"������Ds��|�Z�Ղz=�yM&�DV�ֵ(/�$�L�,��\u��%����m����۷[���Z^�P��.��D@>R��Ȁ|��B��`q ��Z����q�<���X�\��p!�L��cZ�bz�;qc��-P�`���.�]�![��yLq� Ѣ[(~y�໳���	�s���pR�U�2�%A�Q����Q��t��+q��2sh��Vu�J����E����CG@��("��0EPr3(�q����I&6|=���5�{D��k�4?��Y�������7F�G����O�j��"٢�Ĳu1>��Ga6�$��K4+𫤇�|v�0Ƞc�;u���t�E�����BF}xxf�ee�����<��	UIwԹwT�����	L������b���f�9�����
��,LB��e�mj�T��vā~�Z	�jo��mdq4!�P�4G���p�rM�AIa�uU�"E����# 
�f
>��2�ѻ�a�c���e���MԵ��G���R ��g��	�Y��V�,,v��-b'Z�� �y���E*"*� ��L���I?���pQE&�h}�7'N��JGX�ynjP&W�Ǎ�R�P��	�E�W|:ؤ'G�gg��,y�39�6��w5�������{�s�U�i }�Xy&������ms���N���A��]��iݙ�o�/���m�h-�#y���y�ud������!ˑSmf�AOh./�+�2Cu�\K�,��c�e_��nO��L�G��3��aO�����N���3��	G�E�4[�o����L�V���(��_AZ�Ⱥ��O3dn0~����*=K��M�[�۞��@���/BJ��Q���B�sBc�&��Y�y�t��Ep��uaA�T �E�^a�u�t�8<�4��"�mM� ՅG���dp�B�χ7���i����,�)��f�uC=_��MD:x�|���keg2�����Q�'����wH}DZ�ڱE���DC�n�h��lz�>�-a���ѥ ���B�^WOk鮁�Y(�pV8��^�o�σ�!����b���	D=�!ݛu�ڮ�+J�?��ޭ��j��'��H�[�l�����'�R�OQ�	JYM.�j��=ʓ��.�"l,�T�6�r.ք{��b�C�1r�O�M�NW�����+�e2q[�=ǻ#2����x�>�QKE�Z�3��.6+��+<l�>��L2�:i�Xl���mJ��7���qb�,^��\�$'�QK��G�".X�sV
����_W+��0��:dg�ߜ�[1�%�G��Xu����X��W��l�Ѣ�ҡ�"}379$��uM�5,ٹ1\���R���+��Kf\�UG�n������fd'w�m�P�۵���Ң�C�k}m.fL�Y�2
;k���E驫��h�{h$�N=���f��{34kO�N�69�㴣ze<�6Im�r����܌F���ѐ4�X5ꌟ���@ �	b�ፐ�EW����[����.B'�dT�f%I�va`xNK	�ÚR���-A����n{���Y�ǒ6��*�+�41��Y�x���d��݌�,���g� w����S��8R�mw��S�hI�3����ӓb����[��pM�7�Ħ�q`��4��:|U����98��eN}�aw�'��C�G
�>殟;� �o���O��o�1ctApb�:] �:�Mf�_|jJ��^��A
��}��M}�q�/����A��7@W%��M��-��<�V���/XɷY��uP�M_��P�@U���-}�`�_�R�`�w
U�㧟��]ś�s�\�%KBW�
�.7����z�����81�]��Z�jG�	�o�ڲ2���}P(���y����^��"�|,GK���]E{��YѤ0�,���^��y�
1�BG��.�h��y�l�!�ޥf�O�ga� ˬ�L��6��@����(�p�F���v�?o��	X5���&��9Ǹ>��G���H��6Y/���cg���ۿ���Ǒ��#�o�r���U+��[&M�J���%���@�]S�D�^e��jw��F$Y���4�o�V��;>2�a�0�)���5�~�@��/�n��lfM�*��/�l5b��	5�}2]�J3�l(.���TidR�&P�k�x�� ��6�^9���������	3%;;�r~pnsTݢ+������ȱm��١��q���u>C���ćCd��0pHӣ�A�ARke�rJb$��`�vR4+~�x�$郰`��GŁ~e��2�Z��|2�3��PW2���Q�>�2v��6��{�ord��NI���XYުn�6E��ja���8��b�t���wI<Id�O(LI'#�t�(5���z�H`C���E�-L��O���?K��덅��Ԭ�X��h���A��;���Kn#�3�[*��n�-�S~�;��M}Г�����-��tq�����i�5_�B^`4�~����JC.^I���e�Lh�?|�Q�	���FE	ܩ��X'���b$"Y6NG]�x'6D���;Z�{/�L#���ŊfL�!lN�ִN�?L /[&=M��=ö=�F�eo�ʾVUg3q���m|Sd�y�Hr��ȕ ��bW�b�{U�dw��3�ʁsD�
�<k1������֛��r�mT���۝��Щ��͚j߇�o�`x�}JSUqF��Q	�5ڇ&&�`�F�
�Y�.�u�H�]������{f({q�2����q�/'��>�Hx�A��G^�p'�Ĝ������z|����+���+J��� �+��t�и�K��]�YK�ID�����d�QU� r��-BA�"��^��"��v�s��<a9���_�e7:~�M�u�E��EGe[wzh�p��-[��N�@�w֞`a��ƾI�?�~��mU�[�xp���"�����Y�EvM���[8j,�[Z��d��i�i�T<tT�h�צ�;��Pv��@_h1څ���#R���'s@��H�nW��5�
�=���b��f�����\��� ��6[���g	�TC2�8v5����Fٝ9�����-𘪲��sW!ݼ��#��SڨR;���ȵ��qP�h0��r���8˾ڬ�H�T��0^��1m2 �ɚN~�0�zgК����NPk����Y����D,7�&����?/:����K��K'@T�N���g1Yv�w΃������|o/�t�m��"I+8?�z�,^fC$N�T�+�9
Ŝ��T��u�C���#BwP�0���
f�>B��Dԟ��>���P�f�i0�̠���Fa�VȪxK�%ղ�̤+ѩ�:�zj��gW�I7�n�\#� n�Q�[F�S�?"����fz:�b�Ŋ{��F�����k��`�p̬o���ӏ8��h����Yt��>3��[�0�+�������͍/���@
'��} =��#/ �c���'�l�^���Ė�=�f�c���Lql�s���k��{��	V�����TlŰՊC�7�8��}�6�/Y���-��I���13p�`��C�[��A�$	�"��� 욉�Z��w�o�k�K(�#��*�ߤl�Eט-�r�p3����RF?�*�5��$m�ל_rq��i���B
�b"k����G���
.�,հ/�q�� /E�q�*p]��2s�z�!0Mv�b(����?� ��	f|$�-�'�>��&fmFc�ҝ�_B�T�]'�%!��9pxr��c���aWժ/���7џ�yc4Y>��:�o���ٰn	�ަ��œ����R�Ρ7�&#{�ƽs��b�s��
��H� n£�xǤ��+yP��~�Q;��&��k�㞋���p�;�	�ž ��8����%oa �\B�1��%99���k.�C|��Ϝ]����QC�X��^B����'�Z���ե�)�M��,1�|	�!H�΅FPB�%h�.�1}`����NX��ݮ�	x���p���2A'M��f9fj�̴E����X
Bڪ�#�����g�`�烿�3�$,m��+=��6��#��&dg��D^����z�#�9��w��N+şU���Q�Zo<v�A��x?w�Je��<H�q�`&�bc��*"�a�qhr�-XHQe��������J�hX�P8��63�]�B%�B5�\�\;x�(�Mm]��f1MNHo��iV�%�\1We�ܘ0��J�Θ(�b۪ҋ���\`y`�4���]��^�G#|�:�x*�p�(��V�v9���,� �
�~`i(�(�t��c����M�BE�\��ڧ����&J�8`v�l���i僫6Ĩ�ӬA7��1BP^O��2���X�䂎4�s�[w�M��l�Gh^�ڽ#δ{��y��Z��y(dy�P�W�?z�^?,��B�j}��@o�TstX������ZzX���̤��3�4��%��ŉ�e$�eO��M�G��p��|��l��n/�[�4S�=#�է��tkf x:�����t)M�?b�����r-vP��%�]C�G��4"�x�0�׀�y,���B|�t�qo�D�nwWΗ�Yil�Y,��t铰�M��+G���Or�4�J��D[}��q@��������Q���:9�N'EQ18���7뱴x���x��̎ҕdf��3�����&<�a���*��aOϿ�*i���U�Y섍�Fk[�,j��&�	c�{�sj9�>PT"�]�@������M]�'lȂb���ʴ�+WI��}w��, |sERy8,�^:�u>(�y�0���2���r�N�]�7|�䢎�2'�D;�ī6</J|��
ŶӴ9B�ݢ�kUg�܋���ȰE_�k>���:k��*_�=�"�+?���L"��<���;����{6�|6j �4L0��	���{v}9�;v�p�����2$XZq�g�ǠW�CN��c�v$M.�l6����SU4�O/V�=���f��R�S:�����FK�(�f�Bގ䤔���=�vv���$1��W�/��8�|L�[G���f-��:p�O��+��8��ɴ�6F�5�l�@�"mE�f��Z?�H��i����c���Άڏ3v�"[�8���p$��T!�.�>�0�7�)U�j�8�Gr#��� ��a���	d��ߖ�o"�ݞ�U9����[ܦl	�F+�����Hx�����:C���N£�VDհ�1��c׶T�r����i��t�\q5@7d�*���s	�r�Ƌ�S�)i�J��6��{l�d�)�L��ڻ�iW~��� ��2ƞ
��\I����/JN�n��[�(�K�f�sd�M#;�~�d�����@��ʡF6�	��*��=8�SK�k����e�*��nw��'�
��wH�K��rX|p[5���z���BNxE[�D��Uj\Le�l./	2o�2/<�;����6�pő�lsVb��p�ke�s�dc��#�j�1�&��D�O�Є���L����G�K�ՏNj4���㍎jq)O����A�&�2�8�%�4+�F*UR�SJ�=l�ь)�J4��y!��+����v���$>�U��<L�$ҷ���,�Ew�ǂTK�NFuth�B�NPƚ�(oT A.�ww;���a#����T��w�:Ӫ�Hwf8��eS�C� �{_Fo������!���E4� *v@X\�0�rU���>���s
y�N�3P`���y�,��Ov�T�Qa��Li��qnL�c�,�H��Xp���?߀=��F�[�Zoie�ʟO�.�Gכ�u1�Q
�#��ۈJ��h,S<U�o�z�"��?��]�����=����E$RM>��wyp��n>rJ���ŭ�9��J���\�t%�Hi��9|S�z�KTI[d��x����½�T��;)�c[ګܮ��!
r��� ЗX].�s�90�u�-{9Q���-,pj����tѶ����Hg�溔�G��6��k�'KP<�&�CU�|��0]:굖 z��I�r.�.�����!���y;߷���U��0XU`��Y϶���Ң*A���m��A�F_Z� ��7�^}��V^=��v��$�O���0>��(=���g�C��ŜpK
�IY���l~���-t��P���
�u~�#C�h��9Ɋ�|��g��Y�#>j�������f��%ci]����I��@9���I��m �I�抬�P��X�\m����e $>�cb0���7Rpֈb��;̣R���o���fl���X�D��.�"�A$\�GݷC�`u���g���*�e_�m!0R�w�����HwIi������r4��#;Rc�܉��!��<�4I�,Y
����R>�ο��(��~z;��?K�<c��,/�@�1:#���{t�w�s;Չ��~Eh'�����sK�������]j���~�!�N/XS�6��r�m�<���K�ߒ�c�(���g����r��y}ߙ~���Rs\�.�_&}rQ�p�שׁ�M�[�ь��j�f�1���:�OC=Y�ur�縫V�ZI��E
U�.�����T�pp���ʤý�]s'��D�^�A���r$CԬh�HZ��C!L�� ��]�M��ǆ/"��9�E�v�<�H��2R�-z?�)���n�D[�iZ�k��bv���F|0��;]B-݄�:�d|nbz�����$#H]%G�����-!#�ho��v�26�^|� �����|q0������gS*������%/��,���r�H���)�^q!sa/�`���큺~��$[�+�^���Ũ	(�k�]h �q2��W���:dܝ��y|/����3�;@�e�3�c��\J�Y�]H��N�Hz��B�U���
��{F�] ��#���J��V �QBP.�ّ������}K�~Y�z�u@�I��cI��3� ���sq��j�a;i�f���:s~�и ��Z�%�1�{���m������P�ߖȼ��D�m$@z�g���T�@L�9�D�%_ 2nc��(/݀�W�߼��a��J��?	���r���������p	��5�BKD�
�&�*N��#�t�(�w�����Ն4 3w�^�0�e�1�wv�e)��L��E^�i�!YD,bb垮jEgT靖+�+L���l�Ȳ�b@��:zH��F��ZN/)U���� [����<�VE�|4I�,5� ��x�缡���8k����n�fG�?ִbF	��P]8(�)Ɔ0y��,���!�̞���E�k��=�U�#��}ӊ���&w�$�*�B]�<<_K��N��:��l�:��N~�Q�r���F�m��]�j!� O�e����>j�FީN$Yts�6�+t���HP� ��<.�D��'��<H���;|
ت5TJ�@�~���f���mPi���r��֮�>���ğ妥2�$��P��z��4u0s�'!͈$Z�г�\��J�Btg(��r�i��~J	�]_��]�*�vo�(ӻeX�X�|x��ľ�.҆�^����=�h_M9�����r��!D�t\��JW�����v^��7�#�fov�"J@�9�հ}r�$���}Q��FP��(�T��x�l5��A��(��z�/w��&
����#�1�����)r���oP* �Q��"H�X��:Ң>��7~�aǉ�t�>{h���0b��O���죢�3���⑄ਢ�Fcϑ! ��aW�#�+��i#L]�4\���+}䡦"Sd)�Ï)ܟ;ۅ�綆��n3O�<>*�F[i��ý>����x��5�e�_����˹E)`G;���(�T�Sk��Aҁ@F��3'_�|+|�֎G�܃%6���P�P��W�zw��� 賨��BW�Π�8EM0�Y_l�ÄA�#�S��lD<�At��sec�wT��.�˪V��E��9��Rv�jc����YL}����|�3�Hx�M�GNå��<����C��0m��l����	����Ɇ���X�Io�%��/��yA� ���2;"|��*wϕ����+�����PR+Ή�N�T��BR��}L\�e1����c��0M.)�s�f8,PK�����)PGin��FF�)R��E��K�>4Ns��}�� "�.�jh��5c�*-ej�6�՜4e���w�?�6����`��^GYR�^[�d9�\���BIL�7�@"�=p��mQ�DbH����k��m�^��"���(��S���(�nf���������sd1ݰ��jB�Fԭb� Pd?H�\�� ���:�( 	SͶ�g���)ƍ��٣�t$."ꇺ�x��F�x�1y����#��ڃ�2���.(5Gڮ/�7���^D�U��m���/VP2/v�M9i��赁G�h�,)�H�����*�T�2߻9^�#̠�'Q���	�d�oHؘ��**�U$ªY�m���W^�hA��o���B��ƥ�Ƒ�;�������0��y��4�)�R(�;�pUK��,�~�RT�췳M�&��	G&bsJuB�E����3�+� �_���O#?��C|��e��6B"3�!(��R�y���|p�Dl�JL����M�M������f��"j|�k����ݛ��Mҝ�C�-�W���P�I�	>;��*�O�[P��N�%׺S�]���/{?"�uy���9�mG^|��|U+{)�xa��k�{t@
Ŕ�ol��1$8�y �,��fXVT�H�b�z�,���wp*�$4�E�,D����ؑ^�/�J���!mZ��ΑI
}��r<�ԨX�KvwA�����XY���>	������R	�����W��'G�n$��Սݵ!u>��j��xQ{6
ҹ����Ae�P����r�&�k�jc�n?ڶ/��_h�o������1�z��i��4V������1� ��'��m�il
�}���.�S�����@�:Ŵ����������Mڐ	�&�rk��M��<�V!xW�W�T2B���~N�޻�5����(�PX�{Ͼ������=��!�B���b�MI&8����&&�ޫ�=VIuzzsЕ2``m�a{�����"o����
0H����А����1�]3倳*�Մ.��BUL�y]��=4��1l�>n���yx�d/*��z��cnd�&�*Ҁ,88��n��3�ꤛѤL���Sɩ�H����瘝�Ui���$lNf;�"ӄ��9B��x���5��кv�{ �I�~:̓k����w�x����D��`�٫MG:���������AT�@k���a��W�A@mV��A��9�Y�J����
e��Kx#�����2��k��8�{9���f�Q�i������
������BHv��qP�w�C-�OL8��舦BJʳN;���C��A��� Y�S�FE�wbڸ�1����ox;l�Q���4cw�ן�I����Rɧ�?ۋ�:���T��K[��\�wu���1w�i=�����k������p��1	X���f��q������= ��G?�UƑ�����G�;�1�U+GH�N8�]�����U�9���x��I�a�M)b��h�ǉ<<AG[g�;ٍnyw�jKi��% ��~�9w䲙�ܠ=�@����\
�w͎@hQu:��"�Y�mt��[a�G�6�<	�f�ų�+#���g�e�5Ύv
V���6u@l%*@�\�������s�6����C-�by���n/��8�|K�#GP�cE���Uo|#��_ߛ]��z�Kz��K1��Ws��fK�IaD�k�@*���t	�x\����9/	 A�8�s���5L΄*��B6��ݙ ��A<N�(p�q�|��)&������~Z�5�4��| C�+M`�a���7�|�y� �VS
���n���̥�u5J^g��ȚrS�y�U�t��|�_�?`��S���LX�w� F(ʿ�LUŎ���3tY0���^y�3���&Ϊ1yç���[�����@uۘ@(��Ɔ[�\�dy(��x��8�2������v�B��ȁ�e�W�Iu��zzp/y�c���7���E9�Xq|Q�C8g��kK[2��׼�Ld7��~���caK�a�_����}1�[@��$�H�(�V��qE
�S+b�ϟ��i�n�RC T�3e�65f�sn�
��m�]�G�� �m��ۿ$�~�A���X�lTf�߉!��aC0�-��at�2pF��l���Q8�H�g��w4��c4%-��ˍ4��}o*W(��!3�w�B�Xp��i9a�{�:&oWy@�	vCڢ��(q-��R�H�;?�MH�rI�}��d�[9�\��nڅ�jn���I(�����P����;�|Ԋ��n��ŇCA�2�!ǟ�'�N���_�!�ӿ��jR b�릵����0oR�1SJ/�h�b���n�G��N�����_!-���nაJ���Y�Zt�^%n�2��/lp�6���/g�C�N���cLn�ݥ7i �Y�<t���$Oq�B�6i:�Y��@uP<�W��*��zͥ�5�Pc%a��0]����/�KMQ��� ӫ�8�R��M����2B�2f����<�'�W�����,es'S��tQ�7��FW�[����g�g���<vF7T�=~���O�k���<��"�l ��ǈc�({��q8Y��W��(��<'*�YE��ڠ[�,p�F	 K����p^TǢ�s�ȅ^dzgnK��^߯teQca�o�l�I�L���9��]ڮ�h��!me��a�/ەb}�#��B�2J��{D�����8�ǦJ��\b/87��s0��W����G�غ+�"������w��DdX8G�y[{f��OTֿ#dt
�'�jl�'k������>��k���#:���W�����<�xF�����X#;~58��/b�s�����Y뢪�j#@k����e��������#�i1
s>���]�s�L_�<auQ:R/���<9#��ә"��������M�0�#���+�]L���4��ӑ �bG0�RT�0XJpb���JM��&T�D�]��VK].7	:3�E��[ex���dR��-m����FΐQPɺ����&Z�f-s�y�! y�ݣ�6�vs�+m�꓋n�T�Ez�Yݯ��~p�I�� �Z�v�
���WP}�3�Y����	T�4`��&�O\�"^������y@�ϧ�AB&�a
���
�Xb�l�n����sC��S(
����w�[�@ѬH���O
��D���%�`�~U��s�X%!��rk�arn�A���+��(�^����Ƶ��!�(�`Hĝ�|E/�����c/���[
+��"��G34h1��7_O ��B��/��,�*%GOZܼ�P4ߢz�e�ja�a+�����ixX��		�5�(q�Y��$� "�A�ÿ�τvR��M[Ji�<�N���f�m��b��q�O����X���&r��[���1���HԷ ���Cs[���R�r%�+�܉� O���5I�m}&7�;;�^De��@���C��^Т�����W%Ф�P��Q�MM��:�ot�/6Q�B�]�aS/�2�Y�;C��	� u��w��0w���=�R�E�z*K}�4Hٮ�˕�N�&m]�)p�y�4�N�Ba�m��
%��Sv�jg�qPx�u���厯�n�0)*�T���߭O� އ�`»:W�/)`@z�v�is*���Z��$Qxn����ZD��7���8�b������pUy^��%%D�<e�o�xF�ca��e.P�hVbU����^l
aK�I�&ξ�fq�����,(���t�:�F]���fߤ8ha�Ff�k20��|Vp�8.��M�i��� h�zOUՇ�e ���8lc��DXPil�s��X��\P��Q 4 i���q���6���g����+<���[�,@�\�@��e?�^��I���|�"e�}o&v��ww���?��2�v��뭗޲{a/������k�W�QG�7��:�w�Y*�^�e����{ª�G$)�D5a	dIB>}������/��=o�M�6�x�Nl������^_�����K2\�&1���g���ڎ�_)=���k!xɑ�T��eq%S���W����wJ��N��E�w@mSw�AϪ!Q�4П��y�! *��$?��������s�h��9ӫ�?F����s�[��.������us��-�z	ӫ{i���g��L<�r�>HX���/�9�%5h	�Ň�V����G�w��lܲ;����6��6 �����x-=z��L�E͌��`�����bV �f�}���t�l1�½�:����;�Ż;�0��!k��W��'�5�cO�JS(�%)\��r<�����Pi�Ml,G�WD��nY������A���Ux�������0
�w�!y�@8��5�=K|q���r��&��K�SE ��|T��<�����@AG��@s��g�jNR $�#D�%��8��Ⱥ�)AM��dz����^{����r2�O���3w���[;�H�Q,�,�l^�� Y"��4D�&��ub��L�dʻ��h�/��/��<`'��O�2O��_����_Qo��ԙ)0���h|�^�ki3p��60��,��^�P��ˏ"��3�p�,��k�{/)H$c�mjT=g��dYE�#��;�o�@����@ ��5J(�"}1�g�
���@bw�ߠ�c�Q���S嗊�P�H�9,�=CR�#� ���r����J*��?4��>۬*?�S,*�l�@��1Y4kq�Sfէ�a���#����8~�RRN����v��#�RE�<S�HO\�Z�X�_'��VptD���(��r�zB�Q�7#H�s]�	"�� 7F��[�������`���I�?��V�K(�Mś��J9O��?Ƙ��S��:�
�Q=��`���ſ�A�E�٠R
ߍ����x��kux) 3j�TK�}RagZA&LY�-,Y@�Y������$��b2��RXoh��T곜����d�q!�@���f3)����&��rΣޟ��v٪�i<3;Y��"���wum�[��g����Ǎ�	q�����ou�&eI���ɼwtPB���a�H>�qF���4 U��t�1v�������e�����
�v%uᵑ��:B'��$Ż��_&W��b�|{�E�f����v[�K��tm�j���⠢<ԉ��ы�:7w�[E1	r{4(�4��2M&_��]؛9�F�)�R�r�U;��-S�W������]
�o�NI#�F����]}q<�+�,��Fz�̋ ���-������RͶC�)dH����oƪ"΄#�!�ȶt���xc�˞rm��m�5�	m6КB�U�Vꩈ�qf@�grJԙW�kM�V�ug���u��S������t����J������B��Q��Te�¢���:��Y��yk��&T>����� ��PB�;�������Ka�����l9���]��=05r��)���D��J�'{��֥����J�&0|�S��'~	Jٮ��W����8���<@;
���vsG:[�RG�3[��o�RmL6v�������8�'�8#2W���/���?�:ݴ���������%q%�/6oyY�x��W���Ԭ��1���&�P�f��&�uރ�C�sK㮉�#�9�:�̴�C$���/�7������P���}���?ԁ�#L�P��4�$���)\	h�N�q��ۢ��un6f��ތ	����y(�����He��(���ا���m������t�!���ٽ���n���i�q#���)8W�>�،�}[Mi:�;���{���LKD�,���XP�9~ 	]�Pptҝ�<��;�"Q8���r��Ar��)��$9�ɍ�a?�Fv7�Ne@�Q���r3[d�М�#�ɢ�§�ǐ��~��(���(�ݲ���|\����_?Xk�ɦ'�2u~��_q���|mB�Cg���R�}fg�G��U0�G��Ǻ�'��1�,���4i ./�k��~G7C8U�ضE��(Q���T�K����~�-���}��;��x"�}���\|�&��<^7����������N=��d�Z���#�e`�xQ�(m(W.D��_\�C�;�����c�VT�u�xzTI��aϳ�T�պ
��]Ö�Q9�ٸ���+jX�=��v������ę��F�@"1��`�a����Qa�~�? �������=Q��!�-@=>)��� ��*�l�_�-טt��2�?L��(A��n4_/`}h�WV���u˵�����PU��T���J��U���Q�❵Ā����B�:�B�L���I�����/�!n�@�������:uy#��������9�Y�y0�5��Q_��,L� �w���L\X= I�ܪtd̉{��./�6���8D�����,�y�c�|��S�ףD`4BԖ]D�wT�t�<w��d��6s:oK'���}x�ޏb����d{§l���#��"�
�Z��F�9"�C��Q����h��8��L���$	���9I��:��$e.3��FҐ[{b��J� D#|�>�M8�/��\�E��yp�ǟ"A�r��E4��l�;y�d��p<������n�h�/�-�|[��`���}MO���0�2�{���ܔ�rqx-�X�t�
���P'�԰�!Ue?|7��\�mO|//M`f3�/��ݶ��2sh�v����k�s���<���ڬ9�6��Q#�(9.��������!���"�g�{������ở�I'��J�9*%���_:�s�E�z��a~D�i�a
��E%�恝2�|��K?���?�J�%u��]�}C|�}yQ��<(`�n�5N~�`�I�ޭ��Q-�pO��v�ycj��nd�w��Ww�H�eF;��.��5C���?�Q
�6�َ�@�s�LR~�ă��ix�L�:�����z�p� :+�W�W[��u�FTUW���(:Q�a_��L}���Hxɉ�9�.�3��{B��}�������+�2�j���)L�|b���g�U?���?�؎�Fo���)��2�Iuڿr<���n��o�M�#�^6���I^Y_b��}�;��J��y�ͣ�u�?��`�9S��<b�r�>����z
���铡� �ԩ��9/H/_��ɹ��X�{	�*�	��He$��#�ڏY��b�#�A��ÓV��W�
ty�g��,���x����j�����6	�d�����wIݶ�j
;2�ݺ�S�}��Tz��d��(����B�+��o2Q���>�+9��������܎|EǠ�e�3��f��U��{��N����g�U2< `	PDOb����D{!)����=��F�����9�i�{vy'����1�h���9��ڃ@͉}�+��A�'V�KEn��^���5`�8����s�E��B|lg����%O}YW���">���b9���
�Z��.&��!$�P�N^��$�:[;�Gc�\0nE)�H��^E���~�B��^C����f��F�g�C���fϢ��j���Tc(Ug��V���,�)�*���c�y����j�Y������&�<ľ�.f���Mo����=&e9��v���X�FŗI �Y21'`�Z����ئ<0�9�FfYd����8�Kn@�Z���n0̋%�<��U;WՀ�`��ks�I��,�b�=0}�����Ec��[�>j�f&dR���^C~�!�c[�"�2ݺU�O�˴�����*�wv�B�r�*Q��� ��?��B���l�� �ո3�T�.б6}T���l�t����޵��'(��_�,))ٷ	@U����gũ>:C[0sǩ�8P-�E�pux�%!��#[����81�%B-^������I���3�B�E�V��D;`y0Ł�J�,ܦQm�Xj,	�U�Zh߂�
�'�\�;�A���,n+��7DFx��L��o�#��������+@4�
l1L�^��7p�ļ@�6O�#��[�$i�)�z�����-yGw�]��ـB�r^Gt�gU[į� ��O���+���_eO����QF�]�n��)-8\L�e	`s_��,_)$X�i{n�A�V��v�ͣ�%��{G�<��Or &
>�a�G�=�nrw���y����w�O�l�*���uf��.�����x��Û�?�ErR��*-���%ـ>���8I�Q�-C�RS�M�.b��)c�K�_-ɦ�]�j��^� M8U	3T��dn^|N7�E =~F^gE9�+�CBo��� ������E|>�)��I��h����V�+�*��o=��e3�5ޛ�ɔ!Y�*	���r<�# s3��u���<"0�sKj}�c��K!�ݘ &����IK���_\�[��|�O�1/���^��M�2��B�?��"s���H@��Ԗ��!:�C���������Z��3�l\�*�=n�-�!j�7�6��yK�o�Y�� �u/�C�8��c�Ϝ��.e1�щ.�J&s�չ��'�X1��p�nB䱜��8\�]m��<����H�9g��p�%�'���|ƙ�e�o� j֞˺�ȣ�L:�c`ﱘ��e�'�G�_�b�����r�^�ID7��h�xn*��p�GL\�Q��9�u;>��i+�IK��~�N\IL������J���?3��{T�6VG-e�S~��Ο�8�;�y�,3����m�Ԁy��R�-��`�"*����*` !a�!�\H�&Z����,�?��� }�����y�Q�#���(^����4�ߘ����V��#�O�0/��_%��"���#7[+��(uB�#����W)�$�9h�6���?���lM��P%�4���Y"������@�q#S����\��"���7�x��ji��b�d�ohWɁA=F���`�\e��6�҅W�4i%W�]@�z3@s.޼� ���.����/3E+ׯ�/Oѱer����7�!r)�K�ţ��o�7��V+��T4�3�zό|�J,}<�O]�o~qy%ys��O\?Cּ��
Oa�K��6��L{;�>�ч��jL�}�|�,T,����9�����[�۲$ �HE�<])^��0�"Z�)�No��ޒ��SЅYo b�Zf�Ӌj#h��e�7</��r*�P&,��������\�x��˗�
u=ۄ=�!���*�?�x�J-τ�]�Sy�!��� ����}ZҞƐ�0!!���!��ڄr5U�򛸥MZ�B�jy����?/�r8Wqj�O\k�K�tn�C��l��7�ƢY�n|4��6"£�Z���O�%k��k�@-��7y_�����B6ʧ���&��_��mE�
K�h�&aɏ2��#�o$��=eep@k����+Q��O�i�0q�X��_*ʲ��.s��d�U��>�G�§����b�o���/"�=N���fa!���R��~�Hz��L<Z0�j��eTDܮ�	;`��<��h@��g���Q�{�m:��d����iFR'�1��ˋ�L�kk���u�."�������u���U!�A:4������H`2!J %a!l��/�Up]���KG[����s��m�f8��l��|�C���e���Z'e�D�	���QR2�{�,��#&?�8!�H��/�S ����.���ՁD�D�n��Z��*V�~1�|��hâ�sK�#�s�%~8���/�%���;H��g�>�ܦ^֝�E10э�yx
b�6��IIE�>�<�?�Ȥ[����=ٌ�V7 ���tL�(�[
�A3Ā;+m�k�Xl٧u��o��Dpv8��  uIBZ&&}��@�J�T���!�[���$��9��w4�)�r��r@ٟ�ȍ/���`�gʫ���+� ��u�qO��<�'Dc�@P�-����2�<x�4xYP%��CJlYl嗵����;�|�g!����<�.p�� $f�M-X5g�h�[YS���Y�n�K1�8��߱��G��cҏr��G�W�Hy�y��= ��C����{G�A,[�`W�2-,�)�C2<5xQ.�'N�����rqj��WQw�Ҍ�_�_��\�P9;M�d����$?��Q���~j��J�g�	��ff�-�r1����m��eL��d�]�q�q��}�}��>�5�6nc��������n�G�zW6OS��^F+p�\�X��E��P˧c�n-O��NYHց�-):��řۨ7��Bd�{�ب�ޱ �LY�2@�G�(&��?�V��I�Z#����V�;<i|=�o����)�@8�0�k�\��0aLL#0��՜�+�&K7��6|G��0��w�сe�yu�����$k�e�D�5����x����\j*���
���ݠ�xxϳT����w��q��+��dOf:k�fcq�/��g[(��ٚ��`�N~��Z7=Ū�p��(�X?���u��l~� S� �A9A+@��.��FB䩓��WR�#A�%�?hJ.0h�asc�cڄ9 �͵�d��� e�C���߷�K�sT��C������y�l��D z��f���\���6ն�0��-�ٽ��q�����J�X