��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0��F{��SUD����ª6��q�͓C��c�qֲ���L���i�UŇ��F��O�������7�sN6H2�eo� (MZ]uM8[�N?п^wU��E^B���P�������=<n�	o˪lr,��:ɇ�C�k_ۯ&U�t�Z{]`_���H
�%�-uV����[��A�c�a`d�L�<�:]ޟ��!v�<ފ<��3W�����[}�:��bS>`���v�%�E,T�π��mO�qؿ`5� <g����'XM*��ŏ��T-�W7���A�q�n�[.n� ���\t���	ݬ1e�xKP���Y�1ҧ�>��3�tO�����L�y�4?��-�`i���|���(���FR50z����$��h�?(K��������J,9"��+��'l�⬏���f�/O�rw��R�R��N_M4����ԕ3U���&�O��Q;8b�=�\��
~���p�۝!��P�@��O�?ð01��/���K���,�J�;�~��)q�Kq�����6\��e�q���/k��I��m��J��{�ꋕuz����/�5}�x�(���7�MX��Z&��ÇV��cN҄�4���u�0���-®+�ށ&^߯p|6�f��d��GXS�������DԚb�in��S�H�3�U�Y���h����H@�g�NVz���2�ͯ_��o�eZ��j�o��9,DX�Ut)]v�a��@X)4�/©vս7֘�!k����Jl��"��@p �?H1詽k��K�A�I�p�i�	 ȡD/�Y���n�A����[�w��(fʆ�,`<%��)�[haf�t`y���񌴸�j�a	�:��%[|��l����=��d˺��?$��58?���l�
*���R�̝q-\fC��5p(�7�c��3_��hg2��p��%���91�6�	�Ǌ'�=cԤ��0Y�h�=d��<o�m�w��J��et��I��C���R �d+�r��HGI�G���� �8��b}��Wͯg:�Ȣ��?��\�!3�ԓ[5!g	��B\i v�����zY��ᾀ�O�	�^r��@��,A�F>خ��aַF�.�����U��]8��a����
��C ���L|���J��᪌�6�n��?�c�����M&_���|�=b�~%�͸�f��dP��\ak�J��ܶ\��U��o�ҜT].���bڑ1F),���A����l� �=�D[�g�b���n.�qM����W�#�i�o����� /�:�^bHFv�|�Td�-�>�3�>�B��~`�Ss+�~H�Ol".�7�ɞ-]4I�)'��i�M��BŋQ��̩�(=��^ݪ��۸�E}F����Νv��n�^o	������B����#�z����D��O��?[��,ֆ��ݷ�Dvn��$.t�Ke�{����T-�z��횟n[���bLȰw����[(�X o�f��a���F��&��/=�V�旯?��c. ���m��Z�>��%�I�Gy�yk��{J�f���ܵ�+��>f��u��k(;N��$׾����o����5H}(�0/r�!�d~
2�w�S�y�X���������'��QH�pY�
ԵLK'�1����n�� �)�]�e+:��ɢ�4)=r(�%8�>^.�/-㋉^�]H�e�"3�H[�R��7�X��D	�`���3�}��?b���I
�����x��g.f�����\UB֎�x�h)�"�Dr��O�Ö ��ۢ
+7�i|a�Y���rz%'�4q�	�M�/֨��(G��r�������\�
��H��k���bI�s,5ClW_��5�˴?����-d޷Gz�5,�x�y|��}�����<�P�=�|D�=��8�QI���I�U#h(!kE���6�w��yy"@x߃�Y����@�u�Q��NJ��[H�t�r1|͋�y�}��Փ��!���zFO�r�-:Į��\����z�2}؍��1���y (�|�:@/���:�S�T��Z�$�p��mQS?���I@��j�p���-����)b3(A�5�.�O�@�Fl�U�	qV��6�Eb'��y<������wZޓ?�g��Β�=�|Z?A|�sY��(^3A|��j�O5W]GT$]��� ����d��']��N����VZ))C�ee��9i��͈��x�� �M�㰩y0<�"��+�:�R������e�1n�@��$|!-u�E�U^"��8�������ۑ
m.��󩓕v�P�Z��jK&�E-�վ�[c/\k�����ڏOy^�͗����e����;%��2j��q�a���w�ᯰМ֭����Ѐ �m�=���śf�)P�\$�n@�V��kh4�q6
B?�c��+�x�-�݃�;p��D��� ��⇨���>�f�Y���dɮO,?���PxR$��iM�eb�����������Q. ���
�'�a��bD�'[��~��p*�v�k�A��}Ԡ˥��(� |���m;�ޠ�$����<6
Bp��x*Ӫ������9�����V�.{A�$w
T��>��A��}�9M��c�
{?	L�������a�Vd���R��(���G�i_L�0��&JB ��g���E��c,Gؐ*��-�� �_d{l���.�:'Fo����K%��K(����x+�_��oxu9zx[Yi�u3���!R#�l1Qf�`m����Lۣ|�YɌ⧤�#@9 �	D��pcU�x%�>���c$j�D�9�H!�h8p�*ۦ~m�X�kd¼�rǂ4Ka��}��?�\���=w.�s+���}{��M��W���h��L�f����׏�9>�.=}H�����h�6J
+y~���M��Ӈ��5v`�U(��OEK�Ԯ��m���lRR��{�����Q\��*�K�����Pۘ�
�v �P�P�c󖪳i��w���c8Zl��pR��A��`$1;V6�=�"�|��?��r������!O5����O������(>���Jo9Tf|����φ�kq�BŐW,#G(���f*�4b�%j�aC��H��cJ
�\����ע�83Nv~H������4<�2ʡ��Y)Ј���W���nÊ����[)(�jYWܠ�v]���Uk�{��(��U�i	����c@l������L;��@:�Z�&���Qv`�	�S���"q�	LQT`��yI��Mx��I�yS;,'dפ�-s?�2��HE2zu�~4\�)$�}qˍ�h�$�"�=R������ l����gV�~J� �zl�t����cQ�\��ȡ��lb-g�r�c��~p�M�4�ůD�7�b
Ԟ:��V1�c��T��X�EiRI��r(��UD��#�Zea"��|Q��b�3�78L�����=2Z���UD$m�5���aZࢀ�p>	O$b�
���E�����^� D��%X�Z���i��n�
���/F�dV�m�CUK� `)�R7=�v;�gL�;ʼ�fg��992ڈ�ٱӍ��\ڊsW�@2��W�-�An�/F<.hb4N#����:���#���'U�������ӞH���I�8�Z3�9's��m����D��݈�IG�T��m}�&M��M�=a�p/��u[�U��,*Ϲ4�G4�����Z6�qz0S�䃅���Q�'	:�t���ڸ��,z�ˬ N�d���BbKK0o�<oy�a��+�cѾ�!�䶔WD����Am�+{��+�
�h}v��$�0��m���!|z5>{��v�"V}b�2�҇�Bk� �〵�C؛��v������F%�a2�['���z-��v]���7.�l{{�$����w�_�5�g�g�.��X��X~��<���d抪�b�<��ʝ�ux3Z�Zm�bd�����Q$�I�'���lO�ߛM�π�f���Y�	Iy����f(й���%~e{�T^�Q��ꂡH�%IPb�������!���Q�sI����\P�i����rm6�c��g�(���Y�+���(Ѵ������9����p	>>��\ZN��Ɓ��;�dm
?V���}�Z�c6�7�?�B�]��e<*�T����wl��_���R����c#eu���lG�X�#@\nMچ��������gOܴ�����}3�O��%mT4�:�P�Q������N�
��2t��z�;D,7f�H�OFb�R�(y���C���+��/�[u�Z����+�ɥ���E_FJ-Xm����_�&��T����u���|�+[���Ǥ.22���5��x|��|�wpp�ȼ��dҁ�	�%x<f��jz҃i,��r�'�RN���<�alFiI"�Y�
�PԳX>U٨�6�,	}1�%܊����T��@ڍ��~qM�j��F6�A��Pl}���h�xA:%�=���9����p�wF��+�������o��V��Ut��T
�+�,�Ki��&����k����y��o�%�G��h܋3��%�i������;jK�U�E�(��D3ˇ�Nc>�otL���)U�l�.2c�eb:�!ҘF#B�{�q-Y2�*�}�{P�N�\��P�{��8]�[�9�X:&Y���;��GR%ӡ6�NK�n�ꇜ�G!��*��:D碓kl���Kx|�[�� g�1�0!C��������T+(v}*�&D;��9�Q��n*�428�����4E�4Y8�\�
>D�v6����
�܅QH�n4i"<��A��^�hs�=l=f)�"��_8˝|,P|��Ob)G�
~�ל���,P4�-� e�$�����q+r��D�*PS�di�`�$���'j"�q�-�;��6����L��^^;]�;���-8�p�ҳ�/[ѐ�	���,��lCp�x���~���=�U��$H
�d+4t�y�e7�#���ymp,��{�kD��]�u�_R��߻���
��zq�����_3�)��b��ٽ������R��%^`H�sp�r7�e$�3}��u��­@�kn����k���ʩ`1A��&=���0�=�8�C؀%�(P��3���&T�����F�Ul�ql!�.?^t4��P��}�ٲ7��CǽGg�8/H��D��U�XŒ3e�����P�/.f+���)�Lg��(l�˲���kUe�W��j-y�pB�����<ʑ�̸1c����Aŀ�Fn�U��4'o��t����/��vH)��j�r_$������yѐ,��%�F$F�����[e/�޾�~*����*c8�y �$�vf+���ZX#$�Hw*����^�7�0���7����*y(óF�B��.$J���	zl�m9-xt��+f�!(J-��	�ަ��''J�z��}S�)6˭/��]^���b��/۷z~������f#��x	Z��:�
׃.��TFn��#Iȋ��v���3}�n��p�/	��.v���t��{��8a��ط7�_�b.�U� ���C�aU�N��6�p󗈅xx�W��[g�b�[o�hU4����B��g}�T��^��e�r�G:m���n�w��7㞈���aХ�����Q�^Y2m��;��/;����7�+..�$,���;�<�?��v�o��۱��. Yg���l+�����;��+ ��@Ȩ�4�H�љ�").�뇳�q���lwm!>	��⽗bCdxW����6���9"F����B����h@�|��/�W����lZ�p�^Y
ݳi�Z��bUTcK�??A�y��8�<�
)$��|�B^8��"����!�,�]�ȕ���o�%s������q�"��ȠƷAb~r��ϯZ��4��8�OGEt���]�);�U[�8/G��L��&�ˎ�9	GH'��{�z�G(�S䔑wR}� ���+8r��Dj��'�B�`�V4�uBq����(����P��"���x/���$�e�z�7F׬�9��8�H_l���;5��aBU����{-c�߀�d6r�]���CZ��ng��O@�� {$T_��`(�����;"1?H��|]������a�o���RJ6�.7��b�yNh��S���̟
7��U�6� L�üߎzգ1�E�
.i7_�4���;�Ҥ>���Yx����d�B`�} @$�r�{m�H��V�\�����]ʯ�Tʮ���O�� ��j�rB������g�Oڭ�g���y<�2@��ۑҘ�/ �Ia��rܼKQz���_t|G.˴#�k��%��x�zqJ�Od�8��~��?~�֣O��VP M�ݬ����~Z¹��;�uF��j&,�㹶����2�mv��~��P�E��ğ��@�EM��(͋mX{T�"��J�7�0q�ƣ�6[��
�P٧ �v����0��)s��'�����e\z�����+4������-Y��������R�1��*�D*ۙ��@�,����g2Z�7�f*����H���q⠺K������3Γ�K��H����S1����s���рf��?)?�[��� ��2�mPtp�6��&�Ua�ۣ6!�����4�:�5��u�|��!��],�����
T3p��y:1=5�Vr���׻B���}�8=0�s����o31� �t?z֩�(��O���q`ygϩ�5�S6�w�,Jޞ) ��,ؘ�à��K"�z5>�噸�I=�SK�fӮHT�=�^a	+�+�
)�th~3����w�͞6��n\�;67l�["�ɗ�"�X����WY
-}2��G |T�#9�о�nI�R|�np������W9�`�->���݇}�PZ��V�Ճ4_�qD94e'L3&�ƎS]T�`�wc���a��5և��u�|?J�u���	�&QA-d���c6�G�
��*�e��].Oy��î��������;��v��B]��W �ד�f�^�.D�~�LG�(!�"�*҄U���C�ɸ�mθ%qڀ�XpW81?��D���=��=<R�T��M�;�㉶�7��Jh�����V����ŊQ�O2�q�����x-�.�)���$��G�9ѧ�Y��jϮu2��f�
Xν-C˲�@(̈��W��(�A�_�����ᯮC�-t=?߈�BO{`��2��#��Mp�X`cV��@��vq�[Z��6=gX���z�S�� WW�9g��p��0<��H��5�D^�&?�5j�$�
v�ߕN>����_��7��#\�мw(�u"�7SV�>m8�"�6�������\�b�tk��}!���I���۬}�ƸV����������Q�A>��B��iW�U
Nsw����ש;���E��i�e	�j��
s�dϮJ�w3�sHq��^��+��~��t)�f���T�5��9�Β�/2zt�W�|�D�,���F��f� ������[�r3ȆwvP��ʵ8N��\�w��^߭���د�Daa�$�;^Wy5>�լ�ѯ�K,	�Z>��O��!�b����'�6���R�	�	e%H��/ʎ']ImC@�3mq���@��"T.A�Jaa��N��pgc��g�1���MlD��|2�K�j�����Cٗ��z���ZY�`7���3��d�T�5'��w����{z�3�L���ۃjuxl��,����o���&*OzBʼm���ˆ����fP1?���K�7y�կ ����y�c�/�� ��4T�X��=��mܡ ��?���c�)f��7�>��N����n��[��s7h8�0\%�6