��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��?x�?��Qj�2K��F,?��D�.�S�=!ʞ0]>��{���|���!>�Sv�e�x�X��O�H�`Q�������c&������\`�
V�	o2�f��.�Qv�nk�s�*��4���<L�Ԝ�Z�$	�
f]9G6-B�����>�A�v -�:��;�7n�G
���ٗ�#�yء��ݶ�n�9�W_�E)�">�8����TY*$Z�ͦ��H��0>p\˸�y\�&ɷXP�W4�^&; �{��rZMY�CH��������z����� Է��!��JB=T� ge�"sF�7��P��CV�ȕr �����s��4eZ��Þ��ۻ\�y}�Y�A�+L���A[�\�/�����`��%(]�P>�N�S$ZDF��|r��<�$H�t�/���*�V=��_Q�G����|�:&aHp�f8��}�Aϲ�*(K<9P\��?S�����!X��v2�>�sJ^	v)i�k��n�t�3�:�b�Wp�n婹���%�TI�� O.�C9�X��/�c���*W�u�8<M�׮J�m�$}}���dR�o�XGOA@��������p��(s k�/
��$��y?zJT􀩢OѠ�"`r�*l^?ɟ�E#s���~K9�Bzk	�����p�"�K���B�\����a?�kn2OV:�,'ݳK��v�i���pe�I7N�I�+�/�&u���"tb�lZ�ה�����C���!vUCZW���&|�e�;�����.S��51�7.��$�3��@�������)JN/R/��K=���'XG$\�K7¨���v�ʸ�x=ۤ�@��ָ���[�����'3�L���M��Ŗ!�,:J�����'��9���mQ�0�B�ju�љ���s�W��C���D�a��|�4ˤ�	F�X_����@�##��M��5�#�O��ą�W�ŀ�m��Q�Y�ǝ�x��}��GL��n��6��-�O������v$�}^��9F������ؓ��Ϡ���M��9m�v��L�c�g�����|�1�
l���٬/�?����9߫���̴O*:�Q+��E��g��o�\@�<$9��7!y���
p�M�嫁po;�%Q��Q�i���d̪���YJ��G-�p"Ul��=�Uҧ2���)�9��SQ^�j�ݛA�k�:ڈ=)�"[�g��!�l��P�������K'Z��V�YNS^RN2�ȑX�ִS�λ3n�{Ⱥ��㟫Lg�go8sɜJ��� �#%��Ɛ����>�fAaw�l( �p��^��a��M�1���O�S���§p��V��
ƥ�x�CQ����7k����׎P��EJ�9.B���������`�֤0'\w�n~Us`L�Fα?0?[�c��ߐ�,�T1��~�c�
}}8��΃s��cV�x���,�v]u���g:g2�'��w7�]z��9�*����/1H�;W�+��·W]������%I�Z2-�\�i�
]rh@�u%��-'�޹9�l��Ӯ�3�`��ﴜ?���ݾHԪ�z
%Y�S(m��x���ѯ](�����E��.x�	�aw,nQ�܃�q�H����[�������y��/��]�;T��gi��:Ef�U��Y����;��N~-�ދ����"È��O=4����di�y�G~�5t�]Mh����s���l/1���	�]����{ۿ�4�������O-���c(�����!`/��D�Wʈ	 ұf֖1��g%��C���Y/Dc���m ��Ҵ���
]��O���ڧV(c�g��EvB�ڜQL��u��%����u�����D���y�$��-���v*���_�E]^���R��&4�-'��K��otCqxb�����I1
	�/�`�Ɖy�z���Zʈ�ss�|��s:����5m���#����5vW�-��A����V(�.�@ٍ=��,�M  �a��M;p�j��"'���j������fҴ�؀��^/n�;�I�AǳG�{�(�Z���5e��7�Y)J�z��K����A6���	�8�j���C�$����`G�4K�-n$�+�Ål�� �E.��	���N�*�U&��֧_�9�a�/s��0t���!m��u25c�~xX�o�����U�i�y(�D?��;b�M�E)V�T+�5�L������1�(��;�F+P�� �NUi b�� ��)�a��n;���d�Rl?�ɫ+D�2��H���r-��&��:�<./4��L��Ξ�(�����rv�ۊ�B��ыo>�yI�0��}��WZ,Z��r�*��3�=��C�L�����)cZ%��lf��4*f�;�F<c�f�9�9�� }$����^�(`8���,�QX�$�k�7��D5M��4*�.
pg�z"/ ��`v�w� m3ܾh��O�"��V��"�%����T]�e�H�ճ����6��eT=�9��H.�@��`��2Hu�s MB���9����S��l.�=N
�����q�67)>I��;�t��{�b����V����ҕ)��}���f_ �J�w�8�M���@j��N'�kD\s������'h�1����Q���_���;=�T����7�"k:��QƯk�-
�]�	�v�ٙ�w����9���m m�\=�;Aq��m�+1�.�$舡(��C�WEz*�Sv-4gE��:n�c)�	&P�u;9�gV+P1K�hQ�`����vQ]�*��h��ȴN�#\��͵$ӺV�ag��	(�{5�"r
ɼ�ޒQ�/u�< �"�e��a�lB������YNo�j��e�Z��[�U�G�r
����U,���?b��걾T�2P�b�Q�mD�8a���ez{HK��$
p��eŤl��v��u��6%�$���V��;�,��uN$�a
T�~�E��u �~O�xU~��S-w�EqC�#ْ�М���_yBo�+G;� ��؆�6o]�6�k�S!7j���(槥�85�O��wOfU�p�1���2��Ӡ�Z9$`�w@���|9�y���u�IU��0	/
���g����Ҵ�V�Po���޷��g2�Bd޳��\�Vv�����4�^��::|m,��/]�ػ`������5�a[�|�Uan�8���R�m�&sT��������S�H��e攆��8� |���b�d�
䬁r���8���NH��4��%�N:���O�sj�0�-�Y!k�,� }��!�J�;�`	���{�>`��LϞ�����{~+z�Wx����¿�&���G�E�'����Ͽת�����IMk�[���	��XX�].\O�h�̻�$E�T��:�F3/J�?����"��ߴ�uFa���Q0Y���~x	����#+��K�.D��gm>Y�n���[�W>a��R�)eIzÉOc�E��qC�$ב���_gwu~Dbq��Y �ik���E�չ����Nȫ�o�Q��[nb�x�H�cn�)on��Zh&����ӢZ��(�o�ׄ�Ū�Sߐ�`�O;z_1���}�SG�A ��a�cǆ���\��fP@G�S?�Ei�jl�yXnLʞ����@7L���E�ܧr7Ȼ|"z���a��c�w6�%5a��È=o�d�tފ=$��=������D*::�z~6�E0��ݜ�L��l�CӾɸ�F��MͅAY,�v����B*ȥ�
�O	�;�b�/�Z�x���T���{��%�&ڽ�@��My��ɼً���c�c�-��`̼��5�V���q���N� �=��]2��7U��dyd�W�,#�-���J!9X+��&�:���m��},
���T�f:\3sA瞒���%u�5���@����:,MK|�"���e�g0Ը���ccu�\�9����]�pUC��*�+�Z��\{Vd�ӕU}_��,��.���q5Iڹ"�Lp5�ڧxj�_������	�x�bT�3��rd�������3ት=����/�s>�#�N0�h�I>1p�xh�O�{�L}�ƲP�o$�ĩ
QB��a]��}?� 6�\�[׍��%W͹?�?4�]�lò!��� D�nx��=Y)�4�E?d�H�}��_�i��������jf�7���U~8���j���{ES��ON�a�4}>�X�l��~x�|Q.n��[{��Q]�k���#��o�&���q�{�/}�r��K�L��W62�Y���MG/�
�H`�^}��G����!6�
b�q��=h(m�����E�k�1N�����Q��V��o�hC�õs�[j�(����V���?z6DI*�����0x<F�e�M�?# �ýC9�w���O�����M�3��3s�X�D�u�B]�yRBm�)��:?S4��w,��&Uz@�����r����-a$�5�,%��ЙcoS��)�p����G4��V��=l��ߴŘs����vc����u�ш��������ͧ�z�x���fP��(j�T|w{�o��-�e�^�tL&���q�%�a�K���,Or�$Iɧ5/�G��ڷ��->�sgH1�?�a^�PXK��2�����w�Ty��v��� ��_��Ŧ9w�5i<v�S�ح����sU�j���0��:�-ie���Pk�w�V�t���0 �^r��&�pMu���������w�B�0z���z�B&�}�i�K%КHm�D�+�{�c�J���~�����O@F�{�2��@�ҧ�aN6��tF�PJL|�ƶiH>;p�*��ͨ�8@ۡBh�8U�U�9#gx��u�"y��TJ�a���Jì���E���F�^�r��";�o�s%@`�!���%�`����VӼG����zf��M�A�6�	2��F�����ío9���J�{���>�#=���h��-7�h��#=p�������x�,>��ŕtSg�jt�'���>�c24�/#������>�*T������ �W��}�
5q.�$k��LU�WB�E���޽.2'���vr>��׶L]����ԯ�p,Qe[�3D�J֜� :S�$�Ο}��$��Aix5l-F>~~iAXZ�W'*#GPr7��n0�4_ם���A΅�+���p'������{q�>*�GBL�c��{F�H}�������&�n��M"�*�,��o�Kh�1�f�}0�ZvJ�fN�1�Y�h'0S����>����ZRE`��|p&Q}���8ֱ��0Pd9.`��+#2A2�6���f�(T�iV�g�v���{������/��<�����u}��w;jD~q.�ѩ/c/�u^����u"|hr6ʳ����[+D�����Z�\kAW�ޏ���!*���MDb{���w�4��& ��7���qѫ�������G��qx!&ʚH4o�{0R�ZcH1a�܎��Q,r'!ZE��b�lpu������;4��
���)n�A�ԇ�P���^ל]�$�x!��,�)�;�/W����ް$���ӽߨ�Ivp1���0'g��%5�=~�G ��T�SO|c��ft������tp����3������[%G/o
_̤n�4j]/< P�
���� �4S��|Zހ���{|��oI�A����������RLv� ��y���fcc��ɬ8q~��Vk�z�cF>�گa5��
v��k�����p��E=��ҤD�ʏ�s/�%Fݩc���*�a��=�����ƺ[��\�GiYJ�P�=����T�H�6߲�7�8S�ߙ�еf3�7�(���9[c��f�4�]'`�V7-5��Z�U��_�*��B��Gh!"�Yv�K��(r���,Ȥ���oxΰ˷;��Z�H�l:�1��36��#����/d��������r��`�����3 �L�����R{�?��!�T�_8~�"���^`�3�ri��>*� =_�������݉�v�77��:��J3,�|�-���3��>�@�~����8=(�\�"f$AQZ�M%�m�(��b<�M%�b]�� ��,��h[F6�M\G�j�r|��-�ɤ=��>/]r-_�F��6��E�7�l��`dpV��pC� -(T3�
�nuY��+���ocVXkn��XA"�h[��R�A�h���D��O�=�\|�HD��m�_�
P�ّi$ƩY^K��C���In4F��V�*hx��bM���c�m��?��;X�Jͅ��nbyP�tT���R� ��9jX��z�7�*�1��-~.����lZ�#���*��ը]%ف���r_ eN;����R\�ōe�ձ�i�R>�Z�h/�W�v!Z��>K)U�6S4UI^�ͧ2P�[կ�?����q��#PLV!8J�5��}2��c�n멸+���t�8}3��;E�c����ev?/Ϭ� xf����7������dЇ�B�?奛ʖ$&Tɉrq�:���0H��C�WJжW,Zz� ���9�V��1&~��"���U�~o��� ��	���y�	@x�+D�;���M�V9�b0�V1~�(cK�"�p$|���\ꋊ��Oaw[7-�v�Eic~�V��z�(����k���{��vRa}�H�բgN-8�G�I�g���x��PT�ÿ`́����t3M��޺2�Ͽ),40��Q��j��G:���H�2s�O�O�9��A�M�8T��5-�׏�4Un�kc�q�s?~��O��o��7�����N������������:-Z�s\j.���-�v\�?r��g8���g��:Ǥ$~$R���)�?@���rC���)��j� u� YcF�u8�����G[0`��㾰�_����PO�󴯚��4/�[B-ɔ��3G��� ����y�βM�l����>j��j�y�E8G�Cr��x�c��Q��b*`�?�yp�,�R�X�t2r�k��3N���4p�'^_�ϓc�O���
 ���TX��J�'�vǺlQ"Ҟ�1K��v?i�����sjG��;�$�)�O�3bi��qt+���7��EA���@5�,��G���*���i̫hd�L�D<HS1�P����A:���VR^���bF_��"�x`��+5��.;
d'�����XW���4N�~�V9���l�<�}���:l��b�Td1�!Q��	�&��E���+�G=��ے'W_h���,���ͭ+�8�(��+�6I�j���9�U�%a�M?��-l�P�?3Y�t����d`I�3bLFv:�H�a��T�SS�{� )�שT�L������#��%��iD^�}�N����t����	?�q���UnP�I;7S��89�^G���P�9�,�*7.�e�(D�h�̻]
���� ��h����sCCS�=����9��S�/��o�;؅h]P{���+S"�Wl9S�D5W?i��a^�8��$�^Ģ.����t���-�מ�|�+�]g�A���L=q�X햰u��BPg45��;��M���oљ�m�Hp����yy�E��7-�0�+�{=x�lR�� d�L�	���7��FL,�f�g�(E�^Mic<[�1�:I/��x��恙�ˑ<?����]@5�������@j��9�MZ�@���|J/����I��?���"�ׁ�+��јX�����"M~���Kp�R�N�gXC������b���qZZ���NPi�~�2~��ә賁_�Z��c*}�B�Uw��r����`�ȔQd��l)VL954��黺܋�D0
�cS�e����z�<K����� ���5X������ׄ%�X~<dI��٥��Vs_����H[n����Χ�Q����\6���{�5K�.u�n����1�x̂�fÃM�2��ON�K�ZO�qJ=K=&K@�m�|�ژ*���m������IE`�8'Z��銲)��q��`R�vbL]���[��it�Lq`/�w�7ԕ�9���m����UG�8؝h~	��ƀ�=�	H�c��g8앾�\B :��'�(e�?����v�l����=�F��x���ߊoQ>�P�h��&�ڙ�"���̣u���8o6Ҝ$��F
�P�ʃЊ��Y�~��4��
�V����W�#�rz��C�)?X���&w�k���~n.9��L��5YJ=aL�:�� �'Se������W���������82|W(\���r��Bs���z�08���)? ��^3�
E2��)i�on|�'&��%6Xoq�<�n��S��j��s]�ʣ�F
��n��'����$���s����ᅚ�mȸ/Wod��'#Y�$�k%�7p>����:
�
��ZV4%��
[x���4�/1 |M���Y��)��>�����獌9u/����ڬ>e�L�258�a��1[Ay����񌰕ă9)���a���ߍ��1���~Vi�hNϴ��#鱺;eՒN�+���N���٭`zC>o���ٜ���^�l$]z]�]�o�c�ۂ�
1��ٱ�ix�)-�`�|g��!/9�e��1tjͦ�,�9,��<d��V@�a��Ps.�ĥ�m�9���r\��3������bz����^�"E��MN�6�|X�8-�^Yٯi�LZupL1���p�B����UW!�*uD��V`�Z���UU٠�n�4�|��._����%'Ʀ�x�"���{j��w 뺕�"�׉�D���u�=��ő�5qA7nVj��F���b��2޳l����|�sߔdRN���>��P~ZB��OC�t����s�]���h��$N�P��(��&(+���G<�Zo�}�~��UN,NވI�#�/g{LNഖ��Z�p�]��Ⱥ�P �D��oݾs�2�>Js���'��@�~�����r'Z�
��#u\��SЮ���y�!C��Ɲk��P��/�(}��(B�_t��}m����>�gbc�j��:�Г��4���+��G`�)�y$ U˘��BHB��E�,뙾�U��D��SF㔏�|#����W��J!�-l��5"�.X���x5���9��!z����}��J!�9M̺{�����#qr��qf�fCR"��7��5�Z��r��������e��2s��g��9'}z�Ǟ�r�3(l���cAc�$��G�@ 5��lU�P��I��cL;Gm����?����WMf�Yq ql��j��Z��P��+�\�	���t�k�}���X�$H�k{�&P���5�˖�tĦ�(�-���X��v8+b��N��l�7W�U9�*pv&��Fl'	'o�Fб�=S����|&@,�uG����h��_�g�Z����L�m���N���H��.���un����V0jG�㛡1`@GJ���ͯy'���
�|R�U9���3�_`)'��=`�/�q�c�e]�9��]$d,C����D�)sSZ4�&��R��!��߷��V�5d����:������A_*���p�g8
K@�܁��f���ҩ�X(�$��oLLP]|4�0/��R��S1A�c#u������wUf�6�~6�ťǹI���}e��Ae[�z�<u)��Tz�Q���H�"��K��_ð� �[�������m@f���������ഗ�$���ل�,M�d��SN��v�t����g�$����`�>fS���TT�M��/���ԜB _K˓���'�*<�`F��cXv��Th
DD�ݵ]���Dil�]����Ml��<�W�O�!�B\��@�,��O����n�f�ړ<L�颹j �":G� �`��f2+1�7�V��-�F�w!��C��w\	�.�w_����T�K�w�*(�5�nw�AG�L���1�\�w�;����ךhb8JU@%�?�Z��r�f��y";�*�:�e����>�=Sc��C��b<�Y�@��nQ�vͭ��-E�<�]el���I���5�Q���$�^�?���C�hO�~� |��4����S�:�>_S�]*�P��չ|�e� �щߜe6| FOK��d�H[�g�-�h�"��xɹv$ʰ�Z�U
aӊ�	Z�\�~|L�Z�زC�g	�2����XݝW��ו�QSR8�1��)pE�͚�ǺA ł�_��'
�x|�?u
m�ĉ���k�v�L6��y«�l�m�=�i��R�b����P��'�hx�V���j��
���nO��E��w)��ZV���t*<�"�]���`��O���7�b���#	^W��M�@�T=:U� m5��I�5*={&k���/ƹ�%���)�t�0�ǯ�܎�m(o�<����:��˳?7�3�+ga����'�+���� 9C����Al���a#"=xB�CM97i�QP�q����8��@�`��`�@-�8͈�0G{��Vi8���e�4��/BO�������<rQ�T�[<�l�� 1P�QS������12�����$ �2�L�*�=d�y.Z���ӇD�B)TF����)��˒?Z�s��rm�ǾC�05{|�o-�������v���8��뇓n��F���u�P`-x�n=�y�T���݉!w�^��7�}Lk]X�6��.���?�F[4)Ի�W,�ɛ����",Ϫ�q��PE��mú(�W0�F�滢�~�[u�0E��͊u�=08��j�Z�h�H���.�V0�n�}z��d������x@��+�@Ff~J�2��8�,�EI��!N0te����)/�*�p�܏�X'~8J�$Be����6������m�Bg���a+g+�<0q �}�@�o���J�@]H\�f��̨�7��tx,�R�#:2ެ=tw_B6/0�J�>j�_�k����XԹ7��Q�R AoJ�{���iȾ�="��B�0}6�K�C_�Cq���:���	�e����quEY��pt7�ǉ���'���c���fl����7�&!}w^�<Et��ʙ)��,?|�2��Ŧ�_)ꨜ��� Z����������V��.��	s��_��\/���	F��s�w�[�#ǘI�6��b��l`�cY�|=�ڐG�#�z�m��]�
*J��	"/�2u��]�2ƺ��+Ϊ���#'���9����șD��ڦ�;�������Բ�$�Ld~��f���3YZ��8���ܥ��b�G=��/�)�3���#�t���F:Դ����)E���p�%�Z���j��'")�/M��A �������!Q
W>����0��.̙
;��Ʌ@w��hk����,:q�^�ͤ��e����Y����@�l�S�����<�-X�˫��fq���p�T0�����4�-:���b��+�iW6WԀ��L�3�bBHa���0�hY��C鑭f�d�܏?�V��P$zf�W�)X��F�|}�rdg0��x��|����!����F��w1Qg#tcdq�ͯ��Tut��[uՀ�{��H�S��V��IN�C����3V�Fj��0�k�^�ꎺ�:��/�G��Y��-�O�j�XQ��!3!n^#��~^'P���k��� ��@7[��ܒoF��g������_� �ˊ󁵤B� Yۥ�M+���U���� ����n%�x�#q�{n����g��ә���X{T� �@+��@��#�Ӭ/�rm��!�w���-�I���������SW@E�  ^�lc��h�+�p�D˿[�#��L�,��u20���tA=y���F��	�&���τ ��`.��(h���Țph��U�e����%��˝9�<_Я? TPÐ�
	E���0�TU0+[zmۈ���O��I������;�oE+A���BG�"�}��a������C$��!���Q] ��hM�w��]_f]~���fsv�V�����.8��� ��:�}$��Ω��[�|B)s��M��+H<p���9�b�P"���R�=ANj�6~�MBƠZ�~G-��Z>�uؓ��n��dR�k��T�&�69Yto"�8�Nn�TD�s|��\j�CzZִC�Q�^��(�,dOdA�	6�2�C��'.�i�<���N��f�-�\�� ��%p������{x�ډ��G��%:c1'��2֎w\q��N���S�T]����ގQȴ�Ψ G���E�7���d ���,[+q8D��a���	7|���~䓙��P�B"&���E��n��U�����CϢ���(���6�I)���-bK�v��1y7�Q�����J�l� �$�Gc)�}���(
��9�[�D�/A���!��0�˞{T����l����SG!�W���Ġ�_��ѹ�W�f��V��҇�����}t@Vw3jfgߩ�U��B"�6�.D`��'8zX~% �os�7n��eЂ�3݉GJ����z�M���1&3뢋�o2%�(,�Pf���$�bKɜ�����P(mMH�TB��o����Q�����H� ��ْ������v5�s n���LqlͲ7�mdN���EeC;')`?�t(_�x{�u�h��FN�� �~�T%cB?�,�6b�I�k{~��[�����i �/6��辘�������=��P���bi�9�Y7?\Czv��ؘԸ�����M&x'��q�G�|�ꑇ�}~��I�BSZ�eg�=��9�WOu+&�h�&d�r��F̔T9*��%���Y�6���=��Lv��*�P1^k�"0�R�8� �q��$��d���w8�ep�"�@r]P깜�H����t���*"�_�^1���5�k]���R��tO]�k�g�5��>=ra8�<�[	x건�G|H�0 ��������ꘅBgyrp�f"�{7{s�0��uA�ɶOCH��J�����0�e��&l<~�D*��C�u�H�ng��.����h��xF2F��>�)(64�"<�u\��اYw�e����iշ��&�>�����D����%��GҶ�x3�������Ƥ�b��m��ٙI)��RP�j�������~IJ�r�K����G��TyH9��� m��X
��i>��q�UP�֣�D ґ��-�J����l�b�;�sa�@H�Ü� X�RP��?
�|���m�l>"��J���5��ꐗ�r Z2���b=y	�%�>��t�Y�!�|(��>t%(iU2�z-�kyUZ ��(3�v�� rp��l�z3��^�ʊ�G�!*�W��`P=��cI�[�����/����wO�$ xO@q�׏s�y���A ���c�){��)S�#��*,5G��^�^P >�jӭ?E�)A���A|7�����zx�����&����ҽ-��~j���+l@�nXL�w^^�r,�����o�~W _N�־򍸸�k�j�EkG��lP#�6]�sI������dr`pSZ��d���i9����-�q�P�T(���?��0c�����"�����Q_,���^�:��h�3�?�i��'{������(�����$d�E���U�<n�b�"�������H.j� \#�A���L�F{Щ:z�*p� Y:d�K߷��qLۡ�g��7Y��u�67�����7��u{F�[����к&�"���K$@K�2ⲃD}�TͰ%��g���\J�I{������PS�;���w?-K��e*C@���4l�K��r��٩�g��H�s�_�:�����L�K�� ���ǖI�RR��m{�3��4`�^��tX61.�� /,?L��՞+ӭ��06��i���?���ZD�yA�ޯ7���S9����*�d9�Ҋ mȪ�o�����,�\v��rv�2t������?�^�ɾp�G�Fv+ �sS]���/ҷ�DGü����}��f�7�G�δ���:�ķ��ٸc�)(1�&ݠ��z�-���	�+�(���;��e�pE�o���9�t��O�O�ϙ��:���5l��=����M���(A����l����7k|s�qb�*~���m;���M�����"���[�v��M?�\�"���J��>���W���5�?SuO�?�mO/V�Hc����S���j6���IH���7�w
P+%�C4�.�����}��.�:�l��'�C0��-��P�%(��)���jS�iɟ9E�M��#Hx��i��-=�	*ڐW`�P6�F/ao���k?�R���X�� ���cW5�bo���\Z҃�F(�l+od��)��ET���y���� i����,���e��/&� �:���ѕ$�NV�תf�w�Dq�'�]����u�����n}:w?��J��>*#bFwB`���sj0��aN1�m���8�ON�-;ow=j�Z\'�%_�F�A����j�2��"x}{X�Z4��'^0��CfW�PXk�M������]��GgU����Z�}�ޏ۔�`��۟x��^B���]���8n1=I�2	�W��Jŝ��̺�/���7I���+�k�2*�7�m`h��e�C��z��@q�����Lg*��*6dL*$��ٌ|�pG��C� Ռǆ�P"��d���m��;d�Epa�r��}i�4%�Ftx������Q��`�/n�n���U���f��t��j��u� M��������-���Qח0���� ��?O�G�Y�IL�AJ@	pn�gaud�MX�,p�=�>F�:-��ᶻԣ��\C����6J��6�.�˫T;��%:0��6��Q�-P��%�S>zj{=\�Q���nC�j��ӳKi�8^��8	N.%ypeuاO�%�w�YiB��7|�1�#�5D**��e8G9�D�BŶ�N�ܓ�p���_kg�}٤f�����P���j����V,�� �𲿾��A�x�c���Ȳr���ˍo�N>J�%p��o��J�u{Q��Bő*W�rT���\%��v���:u�~��˼0�J�;Y��H��sVG�1����L�jf� �v�q�RJ�Cp��Z��rcy\5N���F!<�`��y�^::���y�6��}�*�S����K�1..,G�'�<t;�|0�v�n#O���R貦�k\s~�Y_-H-�FOa��y�r7�J��[�o�:�]ە63�=$O(�~�W��@���I�[�۫\�P�<�XO� S�rP�6�F�{� Dx ���B/��J�~bVDW��h�ߨտ'�;�T#fZX5����ԅ�a6���v����!�	���%#4�R2HR�a惇JY��q�r�&�����6�����ና=k����=��@f��.��x�� Mš��P����C��.t�C��r���CI,�쨆�U��������oF5��:h)�!$��~�fP�e�Ąb�hFGiiXq�2��o�������yz�������1���Zk{0���ET@����J��E�s�g��[PM}�@'�Oem�#80Eקr�����Hp� ��{�\W]�'o�ͽr��
e_�?�DIB�ׇDoL�_)����M�a���i���H^w��F=s&�>�'�+�M�X *��Vi�1S<��cTNq\��VVǏ��m�-������e����*�:f��3����i�;�B�X�U�I�/�O:����BP*	�s���-�d�$*��%����G�P@�׈��	�A���f����Y�v��"�H��� �R����F��a��P�� 7����yS��ol���_"\TC�]��o�k����˦e�=⪑�'pt���������}�]:}�̀�I������=8I��c��a{���I�3���t��a�<!&����:��끲�|>��WV("'��#�8�H؉T� ��ۅv<�G}!;Gx��繅���� l	L�� vj�b���c����iL�[E��v�a# ��;n�c��� �([��%wœ���P�O$�	��#�.H��C
iZx��d�ĵG.�c�H5����������N��Q+�ЊT����6.��sc���-��Y.�N��DY�T��� &`?���ye����$��-Oe�MA�����N�L����11Ȧ�`t�ʠ��}��a	_N��)�֨���G'���Fm��2i�կ���m����:c�1�Y�]�0"�v�,���K��a�e5�ڃ2,��g�8�X�O�mb�I�7������ϝ�r�y_8G��F��qd4{�p��嶿+�@�^`�Q�'�6����Չ��],��o��;Fv���G���=���ī�'���gǜ��p�pl�%b�T�*���,U�E#"A�-(�`�K�g������^/�4��$�?�C����1R��X�}�PH[�yD��� R�'`�nxق"����qID�m���?�rzxw�Ŝ�s��}��8�\;o[>�kw��� ��Z�Z|��!�A�"m/���5��H2>ij��;�������~$-M�����N�WkK8Լq���ڰ����!5I#O�#O�ӦX����')8Olv  ����/�C�����l^��~N�M��<�VIg��� r��ژ�����1��4c!RfgUs�Od��q��2#<�{���g�K�Jպ��6�:_Vk��C[!�і�:��ԁ�gv��D�j�$�\y"=�w](�vz![���� H�����x��6����I*?�sG)5�����l:BB����-$᳢֎t3G�V��[9 U���!�ABIV	H��W�J��i�`�3�bop�7 z�h.& G��+�b��Zʼ����%Nͭ!�@�z��5S}`]���/cP����=���	��Lc��q�A��L��`���Va��>\-�`���A-�&0@�~)��{ 
�8]�v��dbɺh �+�������
�N��S�������Q��b~-�( C��i�ͻ�=�3��7{V�sD��}_v��(-n��Y�XZ6"`�
���A5�9�Ϫ��6;��?��8��X�>�9D�㶉r���h���8t��uM|�ɣ:b"@E��m@v�'��(���<����1�z|��oB�"y��p3�ocF��W����S��D�p�U&�8�U(�T���5��W�`G��@1�-�qq��x�����G���1y��yV��!���4LlB(Wl%���W���K�7R�k  \����`���ng6���&!ǳ��~�pu�����dL�/Sg��������8��R�����e*o#�ޢ��L��fڋ��}Pm�� k����;A�E�iz��O8ڠ��s�4��k�C�-~Y�Ϲ�]����hϮ�TA�9���af!�S��<�=9W6&	(�lw�6�b�B����7õ&l��,�������[���1�t�����b�̦s@�|��:z�wՐ�҉q�dB�l�e�j4K�#��K�.F�Mu�c�	���?e�xҞ�~��6�O9�y��đH(����$�.��-��Lӛ���V�.�Ͽ����|E�^F��Ɲ�l�U-���傊Zş<2%HF��m����R�`�@�!%l :��+%\�D�9t�F�L�Z��%��σӴT�h�BD�	~s�W�D3��u:��ޮ!�&����b���2ZY�K��Mz_:�_)�ZBl;8$��;�-O:\H3�_H.�v$�e+D�6GK�X㐏��gp��V�E����Gv��{���hF�^�ͫ֡��z{5M;�A����R��m��x'њ|e!�`I�В߇�j��=��=4�4:�()㪎f����1��AM+Ö}d��' ��'����BG��y�������йR��R�;�?l�!��(�5�!�/4�Mq35����H����`�I�C!��{�$U"�`�9�����[S41Y�����*q���t�pL�+�)��{0u�p�g�3(:v��J���|W��r=Nr�yf�kd�i���������v�p�� ��Z�G�l��4�;��Y�������4O�
bί+\Q�ھh.�B��{�h�|���v���6W8�y�n�U/��:���k�妒g�!Z�)���*S�{�f�9@8l�C���E"f�CЭ�K���w��w���B��+�Vob)�ב��ѤL/��;&�xݭ�~��K
�JWW�x6��C�K:b`�pN�B���'�Ғ�\bokV�\�.��a7��w|�mQZ��t�5�����CL�r���pO����z�C�� ~ߜ�7j���ό"��7��Gt��?�(�ʨ�R�E�RB��9Q��Z1zu/��@�#�ݵ����V}�<�c�n���}��*�M\A�MuEq{�	׸5���as�/�gN�׿��Y2O�3�UK��5>rߺ�c��o�3��lIؤ���l��PCI��ͲB�?�Q������U�\q�w��h
���I��Gy��hn���F<ש}勨��Y_1T�w��]�+ʲS��E>� 	!�b��<�$�yQ�"�P�E���%��z<��SfK.��Xe(9�Jx�/�㴭���|���/�d�r����s�8��8sp(�Ʌ��4l*�v���f�8`�y���XAQ�ݗ�c���ǩ������:\��z?��� ��|����[�8�f�(�mO��D8||9U\��g�+v	��yq}��aw�S���U�^��t���[�HHm�J�b���Z���z������gbSs�T�
����Wx���2�d���a���Y�/���ؾ\��@>��n�DV���f�q!ʉy������i��ٷ�R�����*�Ԫ����EFO}HJ��`O�m\u'_8\t����i��i�z��8Ӄ��^!=rpV�8@8� Q6��I�}4��Q�q]�-��Y���n����c�-zu��Db	5��"�3ZVF�t�Ʌ�腄����F'��zz�9d���1��L]�ӻV<<R�nOzZ��F�6(�n��Yv�y�R�[)k��&oU��׉n�����9\<U�o�z#�!%�%�moiG(���V��}�H'��
P����#<,]�}/T����x�͏V;RK��k���_���˪?�#	Ui�S����#�>d�i|������k˓� ܓ�6b�E�T|�����5�/�����D���	�O���PRS�y�����r�M���=�oN����#Yp��G)�#sYC���i�y�������!��Ss�n$�5G�(������d�q(9r�혆�����L��uI�=��H78;N#�
��Fܶ[-�J�a�J��y��E�B���b+*�ݦ�Ǹ �~����:��E	^�ak��왺��(q����O"�+O�!(����>�J�J�:��'�;�b��5_�����z����X?��G4�4�^
��y<��H��F��k�$��̃�����i6sZY����D^��vv���1)��h2\qۧ��.� g�6(�.���9+�ޅ��p~�"W�k��5,A8s���!����Lt���"�};PzSJ��߲��Ϭk�A�뭘G�7�@{�(�!��IZ}k;!�6)�vþTm6\^˂��vm��t���䷸�鯬�k3M�X��B5`{{���9���`%�:�oe��Y���v�$K4 �6-��r$O=���.�Xa�z%)=
 "
&�۽A'M
�#�xP,�Z&V��8\h�$��:�Ԓo.=x
r!z�4/gݺ
�%dyjT�(���
}�]���Hq@�X�+5��>?ꭾьP�TIu�z��R`e�`��綿�� z��1U���5B":H̆ �{�����݈�T�լ	Ҽg��F��3��E��bz`=.T��g��_�����
~\K��0@��㴖�\�c�K!���ȑ�dp!�����lZ�AL�&��8B�nu�L�퉷��H��I^�g�:z�4	�BXn�IT֛�#��7 �f�Y�`��BV<�x°C�=>�4 ���^������!}?TB��\C��E]�޾�2�D�SWAm����N��{�R}Í'�@�_m��*����ݜ�H�P��9�K���-�R�{l̕�F�q�֤o�&�(�[���<�r*���/�����zMG*5�'�ňV��J�D�������~�p�N��z����ݬ�~�N^��*���������kg�Ze����5˨�S�x�¼���t ���~����"�K�J�1˱zHD�x���@�N�J�/��9Mx�}r:k��˚g�=�'�t�-���L.ߗ$l��,1��/�q���O6xpsv�B��(� ���藈+xzp�E͏$Py&Dc���������3&v[5�o�� �v}�OS�0��i��\!��?	�������d�L�s�v�>�\NxHȕ�<{�/RZ�h�V	�USACƽ�R�u����~��0�=�Mc�"��?4�� o� �̰�)��r�_D��p?�˼���|�������(�4I\V�\f��tH��<on��"ξ�+�� ��PM�DT��۝&h㍓�ө�c���2=k~����vU�����U��7�=B�;\R��k
�9.4������ğ��z�8��SV�iGڎUu7v]V�V"����r���r*ߧ�ʩ��Y�]��j�.F���~��:���[�hlEd"��4�H�6�փ��5�[��>P���*�5!q�_H�b-�%L�e*㈝oX��
�t���A,`&�u���Exk��"S�q��ͽ\o�l�L~���OA��73��g�
H���b>�=������K*q)h��7a4�i�F����~��;�:�(�N�%L�q��h/��(�%M7�������a���!5�x�4#믦�2��!�L�PwJi�/&�p�CvV����;��
��\e8�!I�x=�Y�ا0|`�-2���c�w9��� F���kZ�s@T��a;�v��Q'S�}B���տ"k֪z:xֈ��[K�Y�Ԉ�[�=�x�*���f�"]��3sNN}?��73�Z�X#���#u�&O���Z���ÊH�� ���&��.�<����V�<(�v�$���2Z~D��t�Ѱ�-�*g)��������_3�=���$��o��e<�U_c�RK���+Ƕ�+�&��WRnGOEE�:�1�k~+l�n$|���x�"�!��J���c��Q7�G���{v
Ӆ.��boΌȷ���qG��c�|ZMq��ŜFt���p`/�ls��T���M�w �u'��G�6�֔&�,teCD��4\P���B.A���Rpc���	6���0,�M1j�	�Zd*���0�/XG���tfє���m-*B��~�35=�w��4E?��æ}A��q/�3��yBx� ��h���ժ@F�w 26q����;�'�1\Ť6f�X��h�ҞE�7��-Q�PH� d�~C�?B��'�a�;�����$�+�dj4��D5�M�ˏ`F��)����ٱ�|<����uZ���w�p[R�p-��X�|�5��eR��q�3�u��:Z_��l�[�g��zA���GC�{�Wȅa��d���O�e�@j�f/C `��q��$��	���r��Dr�\F"�@����:�&�lWD�� �.�Y�V�_��9��i�N��I�����?�pZ��^8&޶�p�s��6{��RN1�ܫG�c	"⨌C�o͖��f�M���h���q}-(�`5}SNR ����Ԇ�5o�ݙ�i���a���]Vq�;glL&+�a�uP;k������go���8a��gE �!���>$�i�JB�9=���'�C��2h�%�M+�Ա���)�jw�Y���*(�&y5�p$s^�/��Iv[,�������\X��N}/�/��̂X5��jV��RTCW-��2`�ELmU2?�2�pm�P�;��}�w�=�5g�,x�0#�	�u��-������c�k��F��_o20p��(�+�1r�`E)ӡ�o,\�)�c
 �n�i����U{j�ծ�+��FB�l��枲�4�_U����F?g�l;eDjI�+U���	�w����Wd�S�F��I/|��LA2�[� �4(޽p��X�NӨ���}m�����k�0�U�-3�
ď?-���dj�]�|���T��x�E�����\2]��11=�FC%]E��W6�վ~�Խ��4G�s��ӈ_� �� *�첅�:C4g��ʴ�n�k�x#�y��ک�K���]�.cv��!��3�u,�(](X=l&%�50 ��t֙0�^=Cc	�t^�Xe����c�:�
6Z�썎��x=��u���xx�V�qvP|�����x3�%aB}���O+�����{�����r�^ۥjy��ژx�N�t�)�w��:Z���Z橫Me��7��U��S
æD�6��`_Xny����]�E�q�A��>�Xm���TDT���t�@Ѡ����}!t���i�Z_���z����U��!w�=��%���z��_ M�5s+`�r�cLX+��������Q��:�t~D�GT���<�G0ɋ���T��8�����W�f� �t��Ɍ�6� NJ�Q���)��eڊ;�,�Y��a�yn����$��ƍ6�͑З]#6�x�gn.��.���G��_9������4�%�w�.<EY[��rfm�9{��k���ג�\�u�
�>j�W�YC���N\�ű��uD��,��{�c�֊5r[�f�I,��޻E�<#�\�O
�Ӕ;X�O��&�m�vx'�H�;�l�� E*��f�B�2{�g�~�.e2Gu�Yp���C�<��`��wm��2�@�L�$*Lc���T6�Lvf�0#<�l��<,�G3�#!�Lq�ӱ����Ҳ��	���p�۱%�܈v���!;p;�4:>Yx[�6Bj:�F���xifK���9���Xl�s*�RY���L�� G4��!�8zL�8�Fs�9]�E�<�`�b���:�d��,�@4����?�H��D��o`ϪY�������udj��DQۦ��r���7��)\^8�3~��Am�:J�sΧR��2 ��k����+AF�� Q�y��t��T��BN���ȗ��7���g�K|�NM���
�hx����cu�ݻ_-@)���	��(~�
Q�3�S>��O�����"^^�v(@-��1���d<Dx�}��7�$t!�G5堇�ekG��:�9��TRn(��:��_ѥ�h�D&�����Ʃ�h�Ns��.�4Y��4@[&���I�tR���NƮ��JDf��Rrd)�76��d�ꪷ��.^s6:��Tۏ}o·�����9�g�0���}}󗨄�J���s��nRt��#�g((�� ����M�H�I�2�=p���J?_d&�%٘{Dw�v?�~�t�9����M]I�x��Ǘ�|l��.w�x���f'OUn[]e�K7�Sm��#�)ҟ�w��z�n�X�D���	�9���.�wF�:%a�\$M�/�,x��n��q�2s܇AeK�^�d�z�#^�V	Rm	����hb{����d��0�|���jD�Y��`����ZI�k���B`�N���h�'~jVX��sK|�KWV��T���R��_?:�}�_]	o�S)>.�K�n��.b&�o�b�ju'@u��{��NG.�� ƆI����M��2כ��@�,��m(�%�r��VG���$��j���9V Y ��2{:ϣ
Ā�P�}缿�?��9��G����S%�!��>�<�i���~Ī ���P�o"^C͕��n��|uo�����7��|�f���s:�1U��z�3K�8�B�����/4F��
�-*vxD�e�ʄ�H�sh�#(X���=��<����9�'�"���~�>n�\��F�%�ι_�L{�MX�#/BF�47B����d�F�������>�ޞ�h�>�4��T�R�3����k4'>z�f	;�zY�N4~��X Pߴ��+M���Q>F �ٽ>W���F!�b�@�+Mp����dn���s{�h>�6>�O�	.-�\�U��k��Mؘ�3�@���r�+��L0e�d��S~%)Tu�k��{LF_1�Xn"����K;wt 9��[	����]����҉PX�4�rE��G*F÷(_�����D�P��m+h���y��!+��&G�m�3!T9��*��S���8���J���ӡ�?M, ���U�H�q�#�)LN�q�2����d���s5�f���7��#j���V�������o����Bk'�u��y5y���z�[i��m6%zc}6��aa_v&��+Fi&���.�����������S�̀WS���ċ�Ʊ���ц�f���rL?/N����;`��.�q�èpn�}F�eW�g��[��b�-�����f�� }�і�u�>�����h-�tPU0��j>Ǵxi�2i�H�^n�}���_�rFҳݐB�X�����{i�H�n�*�����D����ݘ<PO��)$�uv�ʆm޳~/����"�d�|��B��Md�Ln*a�އ������C���T�?y�G��Q��H� �Tk��4^D0��o$�>�k�i�oEʔLl�౷�~�,s��ϡ�D4�~M{�w������N��.���E&�:]=wS�wg�Pg��M�U��9a������Z�\½T�4�%J�Z���h��6C��"y�Î��9��o�� ��+�.qx:<8�O�d������e�=R� �f0�n���oI�g՚�!�VE�m�P~<����v�7f�x	�|��jbI UF�0D2	�b\<������#��,���Ձ{|�0y4Ӷab�%���������W���ٌ��`�W�M��H�X�[��@X� �!��)�R��9�m� �ai]�hl��1�h���dI�@��o�C��h��W�ML�Z�^H�W~ �؋�K�5��R%RzK��V���]Ɨ̾?I�~�]x����2Te'��~�����\Y�x����
���6آ�R��*��s��C�G}1��D r��F��'Y��F�L������y�՟ba�Oa�� #�z��^/O,C(��kB���������b ������LS����6�J�o����-������9ϖW����&i��Ǳy��n��O����a3{���hU�Ò���u��@:+�R�g��{lbmqH�*�e�Ɵ��<��d�ҧv�K%����&�<��;���$-1�`1�M6,uL���5(��]��n�/_���o<^��nF�tY����#9��՝r��|�Ej8㽏��Q�i%Jc�B����)��V����v���0 ����
��� >5�5m����#P�]Ig�a�������z���j��4=��i��J(Wj�\�A���S�"�`�V�օn �tp�5uǟ=R9�="C�����T�<g	���>*rm@�R��	M�2�L�$!����Ȟ[��f�nw��Ore����E�O���r4Q	�tʣ��,u���"��ߡ�]��|#�+���6G����?��n��m��x� Y� �����!M*̠M"$��V��u�8�6h�M�fY����_;2�@�G�O�����[�;:�\d������*9��� l���`X��Q�[�w���v��dï&-�
�r;�)#	�\���pl%��0�c����-��:h��p�{	����%����S +�\w�$���&�^���j���	�9������ȳ�������(�[��۟^+q[��c�+���ֆ�6���~ֽ�}�՟L�����J�Iڬ}!V���^��⾫f�cw���V�'��v�sP�{����*�懱a��Up��w}��X���쳏n� )��E{�g���s�l�3��R��� +�13!���k�&p���X��r-��h(�VeA��	��(f.�;O2�~���N���gl�|���-����� (��=e��oi�j�5�1-��0�S;��PF����	6�U�:��&��f�C?P�!��\1��]]��33��2��M�s.4�$�$n�q�=�ܷ0AG=n0H�g�PzQ��lZ��e�{\�F�lӚHǲ��_#;�M��&�6��H��4tQ�k���{i�bk?*,%`�%�H��3ݛC(�>q휌�����_<�wv�#Lv�&�Ja���ׇ�9/�z���2��T#P�����#��ə��DN1lzv�'��+e:�]���^�^g���-J��J����i:�������>R��~�r�'�^l��]�짶�B룭�|���U�J��ܱ|�>Ϛ�e�c����C�M�dw�c-޵F��&Mo�Ʃ~n��;n�mV71��o-X{^�`csD<Fw.�ي���4��mZ��.T:K)����nQWbI����t�يL�{�KH̪�S=lih����iU��Ѝ�I;�hf>Ѥ�(MdN z�I��������Ɍ�}[�z���Å)�K𲏯����%<9>�tȎԩt̂�{#�3�����~�q��DԔ}��O��sTe<����so��_���ص�q��4�7��=×^H�o�I+7��t�3��E*x@��إp�qe��$/w%n�g��:���?&w7��Ș�O��E��1�H�y�J�S�2-�c�뭶?����A4,��\�/Z���dZHΚ��=�䡛H��f@��➎{�����g��l�������@X>W�vT��u��
R�y �N��X͑SC�w���0.�΢��7 �8O��JEQ>5�+9�A��9��8���=B�A��c �[P �#*b�=�[ ?����7���e�;{��K�q2���%��̄���ykW ����e�7�MD�����9]ZFR�Fo�k*S�'O�yxZ1�,T���ߊ*2�%ױˢ=l����$���e���:E  ��
�9`��6�$X�^�ӐN ������TENj$\)j
�O�pgo�2�md�W	8�0��ԇ�s!������P�r���(\BO[M�#��i1�:0���������[R@��eĴ�=�x����5��K�!#���	[��$��ʧn�o���������C��)���3r	zx������������\�Ќ��L�0,�ȏ��e���}z�եg$ҹZ�`l-c��t�����0���_$31���[R�=6`��Z+z���g6��m�{�Y?9;)L��DCVi�p.ߟ">_C�7���,�>��� �?/�̰%ӡ�O��vR�(�L�/鍪^��t�z[�(և@�4�薑�kTE����AܻoPb�;��C=j��U8?�1;�עV��\��f�"�4��4$}�OY�'ĸC��nt91 ɵ�J*����&C#HY� ײ����p+Y+e14��AGo��f���}�ֻ���^b��ߦj�EOuCbҚ�S�\]����ɞM0T��L-��K�� H��y�U�c����ȱsŤmTՔ��7�?��f���/p//N�o��j�p���f��ʃ��9�-ķ���M���gܿ�7s���u��>`�F�
V��f��t��cp&/�z���f��\{���_�㗨v�P@��fnN�����`��@VYۭ��#�_���Y�:d��)�[.���nO�g��n���%}�&q�9��j��x�Oc\A��i;����������7 �r��_V�j��\=��Q��kP�Q�ۗ֞İ��,�l�2�k�i�}��m��O8�3�ɦL���T��!;���I��~�-� I���q`���#�q��a���� ��u�&�`@���F>H]�	�\,}�y��BAy�a����a؀0r'�NFRf�p��M������h��~���=��\]8�9&ݝ$�*��lV>h�F�A����@�S���A���BAf��$��s|�WlZ�២���e\`g=#^m��S���q��[F��愴i>]P"�8ͷ�>{tt�u;a4�"� m���:� ����;���g�?3無G��� ^׍(v��L�