��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����Mڨ��˳0��`q�M�'���2&��Ȯ�W�4��д��|�6�K!b�'mY�`��L����T9 �0��6CD�Ux>F�,-0�ZY���J_
�璥�x�>��xk�onb͂��`]��j� X[��c9E��&���r�4���W(R�E
,ݪ1W[e�ߺ4�a�t��2~�_]���>��(�RB�B^�d����AO��Bt��҇��+�l\�H�O�Gl��r�[=)�P�%�@���=ī�4����ȴ|�h���+��#\��VĄz�>�:3����T�����6���w�� ���LCC]'`�^���1�+�֬�4PΉO�����%�+7�}0�+"v>z؇�!E�����i|� �K��n��JC�H,ҝc����E9�s����F�W�Q������l���+V�șR4�^��#��5�o�5��[V��2��s��Y�&�]e.�|�N���&>F��G !N}(O�����>8i�cAL-J�ZL����G�n��o+���q+��2T�[5�6�����ߵ�ik:� ��7J�f�����K9�ku��<�"�
s�#��Ff��'��rg|I��m.�g�(�pB1Xy�M������0ܰÿu��e]@��㮏ly(�m�J��`�Ŝ�Re!b��hx<N`R�o6��M��Y�v��V�eR.�7W"fˀZľU�e��ݠaM*Oaއ>t��gB-�~|��!)X�|0R�P�~W�4�P�VQ�2a���V�V�瀍;z��G��z��S*����-�b�k��L����&M��\|��a�'���<�P8n��7�:����f�׬��&9�B;�I>u>�'a�o��]��4�)��Tg$����g&�_���)i���jKP/��3)��VE�1���F�9���+�oT7G�|����i�C��#��'��qb��)v�Z�YO#b�kmqJJg����?����]�.:��0�x ٦���.��nM=H��d�$ ���]�K+ĳ��>����${ � _�߮S�r��䂪� ���B8@��71��|������(��d}n�<bG�7u�:��[9�;����ɓc3����;FyF�hCˮ��Q��B!�!Q��h�dcB���Ӆ��QΗ1p�8:������k��3lՄ=o0�Q���{t��y�e9Π�P*r�<H�L#`�A~ÒT3F��L.���m�-#�P����K�Gu�s�g���C]fؕ�C�����/(u:�*rt�z��*hA�Vy���1oy�_�e� ���׼�����K$^�rl�ӞrXGφ�^�u�c��U��s(+����gq���F4.t��9�����ȴ�H�o��AO� �o޶2v��ʶ�[��䒥�bk�*��8��s� �b�Ru����ati@ڪuR'��u6��wv"��9|�/�hB�RH%��P�x{�o��r����LJA�'�����ʐ�sHDI	-�|��4�m�Xŵ�^�����D��Qr�+̇��SMq���HGX(_�Cq��a���u��	����e����y i5_੽�aNѦ�� L�F�I�^��m}��Q�%�gi^*D�2�JG�&/�����k(?�F��^��V�5���Q��1>[���/+Q�h}���2�e��.؈f�Tʼ��`�y���y����$f8������5�gc}��ǭ�T��o)@6;�^��R��?Q���]\�^��f�w������&5�e7f��U>%����_�����RdT���8"�'T˝0r��ox��e�ߛ�yOKF 5����b�@zR��
����p��x*6��� �&'Y�#���U/�`����tl�,/B#�6Ɯʪ��}5���J�xV�#Q�ز�P^���%ds �������N�R����EDG��������g���aó/gD9D�8��	�Ŕ'�;������/��xtx�O� �ҖfC����s�=LP
��o �
�9=��b��F
���!�1"�$���LBF���*y���[�I�s��#�\k��3�d���r	��������D����Q
!K˿M5U�{��r���iP������~4�6�+꙯C~À��Ǎ)��]�sp:U��wR� � �W���V��w�BEq�F��(�J��b�ٶ�ݐ0���	�9?���{��3$���TU"�Js/��SB���>J���J�l�D�_rM��)_U���n�H���+4�����*�^�ކ%�;� �~��r��M�!���ĕA��b9���5~\�$�X`|x����.���!�Շ�~���^�?vې�˃=2q���t��*Y.��H�8d4��*na���L&\�?@jA��N#T�8>�2�~��� �VvֹhvgW���6�!�ߔ4�t�D�Q�HwV�r�^�We��ee�)�����P7����{�K��8�@�����/��Nn>��)�-[��}DXWF}��Yn�����Z�R&�?�vvL���̓s�c�lT��Ǯ��(u�)\=�S,�ƋL:vym�*1�z{�v�y�ܩO	R�=V���r�7��:��Xg��o��M��)�O�Z����u�Ό�(���/Q�[R �Z�� �|\���Q���v��O�Á����TY�����1޴.��p�,���/��3'��8A�F4��'�1L��'�ފ�U$����ϩsS#_M4�a���;\g=Ki[S��v�ux%�ٰ!�q���9�qx����D��hs3C��Dp����\>��:�J�}o�@c��UD�4��0�t'J�q�&$=[o���%&u�O:P��
aT�0�B�p�x�'����F�۬9���Swn@�B_�V��fS(��v�1�c��Z�삅W⭀s������)c{�/*�O}e��<�� ר�G>�'�Fe�Z9I���,VH��h>=t8�Q$�f,�~8uڐ��K�r�^f�~Er�7[�,�
nm}���Y��)�@���}��Y�(��Z�r'�a-�GU�Kh�b|�U4�6e�cY�F��E�O&W{�t?�N��g���,��_l��EeEb�4��p��2ϧ� �y*޲j���i�(�����%� r�G���v$�����C*N��G��i���ƾP�q����E�g�OF���������~(�(�ַ�Rz`d��`�7I(�V���_p� (��T�d�:_�!��#hHQ�=foʱ�P�=�8B_0{Bx��VEv�&�8���@��r{#F��`6���蟛;�~>9��x��̣�Z��[/�G�Bω�
�\r8MI���H~��3��]��r�f���Dd�p�J'�H�'��1V:��EQ�ޘ�z$%N
���q�GAwAn"ps��7�E���2*�X������JwpDa�c��T+�u+����z�K��m�5���l�u*.�"��rATvr���)b��c����,�Ʋ�}���]E���_�6�}�CV���xڀh�m����5�d�������k7���)4@y���$>
�H��^����O�K+�/�N���ܚS�d��Z�gʤ1UQ�<F;̟���p�C�A�S�?}�9d���V�F]>�쐪�	7�C欣 �YU�(Q�Hu<g5���!�^�\���B�n��W�'#�J�B�)��W4+��G���{Sx��F��L�Ј�� 3�C��^�R{k+�ټ���4������o*M ���-9�(p�A?_�_@M��O���T�n��AU�����py�:�SK��nH8�Q�ET���`"�`hVg�!x4�:Oǲ�9@n�l-/�nE}��_ ����]*�X�!�APD�"H�J3ˈU|��\Sg>��2��W����v�13����f�hԺ!e��������Sg������)��0�,�P��}�K�d����Z_ҮSݐ�ei�"L{�@+Y��G�g�AEùg��=w��}��;���g	�<�Ӌp>'�T���ߏ��!ˊ��V��~�;�}��Ơ�X��w@��.�i�4WRM/�����T��0Ƈ�J&�W2�N��Y�J�e_Rx���F�����c�vH;�&-�y:P� �N��n����x��AK�'��+1d2^�Ô���普��_M��5�9���`�Y;�P�~�r�_BAw���/tZ����Ѣ�������頟�e��������_�)jf)S�Y��fr���8��41�� �Q������M<��������#�k � �b����l-��~��=���P������eV� ��o� �5�e	��V*o�so#@Sϕ�A�Wܙ���*��Bq�<��@�h�{��į��x:;��%`����f�ǉ;}b<�:<^so�9�A��aח�k�@��$�ǫ���)m�s�%��A�˒�� ��S<���U���� ��R�Z^�4��J7�H�x[ixg$cz�~,�{��e�oM��\] � ��>���"�������qsZ�����^����0T�����.�eIh{�'���܅w}�O�+���K8?"y���X/>���d苗�l*o�2ę��w���Sh�9�^�@A�-����̹��ـ��<M�\$F�v�O�=I�Z��oo�TPĉ1j��=����Ψ!>����r�ڢ?\�O��J��%.�R��ڦm��A�h�t�A)ޅ����#��%��XĂF<�?�������{�i�e��7�v���	^�\3r�.T���� ���S�Ί	�L8!hcL�&���׻�iE�G�:'�'Dz߱r�{P���'NT�>�?`�rSj"ē.c/�yG�ٍAA|Y-�"���W��*���s0]�{������f��"`1B6��_{��f�WFX^q��*:lL��O|���fP��B|��7

�%���|�]yGk��l�4�0�I�>%�V£��Y�(��[ۈ2���*	u�Bꕍ�
@�GҁrGM�kr�>6�����$k�����Qɵ'���.v9�"�需����J/|ᮤP��>�i�p�e�4J�,��YIc�ą&Q���/���#���1RH'�R�a����EE+��7T ���c�d�Zc���Ĉ*dǰ�G
��D)�\Xܤ���v�L�{��	?�n�D�D�9�zTQ%�i��?I{i��	Kie��ϼ���.��X?�)G��ȥ��n}���5�EN���	���]i�3m&�]:���C�G����KvZ�����p�(N�������@�H�E���.�
#�֨�E
�#1��Y@����%j2��.�P=	2�1�+)%7�h2$�`M���f(\�wdv�:�8�v�	���qO����w�5�[%(  rX�>Gs�c��B�D;��_ɉ	S�B�ǁ���2ī�u�\��LMM��ldPU����	ŷI���Q�dTՔ�0>��/s���z�=��x?�VC@�`o�#�R�3�;>�ڶ��楇4/�`"wEf�8�$+��\U F��^ؤ�^�@�;�Q�ɛ�E���������{L��6o-Z�0 �!HIaݠ[��њ:2�fu#��6v��q�ǆ�BK����e��B�AP�E&�,�{���8֯���^��,�o{\!>�9 i��ϗ���ξ�,�8ߨ+�֭�R{��;����n���(҂f}����������/�6t���7��r���,�V�@[�o?���NP��3S�,��=:�xk�#�����вZ��m��SQӘmP�/��'�.�S��0��񌃽�}���w��(��X������9�0�vЩ9����2��x�n�L9�j���Yl�Ҟ	�����S�=X��;F��q^��J-ԗ�'9Eb��KM6|/�k�,X�Y�k�A�9���H^&�ⳃ}8ǵ��-�	,=g�Gʱ����Z�B��@\�CŒ�b%��%�$��g7�:<XTYvT���3"&fg�U�2u'����ƍ+j��ೌ��(e%���1N�W҂�?=ֈ���mڦ[*�'���������$�ژ���P��F����}B��<�؏>�d8R�5��K'�S8Vo�]������GQ_t�\~7O�w��tꑡ��n՝���Vq�W�=1�狥�����{+M���+WTBq��f*���	Ԯ��>��݈�T"�@�(��	�"�a���否in�B�G��4�0��鰸����A����Q�{T^Ӊ}kH5�'邘����_!����d�׏v���i��%7%��>���*��(��\2�Z~