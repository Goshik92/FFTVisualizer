��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|n�\&���X���S��p��0���靻��2]��^a��C}����{�dHjq�9o����2�l���n������P�-���jOpg�k]��[�h���P�u�	ӂN{I@ :(�L^8��	S������H%�q���Q�Q�,��9�ԫBL�V�({8o'ב��\*�L"q�"U)�~="��J��q���6��+c����h���G�1߬�������dK�`bߺT�a���D��֝�)4ɹ��/�k�NR�:{�w�OkM���ax�����'yyK)`��x����Tz��n�?I����2��zJW[��'�j��o7����k��:o%�0��cs�"����f�+u��㟸iޭ���kBB.܆;Q/sRy)�H��V�h��nZ����az&oT��`$9a�
2<�l �Z�z�h�+�QάJ���C���X�z��q. z(Ӣ���� b��n�K���o�{�0� ��� ~�ծ���	�.˞�	h��+e��͡�i���m7������3��q��1�i��u�݋(����-m�53��w�4Q.zY~�8*m��q�E�$�w�{����+��:��p�p�f�^���"�ѕ`~�Gbe@��!_�`�N'�"�k��AJ�3F�XgEy���s��J&>S�M����򆋖p����6�o}5��ro;��F�#w��E�%1�+D�γ��5�@=��v����}\,�uز*�Z��_�X��jd�/`)S\�-��Fs1j l`�����,/���z^���+jc*8?z2 ��,�<-fxE����	��6!;�� ���ҁ��Izs��4d�jNt�^��\c�	�<�ad��OG	�^���y�����j��g�����weSsfS�|�k��I$$#���N��,3締 +:�E��7����D,�j0��o�F�,�u�}�ޯ�Pѽ(�Y�x�k| �%�Ǽ�fA=� [�_*O��Z��:��r��bU�
$"��Q|��O8�H��3�{��Um�О��%��hpJ�w�Ω�V���ǯ�i/J�� �2���Sx�
@�ػ��=H�
m��ϸ�8=S���«h���ı�K�����<�7�(�-�ʧ�x3��5��3h4�<�<�S�eb�x�ETOG��[U�j��(=�ǩ|ۧ��K�jQ��\�p������!1��;��������]%��^�_���֙
�>[Zf�/��!��]�c�\}2ఐ뇤���n�������ƾ&�Y�#��=m��3R2�y��
�.ӞNO�Ⱦ/[��+_����l�{���v��1����ըjCsRw@~+Z�!��Y7ic\��\��m�^�
m��8�q_a���j��lDM��F�2�[�l2��m��#YY�Z�cT���j��i�1��X�2@��Ȏ�2�a:Fd�֢8%�6q��9 s��jP4U5z>	Ơ��K�i{>�s
e��X_�J�{yip�QMuP�;����1�w��u}�Ϻt��r+�x^J]3�(��HV�8��9�z6���İ�	�$�6�����U2٩U( 0:�9^v��<����i��¾����M�ta�ߤZ���}�i֓?�����i0a�X��g��xnB,ƴq���AX5�d�ֶ@L"&�j���(ɻC{1�Q*�;�fvh*��D*���@"^$��|�ܾ�(��z�?���A�7��P����ٯ�Lim��N�f���g�?�í�Y�M�쬊Z�W�t$��<���.Z��[�V�*s�\Q@8������r�h��`
�����u�h%��0�ā�נW�K���8�fzb��|���
~`�=���ۄ\�}�>���H4��<е�(%��*�F�iܰ`��
?!<�Xa��8U�ϨE�(nbW[��������Wb(��y��]&�R\ ����䣖�c���
�ڢ�d gl���B"觃�7x��nw�-�f�t&'����"��R�2xK�\��� U�
�a��	ht���O��C�7rX9o���t{I�r՚�h�$�k�nc �D��K��OW��o���NfIg���C�ҟ��}�&�ё�J��sl*	�,E�@|n�q���Z���5���m�tU���N^}��ӭ�͜�*�Pց��m}H;�\�<���Цd%�/�=2���,5ĀB8��y��4��-�[�r;�+\�"�R���%�`�#"��")4ΩϲdO�j�Ojlv�՗�4ef}^�Ck�8=� ��(���Kv}�]]��7y��"��Sӧ�_Q��<����o*��~�%��H������lчg- �~��5P5�v��"-n�e��^B	��iD,��~K�����P�( �{�7�֡�/fް$�ɨ~�W���s�)a�Jn\#��$�t������GN�L�d��:�A�2�³�=|�PJ�<��<��׻�V�L�U$�H.�OK�0% ݅}��qG;�
����Y�J&ԹF4�q����$환�w��Z��E%"B;i�7}��#*��wN���:�#�Y���1[3��S~}cn�=����J�Z3�������t�O�!�>�K���sR�����L���rr��<�6�LQ�o웢��_�����hɎ[v��mAV<sE��\a,�!��	8Vu����>P��rMP�r.��A����$�ZC���LtQ?�JF&�`���K��H@���Y���8�\���{�D��w�x�N�Z����>����At��_��31��\bq�$,}g��R�^Ϧz�i8���&�X!��0m��B���=��[8tØE�|/��b�3Cz���`Z���\{�'�h�������kJ�?��j��۾JS�Y��o{�O����������P&䞝��i$���Z�Ƥyq��E�V} ;0�i�qT2Q r���+8[����H�H����=���!$�a.���e�v�SB�w�L,��8���W��}��j�����p?_���=�Prr�8���m�o­q�
�al��r�u<ַK��Ky�u3�9���-���"F��aZ@@ "R��@�J$܎�9�"x�K79����e��?䲚�6>�]��:H���L��~n�)�*1�����u�,��c��{Is��p�d��ܛx� ;��6�6�{B#��ҞJ�-�H�5�Q/���e�p���I��x&S�|i3{f[�m�qw�&�����G�z!0l*?!�Sh�3..OI{յ�b�]�%[8v����P|�ΔAe����u�T��B%n�CQ �9O*���[9I���Q?C�O�݌�	i�E���F���^߫�\6�vI�����>U`�{X�����"��>mpGZ�W�?Ԁ����!���%��JГ����=��=�ܵ:^���
�+n�]�}/� Sw�tI.n<�zo	F� �ׄTk��R�p��c��k�Y����o�5^��*��L�qo�ʠ�s�d>`��S.
,����h�EJk6�|�N�ML������ӲIvW2��j/���eR���[�{(��6���u��x���׿R�u���C��d��&[�����7ig�����b�qB,�ldv\�v�0��@`qlYE"��֑�b~ܼA�"4q6�CQm%��������r�QX�E�R��'ou�6`�^�xFe�.���q�:IP:�,L/�"JY�����狈�h�WI��L�4P����˕������: ����z���c�j��ffj.��À���Ā L1�?3���eF����� `���+��/*!����"�P��{�����_\�����1[��O].��]:y�D�M��8cps�F��)�aC3Ba�O�i:жOs�t�m�������%����7����`�=����e\�To�:�Ja��T]��?S��1բ:�1Q����^zM�w���o^��T�N��4�w����M=]0�A��o@פ�X�b�ǭ��B��-� }�%H2d��ݴxdG(c"�8������r�R8^_�9 [I�@uIf��o�l^����\,�K����E���mq�KEK�g�����[*}.��$�xO�� ���3��v�������@�[	��Մ?�%�2���h�c�����H�'t�"��}�# J������5��e��0�R�-�l�0�������� ���-yJ8Q�&E�%S�ތ�]Pg֢Z���QIR��J��$'7x�S�=�u��P��>����~=t!6g�3�y/�*��c�mڰ��:z����oKW��ћ���~��m��&W���	��_���W�F�p�. ��L�j�^[*�IY��O!�F��K�F���/��a�=|�q�\�^6]�+�F+��b�F1�CW[0�����Fu󐧨��y~.a�5^������b
Q��s0�:Tw\w[�Ư�������ႇGۘ� ����G?,�W�(�ipºr7�#�ڨũ�G%�*��+�DO�AG��_�+g�B_ B�i���B��/��B��Okf�ٶ���٧��/?��'i�1���(4v�	��߯�: d��z�ٟm�=|EG��J}���-��? �]�M�����Wb�%�|���yQ�v=���R����)SqԊ4��Rd��9�r��Kc���7��Py+؅!O�6lm�>�0���ޜ�n|u�	ў�_��0�|��Q �;d��}&��6<�< ��{���K������є�}��^H����ɺ|[?��2'����t�u��.}�]^J[f���ϯ����F�i�LrȒ�W"D��R�Ӵ&�[�p�%���e�a��tʬ}V����|zf&��w��sY!����'�>�i�j�9À?���v!O�AD��+O�u�y��~�֛�0���D�"q�CrYl춱��9V8����^��܎d��Z��x����1���?i�3��T-��Y ;Hc�� }� �1��c�˃c���w��Zr�HP��Pj*4$�T�mnO��5�6�'�3��� 77��R�́NuO=�}���AB�N����l����6�x��z!��N�a(U�u����%��	M�&��y6��e�em��
�v��q�~w�!j.6���N����yh7����b��xH	L[nZ�4Z�0����J��QpZ�/l���#�eJw�J��~�x9�/��Dm������es�,9��qe�͒����/E�ݾ3h�ђ�v�e�M� G�X�����Kd4�Oײ�@��QN�j6�H:4O!"AYx��T�����m��4�d[ק6��������8�K2'�ýC�n��<z�SU�DǇ����z�~���f1��j'`<�>�g7h��lɏ�%��&L��|�٘��5�/M��_�y�z!$,���4����Ѿ/X���^��`i@:@��J9�B�D�=3Z���g��L�)x��:�Y���@�{�5��^]Q7m���]s����M���Z�k��Mt�DO�	�[�g��Ԍ&b_��V� ��ac�T�`T�H�O�n�$�$շ�Y���b2�QBf�9�7�e	������d�pX��(]��>/�7�4M����-��̞`B�����%�����)wȳK5�����Flc셧�g�zP��R��O���\s��0 ��.���͏�)w:*8Eu�#4�����Ec$�+Ʒuu�� s�+P���!���L�ꈎ���	Z�/F���\6�����AbjR��wcZ"���!$@������|yB��˫8�H���su{��눧��J��w�!q6���p�a�hEz��)���LlgYf&qvKr��{�ޢǾBI����m92�"�)%K	Y�&8+a�b�o�E�'�U4�rL[o[x�-�Z��"V1�B�@�Ds�i`�`΢�$eR� 	�B4�
�$0���/h�ӡ]{c%�V�V;6��̄�%B�\X�Ǿ`�U<�ޛ��.�Z.��N���:o�i7��v��ώ͘G��č0O��:�>�vӶa�Z�O���Ki���P�k
��~��E�r�hEn0!��Cd�X�Y��q̮F�fͬ��7���г��Ӻ�S<r�O'j�!�#W*��ș6$��m�=1ѿ��	�zD>G��W)�R^�=�sR��������5��v�~M.���+��:���~��������6���/�����.�>�Bu�ƾ�,{.cV��6�@WP���;}lɆK���/�=��������k�)�~a6]5�5*In�FrB��*���D��Ƙ^3���.�HJ��K��c�%�BL=�^��}uo�sC>���=Xixſbz�&�i�m$P�BE�{BB<�f�)�g8��"��m�����#��,xؒ����0D�!G �K���F����{��y=醆_�e�b��q�,��P�=��3�c�/��b+E&�`ɹ��0ecP�ą�~������)�'�����������W�l^9��Ĕ���j� ��NP�"�WS�/ch�9HGa,;��Gs��!�����
�v���g�����a5gU'?p~!y"3�����H�MDj�"z{��iN�<�x��SG�iF�4M�Ky�޽�:���g����o��-|�?KC��DGU���T�����
#��./�XA� ��h@�G\����i�8�,�H��P���#��
�
]M
-�d����d}C����A���68�KO�`U���8���S_S�(�C���^�Z�	RrH�ͮ/��h���>{��Ο��l 8I����5� (K`�`Λ��P��ᣝ$�d@5�%�u�����+��x�*]X�3h�$?�hR�OO&f�Tm�F���h���vO_�N�tT?G��W[�h`����|�b�J���$lXl�K��������U�-sz�»,�")�l(Oh;�kU�{p����`-��&{I]�<`��o'���|��yN�����>c�6�m�t�~�+t�Db�6Q3�
(�@��;}#����F>�p�ZZN[�3���d��(K�2v֔��E�'!�@)z<�\,���n��m2�$�xJ�N��uDG_Ub�uLU��M58�k�=����uw��5�, �F���!�O����|aF��@��}Z�4
=�u�R\��N:��RCM:0�X���9���bΗ�H܃��2})�уaӹ�����Ј_Jw�@�b9 s��w�����hs[��@.��ڂ$������������U�^D-��/�b�>}���
�1/���:�޲�䟺?r���d�O����;df�?A�:vl��h̜%+zH`�i�v�m����|o�R�W�h��n�gX�hj�� n����(W�,@�;��j��Y�t><�.
=m���?�V=sOS�P.���[�/��s`�Z����L�8�|�и�Ҏ���s=LވH��5���RLn&�r�Kmpq���x�A���^)Q6�(�'����sY��0�^=����%t����cG��Gd/(,�-����3/�=ؗ&s(p9��g����a���T�w��� ]��ڪ�Y=��5)�L<
��w��7�GCI��KqTf0O����,�3��n���Jea&t,KS�r����/X�}�=�9��cOF�0ti�	>����ݵE�e���i�{��[�����aC���;�JH�+�� r@N���n���Ro7�P��qz�Y���YN`���uq Y�(��ѿ�2��0Κ�9�lt��d_���΄����Ħz��V��!rߡ�V�D�h��x
8�3�V��oˤ�+��z`+���7��U@�����g�/(*�-x��ʤ�3BK���cg�w�saƽ��z��8D!mdQ�_./�x�k�G^o�e������y�ÿ��
�2�6�?Q�#GyX3v�Hm�.���f���ԍ��J��f6	�p��鑶SKUp�{��OT�/�3݁�6��8y&(R����Z��5�K� `Z���	|�b�t/l������E�Th#�e]s��P�Q�o��R���V�&t���������}���pp6ʹOZ��ʤ�������a�c������Mk4�D��/���%*C�`�_M���~ȥ.
� K��;D	H�� �������.B��n$_Oa')	ǹH*� <ϻ��Ft4�L�̊�������!��WI+LS��O����h?�Wݱҿ. U�����
�2M�{5�p�/b�?���ux��H���l?&�P�-��/m�r^M��~�F������QW6�Oꀮ*Z�{{�[�Mҝ�+L/��
�b�,�x�h�Vb�m�2�)X��B�R5�w\+�#�!�"���5p�*=���&<Wɏ��꥔���N8"8��������K��w8=�I�4�]�@M2��o��&byS���+4|ԧ���t�2$=2c<��!��2���$AI��Z�Q���� �ǰ��� +WyT^�z�C2[��x;3�1������ګPZw�	�wė��?Buu��e�J�p������"�Z:~�4��Ѩf�F����
�ͅ�[^�]'�����5��B$E��'Q&G����Rc9�3�L�O#�˖�'�%rp�ޢ�J%�N�E�O{������K�PA��M��щ|��<�S͚Ѐ�q��8��>ʺ��RL�=Վ���崘&��!�e�k>��6��ֽNB.&�y�F�3�ًi�������)�} Nj�������5�qƀ�Xj#(��ྡ��X6�pDX���G/p�b�<��T�m��[(��&Fw�9��h�14v3�^�;�&k|�G�0�8�hR`�!oT.��B�4Us���5��~jn+C�~����k+R�U|����ӦǤ��ŝ6'�_��a1p�7���s�|i��f؍b���<@�1��p�&^�%'�}�@^~ܷ`�!�ڲB&�����`�D���o��R�ʢ2��P��oc�Ҵ�>��42�
_�&��Ж�����֓#�Y�R���
�@|���v�Pb�(qy���oP\	!ۣGM��E�
P�X�j�1Y�i1���F$�a��U�U�%�{�h8P�eD�iX���%��'y<dl�Ќ��>u��0Gc�C.3�af��VA��F�fmO'u�-�g��]�Ӆ�i�f��	�d��T8/U����[E�g� ��a�Z1 d���˶�U���,��E5��!bC�-: �g��0�@x�@�y��W|f�����m�x9����+N�=nB��[� =A�J�r%0�ވ�~�v���#�~!��W�)ya���m�����č^�g�R��{��"�k��|c�z�Jp�f�~C�G�v@Aʞ	�C&4=/�t�8JE`���9�޴Q"��h�yCp����5��c����ػ�##���H�R�����.-��HV����7@~W�EO�e�ST�6��b���d�k�	���Na]Y����!S^A���lW�����{�!f��O�WљMg�,*D�{0Ak% ��Z��0v���'-��+�+�����UZ���i����Ac*�%J�z���]�2:��pҠq�.��̭- �=ڣ.v ,�.3G����J| ,(/�9��\�B�H��B_O[<;�Qp!k����1�:6����`�?��ZU��␚n���d%�9ƫgY�9�s�`BT��I�e,s��uXL|�Eb�1�I�v`��u̓	g���Y���Z�����5�]v�/�1�g�8 |��p��/e��G�-��V��}����	$�Ń;����ZЍ��M뻿4$ �lg���pڜ(�-:���&U�紹̫GEQ?�?����]�;l�)rp�W��Der)��m�ӌ�][�G�
)y��dKv�u���|m��
�����q1Zn8<���`C:W�I����K�0"<�)��cMjl,՜�~=���E�[��z/^l��/_O�)��h_�מ�^㹪�`i��I̼��D��z!��p؎w3�r�8T���>^�|#5J'd�O�����,&�edL��z)&sI�~�˙�D[U/��ЙZ8��G���?�i��l��N��i�NP�p��H�3�����q�B˸Q$j>U7^C���N�����9��Si(���f�G��(6��suɓ��қ�h�ѥ�b5����B�P&TO���
B��%��OUZ�<:;��3��K��߳��	~��:���1�*a �,E�4�3�����"�/-ub�C	*{iq��3 �YI�h��#<p2��.+�X��B�W=��g�I���Qˊʀp#̛�M���́��VR�$�a�[����Y�����H�ĮI^�ߋb�ktG�h�3q
7�d`k	u�5���\�r�D,���R��3i뗏�Y #e�3��me�1���E�~���U]L��1�-m�Bh��p����w�7�.c�â'ߺ��)�Gĭl-tp�1�6�Lx����S�{/�?������*l���R��^��^0F����\,)�G�7D&R>�C{e�a�g�����/H�8�%Ռd�����Al����C�r�Cn�{�r[��I�MH_).�2���@�!�0呉.i���>\v�To^�sW�dV6�W5�w3@�"n�Z�/ue��Q��i�v��N`7GE�ш<�PGo�T��v�^�p�W�۩����`�e����s�LL����� �bjn���vo���Tq�Kj����>,�'#��֊�0��A2ْh����)��f̑�|����s̆���H�C�>.��@5�֭��M侩�����C�z��4�4f郼�.��`�d�~��
Ǩ�d�I*�6�����#��Y�l�y�<M����^��V ��N3��)���Į<ȧ��4w62*����'#[��	�7�����z8J�<j��)����o�ϟd��KZ,g�UC�l
���T��/�Вg
�*�A��Ev���/Fm���>pOh3���VY�ǩM�J��Ja�g��*"�]�D����; 
�nX��r�~�֢�Hki��J�:�g�(�X^O<cD�H����B:�;�0t����b��o>��z!��I�ᛞ�w�Y<PE��\	&r��_IQk�=G���t�ı�{�0�,������B3�p�
��ġ�99讷9�hec����\
��
�wF���7�;�UV�'�Wb�җ�b���o�d���bFv�G�����)�t�`���&� Ԇ�3]>S���f�Y����	5Κ9j*�\�(:��C� �=����'���o��Ocn��4G�^#����4��c�FF*��}^
�j�
}�JԹZ�"�=����!	q,�p�x�ny�y�Z9��G.�.tޖg�E�d�8��N�{����I�,	�֋����L8��A�S�8�{Qڃ	��rl�"����1
F��9]�	:C��	�wF��h��р�H�o]�̃昭��L�p��+��jr�z�ڈ����a,0 P���9�-.l�ՖG�L�j�� 4�%���f	e��h�4�l���*�g�{��7��~A��<=����(��]Ҏ�rϋ�qaM<��0��T�����VǝTS���	���&��/8rt�Y���W"�4��� q��h��n�h[?�lf�ξQ����5�҆�<Z#E�B-�m�A[q��B��:]�A*+o�W�<$��W��G�v��:�I�	�E�p�*��Q���So������IbիʩhӢ���+�,%�����-��\R��-TW'��/:����9G^N<�k�m�=ҵN&d�#W�]�z�]�	�2�@r�|�q]i�� �4��q�U���0��mm�^.c�����|E<3''3�I�W�(鹪1ZTw��z�P݇�u���`���{��B}6�ɭ�Ҙa>lt�N��[�Qo��_�3������xp��:WT�����G���=�\�� �[���g��)���h��O��eŀ��6�~b�[q����a����d<����B��YP\���VT�>�ڹ�-u�E��[�8�6����O7�!�K��G���~���<���d�K�ú�O�
������	𹻧��$�q�DTY份�vӉ�%z���O�'cb��綀c����>���U����(�p�R3�u��k����� Q(�o����=�����Ƭ=N?�vt� ��_�K:��zr6����~���L����e /HyaE��2�l%�P�W�T?���FͪAN���Թ]%�����8��U8�o./��'1@9�~���f��.���A��:C�P������x����#��sSQc��	�)�KD��2I�	�p�T[�gJ�?�!�\�W����%S����%9��>���
�o��	+/��� ��7A�D��	$���#H�X'Q��[� Uѳ�?9�|F��t�#
����RR�1���0�T��Ǫj�,*�h�*F���ѭ�%S<��E�f�*T����͓�6z�!|���w�2���X���H�����a��ẇo��dP,����=�y�q� �<��I��P;�Q`o&1ޕr�u���.��j��S(9�����ݺ�)�R0�F�K��u�r���f<�{iM�[�"��qP6���3�8�W��X���Hkk7;_	��q��Ud��/�hB���.���1�@o]�ڿDc��XAJ��������4�j����]����ذ��2y��Ź�Ưq��m��?��P8B�����_�\w���� ��J&���1��Rǰ1[�b���W��J��86HeA��	���.P����j"�a��@鶾�����'�,I�
_���X��,�e��9g쌘?>�۫�����Љܲ��
��]�y!w '4;����̢�E]�:d/����	�,f1Wwm�Of��s`ˊ��u�5@�i���h8�?V�z�>�*KIp�����g�)��Q�:w�"{t�H�z'M!!�H��|�l��5�ɸ��>�W��me��u V���r0��6�i�	d�p��&�^[�6�>�.>wlѤ��}k������"�����Y�V�5����K��qpX~ T����R���F;�e7�ۈ�&�T?0Evt��A߸p3[b�tSF 2��Sp�~]��IB���7 ��i���͔��q�/���s��� w)�|&֤λg�]#c�N_\�D�}��.�Tr�2a�����?J�����Br�0��}N�a��ր26���ޑ�O���Ɂ,��j@�˂9E:u�tK<~ ����Յ�ĕ�O8�����4J��6'm��������ȋԖ,r?K�p�_H�Uy(s�p FQ,�d\�eṬC�ɰ%`��'6�E�	�:d���w��(�������?�wأ˄�3� 4�*��o����_��e$�gf�>��s�Jì��We�k7����dS�a(Xn��o�P����$�J�j��\�A��:��Yg ��&H��
�P5^� ��gX@��D��(�4�hG�|�i���A���I����>��??�`��^@���)��@:O�h�t�I[�sF(!�x�w���⦀Yc���d�;�m�,������0s'g'���O��A A�P(m}�����-���B��Ζm�Y9[ּǶ��ś#=�k��b��-��tǺ��C�����Un>E�DoQ��}:�ΫN�_Ć�`>�Ӱ\#��o�*���>~�t�C�! �"R�0���6�pYȻ.4�WI�Z\�[`UWr6�t2z��.�c�/ΑZU&�|K�
��񲻙GZ5�)�<�=��s �_���x�s�k ���׫P|m?A2�YA��ӕõ<Ȱ�tC���&���%�O}�9t;f.����m-mX�s��:a�	����A�z�S(ٓ�̞l�:񎺢ϺM⽟���;�Ј������$�+��Α��W�Ǖ���-]�"��N �Ζ[�w,�c��}�8��``�S��R�}����E��2�Ҟ�09jy
��~%��:��V�#(2_:9�/�������[��F}.��i�� v%���ӳ6��F�&��QȨb0D��H��Q�!������{�����>�Lb�b�0=����4m�j�����x���p|�������>$�$�[�5�G�<�R�O���c�v�j��[�R �O}'ś�����u����m~��T�N������\�Z����w��ֱE����3��K�^����.� �w?�
t�S ��yX��s�7ɿ)�x���=�\���R�I����-����e��R'L"
2�h�	�5���U�)M�[�-*��]���$��U�}�#�Kh69 $��{�_��vCV�g94n�6cT�N��j��G�.���&�x��7$�&��6���G�g�M�OeځVvf�~T������S������M�.�󾎅e3Gp�VT#��o	Ժ�R	�!}�I�_ˢ}qrL�%O8�L� 3(��4��%��;��w���a��& �=C�X�d�>����oo���Qh���%*�5?���w�{�@#ӎ���~T_#u�4��Lpc�Fcx:���U8�5vK0�g�v�p��U��Q$�%�,��8T>}+Gj�}�!sEB�6�&�0��#KU���h�U��Z�Lv���W�v5B�"�Ǐ֫Vۏ�&�����!�0 {�aI�,��)F�d"�����=� ��W�܁:6UpRc�#|�
f�V���g<Y�(�ow/[�U#���;�����2�#����c����s���KyT�!��'_��S6��N (����Sh��@�A��y�3�F�n�qP0I���@�İ�n�K*V��(/��ٱ�k�j5�(�u.5��H!�цG����^�g�%��lT�u��hI	���g��9�����%"*!4 ��O3��6v"�b�a�QUu
jF ��ְ��e�t�&��a����@|���9y��D��%�"��+P��uG<֟�~�VWC�Wy�