��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHnX�l�eT��(�*-j���Y��ϓ%�n0<W�*_o*���ſ��S��|S�u�r��7�r��<Q��������{|(����k��4x�[�?���a��6�v��w�ř)Cp.\
=��FE�p��I.�d����<���Xs`�&��	���D����B!�����^�Fb�d�ٻ�8�͞��&@ʹ����O���+f�Pa�芹B �_#��t�U `��h�g�?8x�x8	B���	#�-T)m���p�|��D��i���N���P���H����Rk\ɥ�L��\���R"5��BErZ/�q5x�'+�=+� �����˭�^p|�=*F�ε~�8��Z�ڊ�x���~��<��@�s�D�$�� �09C���v������P�K��2��3���W�˕]��ɡrC22�~��=�S�n�E<���)i����;^�TZ�~4�1 �*n�Z�\B��&8���O`2ŹS"z�!3,�(ך�6,<���e�Ư�2��2�䇜z�K
2Q���,�������aBH��Vl�@^��7�����Gj+W�V���,/���mɊ��}y��v�û5�!l�Q�yL��Z����>���IN�%�V&�z�[�����e0�W�]�IF+��r�B/�I+�컁��9��%%
f�r٪���,����=�����>��*�B��Y��-]�x����[Ĭw�t�u�����ÒD����w�ڱ�H�ٍ��9���fcp	����(w�N�ᑟQ��S��_�ύZ���;������ue�n�-N�.QH��'��y,�9�#�E��f:_�h&S���~s �<���qʆL�����a�)��U�GBZ�����5r�����f�g�m�ۏ�@��h;k ���3OJ���&z} ��2E�p�z �
�f�Į8��(S�P���f�ZVI�6:�7B!"T8!ϻ�t�K��3.�|_��	;�"}^���RsnG'�އ���::�u�3�I��w�ᴶ��ѽ��"y�D��Z�w��M-��`v!����������W��[���CFr$���.�q{�=���`�j��'5� G�{�������!e��#��'�őbR�O������ȷzz�Z�|&k�W�����k�#�SSUQzĥ}��@���"�(�1OuEX.�=�%kR�3��!'�N�$��#3F�}IWd��=kg�������Q�p�Gܞ�O5�\s|��͑���	~U'h��5/S�����,_��OT{�}*��0uh�:�U���M�R�c`�Gy��俾��)�@ *�����d�Gh��{�o H�DKwn� ��� 4f}�#\E�����}Q7;�p��Γ<�Ri��ꠡ�jS�+��#1���lVH߻i�R9)gA��y(���U�A@�3)ү�.FZ�w;�4A��~H��̏St�eU�
��Z1��4 � �U���ﰺ�ZjC�ѻ�w�����_o��:d��]���)J�0�^��iF�}\(����gƮ�׵��>�vG��U"�Q��_�5"������Q����
�jp&��B�F�AOt�����T�Q��I
��B4�TB���s�|d�Z5�+�g��{HO� �!�"f'��
(�s�y0/�(Z�E���Q��`�q���ܺ�9@M>�z`�����*����n��N�� ��]UƁ��k��ۼ��UoJʄ��A�~�q�=�C���O:y��f�� �du��	$��l�ݗ�����/�$��V~,�g!v���'������n�-�t3������4��W+}��7��5�{�;8X�X��N�l�A������d|��}�:��$:A�{̠��'�6�X�y�+�d��5�"��b�ZIz:��3�X-�Ԥ�
gg���,��}���c�ٜy>,:R�����}&�K�Ł}�ʠ8�{t
�w9��Xk�o�����I}D�� ����¾Pzz��|9�v�ipi:�8��A�>т������/S����=�%)�phTš�Ih�-�O��j��ɸQs�<8y{�x'�_D����F���x���֠�H�he�$��N�\{���b��`�}���\���c�����.s{�L^���)��	���Z�qBb�'T�~�� �sjV�f;%� 
ʡ��k?�a�����~�`R�ʅwvK@��L�!�bYp7�M+1���Y]{ߔ�T�$���s]��(?Йm_��9?̢{�稣3�+1sib1�OƊ���3�Q�-.��D�;�,(xI���o3��h�ŕ���㝕+ -�_������Kr9���鯚���cu#\��p,(&��-�72���t����P���$,8�G�O.��3���q`��P^M�����yц��n��^S1��t��Qd��#���jY���?З��`CJ�~�+��a�l�'i�l��dg���:�~#���i���~�`�J��	D��òF�)C�@[g�G����+�
8B��(Ҥ��Q4���.�� �ڎ23l���s�*��b�]��T�hk\�����`����b�ܝ�j� >��FcW�na!�����/k��Ь��?����*Ul��$1�'��(�E鑯�w�a�����~�H���Q���m[�00o>/�mFU��q�n��O����YDj?y5�ސ�G�p�+���6��%�Q(	��_�	R���)�PC	�^�v�0��C?���x���6}�K:��7����u7\�Q�2�}n�"u��B�)2�ŅB�Y�|��Y�EÑ��\��h���4��6�u���n��ʨ\h��!Vkۡ�;�%����%�����3*��Z��t��:�	!|z����$`���u���1�<:2�b���YY����{�+v�z<,�d���W\�����8�W�����t��BQ{jA
o��H>�m��e�C��::BjϹ��B��������$x4�6O�QHL����(3��fӃ�3���󧳂.L�b�2qC�\8