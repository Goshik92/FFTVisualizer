��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܫk�۸�m�i(b[�{�㇌�]�i�5'�`;Etg
<������H�W޵α��wԊ�6�a�3� G��λ�:~7 !�v sh��~��P�'|#��x�C�[�~���{-چ��!�:���)�#aE�C�;� ���&�'��c�w|�:�)��$��Sއ�Y�K��N�4uFLN��6n���)G�Kh\��V��V��ie�� �$���68D�"����܀��ds�ʄ��]�,�',��2�\�m���
��q�w�<����;�jCZ��7p� ��}.fV����|)]"��A������QX�C�s�n��ܓj�R+TlM!��2-�Z`���f&��1v�$ːI�:��`����a�c�_�8�up�{�{�3���b��ӆBˡ���%� ���P�r������goAMp�B�zO�RV�rʪb'�2\�Ok�:�L۳0
m˱�ߠ�4Y*�6f�;9���~��, �7]7w8��ē)�;����g�&Y�mϝ���E�u��T��{��7��m�R�ڮi�8&������Ժ�)�:.�|�q��y:�r�?H/iO`���A����4k|'#Xe�+�3Q�b�����yW m)�����v}( ۼogȡ�C�B �h��C��or�_�ˤ<�����>�?�o;?t�'	���`\��l���7�w���Z6���bKe�'{�֊����Pi<%���C?p�,Op^K�������vrK�����uנ��Zl�$��uV_��iz7#�	��`�`���>����^r��K�ö�5�.D&Jx:P ������5$A���2bp�%��E�A�wBװC��{�Mfsf���/�uݦ��~EH�o�Ҟ�Dբ��L!����%)�]*R����7�cػ��=sp���"���oѡ!׳�Re�[���{�r���"D��8?�շ��L���ϛJ� Ѣ�-1������92�o�u{�<=l���} �H�]H��khu >�_�s_�Fq��1����Xf�9'����-	 꾇k��)�Ϫ��K5�]���Bq)P�)_2!�Z���1��,���f�
���(�#qs��L�	�:k؟�%�9\�Ҁ���E�:w�� �0�����H'oK7����=�;�,aַ��`�Ơ�͹3��OK� ç�_�~����9-ew�94tE|P��7$�8ˠM�y�}Yg ђ>�~��#:g�˝0j0��`ƬC��{�#�Ge��]�^Nd�����(����	�D$#�����~��W��� �BM얓�`ӣok��Ax�E��,�E=Z\)��ΠEpI�l
�?���`�:|!8���-O��Ou�|j�6xe��Td�	h>��?a�ד���@���L����`ZA���q[�`C#��*7>�Fr�s���`��� �_ST��T�vɆ���_.f�6��ZmR���*0�܋���"��h�c�
&j#�ğ��6�u���6�E�Ԋ�l�xQ��)���絶�?h}8��R��K.��R�w�f��U�
&�GǍ�Y� �׫�RgE�_�tz��.R���T%��u�M�.������:��UN[%�:8�^���LH�Sb��F�ݐ��,��&������x��'�$�,��L�殇E�c�Z��لR�k]2��N���]��R9_;/��!N�=��OM~9Ú|�efV�����e[胎�ا��-���i��T�pR���E�*ܾ���S���晋���2>�E;�:h��#M�:)�XY��k�1��BN Y�{[�t8��+A�g��:8R�MЀL7�LrS:���jh��~b��e��k�	up{̶#R ���B��y�4�|kw� ��T��%I�8)-���q_�(�aJ�`�I�2����Z�
L8=�U����H��F��,��o`	���"�L��#����}-�Y�NyT�bb�"Z18�1��t��/'>�N��ҹE�1!�I)�[����'�(?���ꖟeNzCE�s�@�EX~����n5x�� }�q��@�us�n7c�wD|��p�i���MU��KmxAԠq����	�r8�����z�������ԑ$��$Wg�
E�Y?=�?߇�JE�MvZ	���{*�r��M����,bZ��;_5a
����FҤ&�#+�>�_@�iur�oq3��+M���R�B��
�)a��+���@���	h21�͎�?'9��&S~eY>�͇E��a'/;e�mj�I����m�$4����I�WePA8�� ��ي�*}���'k��DC�)��r�����T%j�����������ygeZ�z��2��ڏ�9�@Zl_�c�� �l�s���<<cH)~�,D��p�)��Y���_�`��en�s�p ��I��B�cQK��ԔН{��ǋ�iNF~np�nE/ KOF�K&3L�*�}�q��PP�	��:4�h���ff���܉��^�28`t��'w�v	]�7�̍id>��	Fk��p�;k\�����f5�\�a��Sr=��.�il��q�KnHB�f����<^��D���J��\�/��c�L��"d?��\=7	�&8�Y!��+I�ʋ6��.a�.�.�d#(��F�� ��.\"-���;Ht�D�����`�@��\�wTh�:�{�l>:�7�fV�����8p��v㟔-��P���I,
�%��iF�s&�W�rйOGjp\�`:��ܖ��fך��c��2L��}A6[Ru��΁�^��YJ&1m@@�;+
ǻ�s)9���By���?���A����״�W8��0���NG,<��m$a��}�&�X /��~���3��u�rm/��w�ߎz �~n��7x��6���Wg� _8Z��D��d7����@�VMk��!R	��cr˗ghH�ɣ�Ŕm���,�/��L[�����X���Ñ�{�	%��Ib淍�La�)�,�l[�VP����Ű�v�Ȍ#b�Pg4N���u��pơʬo�B� eD�I�v3v���O�;�-!�M��)*1�z!4� �Y2F��_bLoB�>g����ho�w���t�X���3�޶��J�jnZ�Yp$O/�ϯIp�#J��oη¼ݩ��]�U�Ȅ~̵w�������