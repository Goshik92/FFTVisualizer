��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ��p�oȡ�;u0ީ�^�)�>vys���2{�L�~|c_Iy�K����-��9!��\�Bi�D��{�Ԣ��r'T��NjH��ဣ]��9��|p���4d��oc���_LG����*k����۾�T>x�/>:��e�=�C5!)f���86�$����ԤE���oZ�&�x���� ]1����V'���Hci������I���-�;����{�gr�HR�l�q����~�n�2�����̴S�c�6�'o����f�?L�2���r�����uq/�Z��a['R�)9"+",��:�l/
����#���U\3�$π��`3��J�,�;K��=.�ʄ1���c��ą�&Y+[&��z{��/j��?|��~:�%��?�!M1�3?ߤ�	d���j"VlVg8��j&84)�|K�\�Y��m���TU-�^V <h�Τ�4XU�/6�����X�_A����W!��i��o��>��B��.��9C��iżׇ�2�%>+o��q�(t�
�%�\����·�*,U��y�oxmX S�`���;�F�S7�
�(���!�e�5�I��Ey·���e�`
&NTv��n�������Րae�m�d�9�<]����kw/��׼3`����ǧ=��ό����d%;�4�����"?E����R�m%���<�:F�Z�䕼jp�j7���P�U����AX�����:;��}1I>�[Z�洽��J�(T��(A���ik�sO����al�	�y�7�Ady�3� Ck�ѐ�9���#O�XM��@ŏ��X@���6�-i�� �*D�ӆZ-sa)K�7�
�3�`8�"\��u������Axw|*�>�y�Z��eDJ��rs�?���P�ι��Q \�f�Q)hQ�&��c�'��n.l�.'I�X	�D)!���s_��@U[%�Q�A���"��L��֢��۾����KJϽ�U ��T�/�f�MYA�����������=��D����e��|E��T��_%�����̸;�[�T�J������i���~��9׾$T�r�j?źR�o��*��C.�������uׇ<V�6�ĳ��Č�z<\�^?�����h�%X7�mp�Y^}Oa�V���_�L��������|fMX���M�T�B>�W�~l2��pVS{N֟�c�l`j��p=����:�(��e/"ժ�8�nƓ�#.�6a��~N*4�e;��˖��b�3�K�l�LP�X�7*�H���س��������u��t)��^H{
^V7��b�6%t�"���9��mG�hDc����%�@XȪe*��������}"���[�U������<VX�<�ˆ��uY5FS(~.hnsXPGw�8�����8����ћB�R(F���4Cu��wU
�L�Oț��}T���+֘e��G���
��Sl=C
`�<�u� �*v�xeҍ�ʫĩ���z����V�ޢj�M�#��u�-�M��7�x���ȦO�� ��u�v'6!�dC�@���(o�P#�-��v�/5��L)��Ww'%�l���#�A��0�~yΡ���M:���:a�<�z(�t�z�}��DG�q$$��n<p!�켒��_$|:����$��[r9�
ĭ��F�G�O	woz���UH{��$r|gN
:���	ߤ����v�X��m-F��`e��^-����`7�gI��-z܇F�u�tV%>���OKV��l���^�=r��v���ŗ����<{`���_�)u�g�Q��F)�ԥoT-�4��m�mqH5�@�AHğ��%�@�q��7+v-�"�f�ϐykPŮ!��p�dXA�5���5��q�}�pi����U��Aj,nv�R��	���6�i�N�.�Tگ6�v'Q��چd��M�Y��4
`�󒰇�m���c���ޟ_F�����p,6��*Jf44O� ��h�Yx� $4�u6.����}��\�^|� ��гgt�wd*���w\i�7U4�f:��,�6�:�XY>�ï'������L?p|�{��8�E����`4�����˒<Ȁ�nC��!�3��[x��e�8�5�AO`.B^�'�b�e�zI���ʁ�qF�7?K����Zh*>:@�����sPC��}�.�M�b��� �yy��q.Kd!#|��z�_����i�Q�Ӡ���R�Sܔ�r^!p@�����ɘ�<�`Y���E�u���M���˶���d��m�FpA��J@@_LJ$���6;w)��=wgU|#.
�_ߣ�ْ���f���s�l�)�~I�>�*S��,`���;*��S� CQ�hnZ�.H��snb��i�I^$K�*�;l�� ,&"Gl����BT�����0����5-qD\F���4]�WD�U�u��iE�9M�l���[!(Y|gE���6�B��g�ň���������"9 c��Ռ���6^P/��g"���:s�x~��ʺ�?$h���Z��^�$=�B�U��x�#%�z:棥�VZ�YN�M��f�(��7.����)V�Lfs���eB��m7��籽�M�#L=C�]% OR
��M�x-mX�u�0���ʻ.,' �b�"D����'��E��|ni��OA*:i\�ԙ�&��4���e��<�� 	���Z��,WA	Gc�yS��V��b�t���f�q��!��0�g8�o �&DN�������R�pg^�G@cj�JO�(c����H�8���s�g�.��6~����S�Ō���C�1X�9lQJ��0�!��N�v��G8�A�[xzVru�b����!�*�x�Cj2x�c0q�+
���c���z+��A��4�6��uC�c����=�rt��*����(�y����m���X[�Ew?1�t� ��,��[�%��]��;�8�^�'�N[ᢟ���E�7��ߟ{�L3�?(�G�ʭ��[U[4��)l�R`��[G�è��4���f:�sUR�J����I=�)K�XA�ܸw�ߟ�
iA��#�[���`;ݰ�²����
Kœ��#_�2�GK7%��t��ή���c��k���z3�(qE����y��s�_�O��_�7��ژ̉Kb9UYfm�9.t�a�� ׾~\���9��gVh
8�1=	��k��n��"�S[�9V�Sd�������ɖ��]�^,��>hB�z�PKp�8�,�W%6�
�Ƹ�e4v'uG�-̅�xD�Q7�L1r�mt��y�*�Џ�Ǉ�5^�&s��8}i��:��	)��:<.d7��!o}`�K�H@t��ot7ԟ;-Y�ʏk��-vA��c�1�e��:��ޝ������bi�=�f:�o��(y_�ӡ���#����K� [�����P��*��(��<@.g�R�{�6��'9)ii{�n��t�Ľs@�p��c�@�����TyU�Ҝ�h{k�n��o���]�Z�.A/WՌ����a��<���`s�y�yR��Z�p �2�Q�@�.���� ��΁���\�KѾ�4�y���������W��;�e��؜��T��~Ja3��auBizS��^-�t���.�\]j	FB@�����We�['��߈��U��_����ˀW�p*��\��i����*tst���\�R�RbB�)3�<`_RlG��gׯf=^ _��)���D���iD���V
��M�]���.����MW�G�i�KS�u�O��$�}�u�"}�$�jo����������V����l�j��s(̍�w�6�-�f��P�ŤL�=���<{~W�W@�L���n=�iU۳�.9o�#��w�X{n��$�F"j�������O~#�g>���LT%�RUV�Tx���iizhLTwj���Pȓ$���xjWI߶��H�>Uz��o�y�ngd��.ȩ7��8�F��C���Q/�����Hfu�"c{�	��p�i9>���yn��g��Y i%�ܜ�c�~|���．T��r.K�¿g����ؠ޴$6�h2�\�vH����8i��+�"�vI1���1���b�7ͿS��}�bF��D��(	&���'إ"� Y0MжW˃�o����ϕ���8�R��׋�B�害�����S�ၗ�uC]<�KRXdͱ�G�qŨ�zp9�-��94J�9ĩ�h��LT� ������Q4I"���a�W$���$��0є*�E�m()����+���y؝�g�V�����L��~bV�TCx�% x��y�6!�(5�7�P�?]vܷ��r,��g� ��-���Ֆk�@:���k��� 6�P�/��Xt>I����A2i�`)q'�k���$���9�˿Ό16&И��t.�E��a�Fʇ��E'�Y�^6*y�/��J�P��������E���7a��.7�B�7�|�s`�7,��x�Ky��t�"�ahger�C5��n�$�?ԯ_��~W�'�S"������L��ǐ�������,��L����f�F�6��j�q�^,�Xe~M�	c�O�&��;[������ʗ=��Ur\�7:��:�m0�޷$ty�T�J���Na�*�u���������4�}����A�l��(:ON_�3o����'{l���#=k4鶦�#B��GSZ7z  �b�$�3<X��h8�պi��=�;�b-2����ɍ�x�2��n��#.G�ܘ{���ƈ�ż� Z!�ڣ��������j-Z\<��|���x:��o7�g��e����:�����7uEc�&i�NJFi�_+wOcY��d�%�{1+��:)����::�tRX���"�x�ט����Rkآ�0��^mx^��U�?�C�"௧�Vb1�2$�+ʨ��r�ƺ�󮓎�(.P��ʵ%���3\À�h�DB�K@�L��/3A���?&���5ɰYfR���/����G���JM0��:ө���$�3�kX �Hވ��je���3�¡��%�h���L+8b�	�=�N�of'�N���3�ὰ��p)���#���������j/�c7�
����������"�Dۻ#u Y�,�Cl_B8�N����42��4#��j%��/���@�넖�5���|b4!u�m��
i�LL�C�S3������}�<�Μ�T�'���u0�|C�mw;����/�p	wl�|P�^��Jπ`�J�bh.��|Tp@�>]�Z�z�+<# o/��\��RȗNr��}D9-����z����8&��#���+�.�^5F��k���*�LV�S9͕�pŸd�c�H�=���w@z3�(Y���OWs�&`ufzb�zd�W�$̌������'� ]N#�N%��'|Z]Naՙ��M� �������˕ ��P��)g8]Ж<Fe;�`n�;���j�����z���Z�JPD���N�kw��)}�5�=�سxpT�����6߆3<`:cȒ�}.�:�|���=�) H����A
�moC����7Ý����<۴8ʬ?'X~�LΪ��R�S��jv�S�$m��Z��"�dW��a	��G�鱓��d��{W|�Y/N��������㊿#���	R�-�8ăA�f4ބ� �ihy^=�L���������A�M��ǐ��k��0HҟtF r-���7� b�?�5� b�Nv��$&q��A:�"��!\P�^��z�(J@���K���J���֌�6��d��l�����Z�b�y�j�aA,�t��V��o����!;C�#?�_<�[����s��|QV��o�DQ�D���B���E��(ei��_ �eVC^������bC���h�.��iѲ*p`��l���bE���郕*Q����c���b���o�=�Ҵ "���z!���?j���(�J�5�2��%�UNV�V]8�Ba�f�j7>���	���'K�s8|�Yg^Ph�q�f�UzQ�~�%��