��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn?�v,�.f@�H�z�d������fM�XV#O&.�~�=�����A Y�<�D)��Ϣ)>�Nƕ&���������tFK��)�{i�8����,�M�+����pW_�F\��2љ0�����c���1=�X�����%�&~�5&�aL��C�%�B�ˑ} ��vP��Q�V�A8��O��#$�o��vo!m��P��F���eP�(t���5��A�.���d4���%��\�	G���tj)U7'R�w�A%���Y�<�6�U|;Mt�=Am�l֭?�����V�G�c�7�c��ɗ�nT��b�u���8+a�r�<�v6{l[0El5-�/|�h�E��p�\/^��"XUl�bup��;ic]|b����<�T ���W��
���^}�#SI��G*��8���S�˛ ��W��50ڈgꇗ��1��J�͇}"Um�}��G[�2�Pǚ�E�C���� (���
�a�n�+�T�dd	��c�.rӀ�	����\�{�{�_����M��P���QQӢ��g��,=��@�R�lh>u�[�ϯu��%�@��8��1'�*{��h��rx�x�3n��J�̏�z1;Y4Vp�)7�W�-�!�r��5������)9l`�<�6M};�!�
�ShՉw�^7����u�����uSא���y<�#blk�x�2��]\��\:�R)���䴃��!�@p��b�;�H���Y�z��rR�;;�zb��	�*��'�F%�T�����d:���s0�9Dh]��adh��8�z�dq�0QAJ�$k����2����C��L���Úx@$���!b�����^��͎�^J�ر��!U2�_�Kx��"eݣ��p/�J�rL��u$�lj��^�E4�����U\Qt�	|�awE�/N�@TE��Z��P޴I�{����t��kM�кL�n���A�wP@�;�P�;l�Ʒ3�3K%�՝R5��䚜���k�]'����ǟ�U�{�w�x���8X� G����	�5^g���6�N/R/��
Y�9�]����"��IbZR���j��F"���X�xZǆ^B�Jp��*A�zl����"Jw?�A^��lut�A�����m�>��O�0��f�+���N����4=ʒԝ��sh� KV��<UN롶n��؋*y��d0Č�BS���|s��2K�� �-1YzW�{�oiBmV����"��pe��䩀3
i���՜���p�ׂ>���LԵfi��8�c `^��wZ��V����M�"��)�������Y>/�,�<u�&�Ra���W�j�S�7X��H��¨�1�!�Q5}S�.X-�_`�LԲ����^+Hd�{�TQ�Ɵ��c��R�!��2�!� E�\xB']�ACi�IA_��B����a<JJ͕z��X��]�v��#�U"�W��P`�d.V'����cE��c�tȅcږ��5���L�h'�Q�l�^�u;F��@ut�{�8>������?�a�(@rV���\��R�JC2�|��u���9K��\� ������;bZ��a� w��U2C��@gg���I7ݍ0T5�ӥ�29�0	�� �������{�s�����Bʄ[�7?����4��I��,s���_�Z�0	����]�XD��l�N��?r�y�cI^b\�PN�n�5Uϼ���a��}?ekÃ��*k�\��=�	��J#����}��X��֗�l��ڭz. @��}�k�2�i���������YJ��>�x��3��h�Z`�j�`~��K��S�O;X'�z��'3����XDY�Լ�)u�H�>v��XD�\��M�⬚R�E���6��Ea@W&���+�ۃQ���4��_��*;���A�7Tu�lEg����W3=���Vz�4��WI&Z�o��=��׽=�Lf8a3��G�|Ζ�uYm-A���.��v3?l�=��gn����@���(|���T��ʿ�5TCJ1c��Y��~���3g� �l���2��[�v:������L�E���-f0�oѓ���GI�y��:5N�^%�텤gt�1��y�kEY��z6�Hܖ���2Ԅ�E����2�_V�0�bĹ̕?���w2	N�GՁ���aD/�W�r\�?���ɭ���h�aV�5)�?���5��5�e�"�֐�YZ��w�{��Z����ĕ�nT�%��"���$F1_}��J��O �¸��~�`�� ߓ��P�ʈ�\v�����,?�L-��B#�X.�J����m;�t�R�/m�uZΎk����8��"�w7B����Ǭ�m����������_ɔ�P���
�0�.8wT�T�auE"��%�h0�YK��e0��TkO���Þ�*�
B���`D�(H����f��޲z�<�� *K�G���(�8�sL0~9��v31<��-Y�պ͌�q>V�J.��&�����s��/���S�����]��S� `��l7'�ȝJJ�9j��x��sh��4���������0�l�/�Z2�cYiY�E(�h�kr#�M��Ҳ�	�y�M��n,����A����2R�`�#�Yw���*Y���}y�4k���;y�շ���=�MU�/AR��Go�����_�ةsN�?{ky��(��7z�~��㵺s9H��+�,��gK��n����[MO����p��8��0Ln41�����|� �d�9���*�t���d�#~Rx��
���U&V��-ܩ��:�G��
��a��F�Z�o��[�=T�P+�%x�ew��v.]5��Jt����&��H}: qr��i�7^�L2���C�ySh�wo>����2/���h�#���x#	t�m��\f��%k{N�"+@�o�O�;�{�5<��Y5�\��GKL)uXT�����R�Y��ƣ��o�Wf�BQ(��٭N�ڤ}��&Y�O���8v�
�\c4�KQ{���q!�P�U�ޅ2\(���u�g2>���XZ%=r!�ZBם^6N�Q@�]����(C��{(�B� ���s{ռNQ6�#�\���p�X��;T�8�F� �/��~��"�@�\(`�p��頵�,�ʄ	�XQxjߎ������jr�, h��z�:F�17t0B�_Y��W�	?+���ٙ��Z�,�il�n�I�n}��.��,�[KA�G�T���X���'��d��>����I�ܜ�b�ʟ�,�ʱ�rv��A�쁄X̱c擎��1��5�8@s�����n�;���g,ߓ��5������ �]-��������4�U'�{��)x��1`:37?���c���A���8�E�B9Ձ�Ss�>���LAIa`�ET�gv_檭�	��>f��u���ҁ�G�4�V{�+v%�);�6���"���G*M�b �Ȗ��0�rޟMa΍����WF�+����9�Hxg���F��5��%�ӽk������HX2�K]˟��	�Ǫ�C��^B+"x���
�\&�z��
}w	��z��Y/)4��)R�$��[��c��Mw��UY�O���n��5�������qX~��c�-�xv�>��>�w�-H���;���Ǔ<�ʠ��c�)�ȴd�<����5�1P��/�D�e�����ͪ�����6 ��-��0�!
N�ڈ� �j,v�O�'Y����^����T�i��W�K����݈�EQ�)ym��X1�7oP�!};�7��pzD�;Q���ƙ��?���P%�.�O#oٔ*�R<=-����Ж"(	۸�Z�¨�%	b�j:K�EѢ�Ne�� �E	m�1t���k{|�ӄ��q2���9#Q(���0��]�5ޑ��6�� u�Nġ(��=_�~[��I4�KU���Gt�~ԓ�x��	D�,��ryATk�ڤ�%���w��@G�@~զ��ys�/��4��9�����2K�L���l�.H��$۸��<�8�&<�!h�h,���{I<��X�Bъ�p.�G�cZ��wi���������-J ���Z� A61r���?�X*K~~p���F*�M����c�
k������؍�EGr�MT���P�C2��>f{���Ww��^����4� n�_�3cq���6�)��VҊ=�����S�^�c\�U��p��~�� �U$��k���huH��nNI�KI�;�@�_�]�3'��ڣ{๋��]�bp�G�\�vR-}�� 2�!��( <���������\�V�__3Wq7E�9���#�֗ɞ��F֣K;l���TJ����A�c�6�:���E
|��9Z���<�i1Œ鹘H��*	AD�T��^w����)����G��(�����؏�!�ͷY	�9���.�0R��Ur>7p���| ^9�ԡq9?���҉����h�%3Юu
?����/G,�^k�L|�ԯS���"Mi�v�J��r��&a��3{F������`����B��,�c�y������f�ք_Ye�5�jz���]���y���V���Z��G57���<�l�;�Wa�&M�NA��=[�*e5pjX�ţ�Ɍ�����<'�i��7�b:��J�J
�(a&��_,w1oҲ),��
̻�E),
k������m�`�0(�[�%�\)wY@�^H��brI)�`a��jځb��/§9��u���ʛs}�F<SW�s���9Yk�(f�Q/�\*-S7E�D��g%�b�W;e�����)D�/��(�8��˭�ܳ��}7T��!T$���WK2��_.����������m�Q��fL�GL�J�]	't���7FV�2���p\؎��
�΋��D�����.������ZH��F"���0�|�c-�&�lH��W�*���ĉ��z�|������7,|�8 f�k͍�F��Eoru��d�oˢ���I������
���Z��҄E�Aw�r ēW!��%j��T�_�<fƍSQ�����,����+�/��prQWo�|�1g�?2-�ӭ�,	�r�A'=����x�T���q?6� �����#�;vޱ�ʱZ�(Z�E@���䝧t;��H`'��R3יX�Ǧ�j�E �;f�{4KW�[�����3௼,�㑑8~�� k� T�xѧ���br=t;�E�>�t���$$Ⱦ䫝����X�����Z��^+Y�k���瑍z
}�J'�,)��k}�=�iؓu�I>��翖�f����-U�0Lڻ -�6�Z���Q(r��=V�Jm]���k@< �w]�}��R��d����o�$�+�����s.y*J�v&`m����� ��y�O����*��;�9�eqX�cl�]�r�%��2��7h�/�{P�o����6�vc�-���h��ѷ������[ީi��H�����v���@����Eu$T���f;�oW���?�-���y�LS	��b��8����Uu��֛�]��
�J78�=A�$�f���b��bR��U1�|e[D�d���5ɬ^�����h���ӌm������SAaT���I3Fc0G�\���Y���薧��)����7���ӽH=�G���N���4$7P�>��&�����Kn�j I����~!|d�Y�_|��(�k_ݙ`�f���|~��lq����f�L�Ϭ�|�b�%Yߴ���1jX�&����.Sǀ�_%���"�+U�J�T}	��5��
9j���Ѵ=��n��O�x����w�H�3?��1U�s:CX��.wc�Z�Ŗ��DC˷b��#D�-f�/������^��*|��t� 9 ʷ63�'�V���=N�S>���U@�j-�3y>�fz�Ӄ�{�=^I?�����};f��1��[�-k��8$�&25˔����?�|ZיL�H%��˔T������7,O<�!$@��7=M�
�w������(�ZɗH "G���N�!�/��Wij��ۿ!�M��si
���J�<��K檃&C�un��Q_�"ź�c��F�	E�:J����d!�%���!�b�V	ʸ��$�¤�E�:`��n��0DŇW����|�e�����5�T�<V���zݰ�82���p#�vh|�9.yuО��R��?��%����̵�@'�ًN� ����V�7� z5�.<���6�f�NU,p�ߗ0�T�"�ZTE��A�d˼VA�I!�FLm7�zd�&ϴ>�y7�U��BKC���F�x?���[�&��1݁��Z�i�t�Ё�p�������u^&���:��L��ͩ�]��i������=�M��<�ϗnP�����B��'-ֺ�ڷ��P8k��r��U=��6C#��Q2�������`X�p%�s�/]��	sD{")�p�s�m��h�����_t��Je?�*F3|��^�L��](R��;muyvנ���Qܒ��~�-1���H����M���ON���$-h�I�DWP����B(0`��S�ԐW���&�	K���E��H4,���`f�c=�ԯ���m|$Tg�$�U���/-I�*S'2�7{X�����:�_j�O.��[�ړGwc�g�-�j�j�ĻwL���歠f�Y&D>`�:M��d���r&��f��ϕ����mQ3B?�kzb��Yd<`�"o�s$x+^E fpU~d]��6_9�feY[zÙ�Ty�^��j�.��5���*^�@5�#�,ЈI@�F�Wzl)6Ms�WE�1���bf��I����%��	�xuA2�O�t^����ĕ?�&yEHX���':[�<��љ+���r=7|��&�E(\�<֑%�P}�G���m��$�4�.c�m�:��{WSdp?ƵT�"3!9����~SMg�JA�xR��y �~.�H@@G튦T�w�M[��SK�9�F��:G�����Ov��[}����� �&NtϞޗ�jH��o� 
+`����};�y�jИ���w�k�\�� �{���`6�Z$�IJ��Vs��|ۜ��M�aDMy���@Bͮv���H�W|>E��#&w�B��Ie�H���ӛh Z��۞��� (�M���xoD}�[����仿IM�"�+���x~am�H�8��h9l�i�z�a��Qz�/dk �4Pw/&fOd�!~Z�YeB>LǻO.N}��s�_�o��K���^;{���JF�[����<D���8� ?�}҄�B�n�<]�,`m
i�U�+�Qo� �pd��Tx��qZQ�=�+�lK���\o�q+�u<H�6_m�.�=�aG.eիĶ��m�c��>:4	���f�\B>�`H)�ʰr���CI�L8贿�Մ�ҭ�l�
���q�"���y�n=&�X�aj3c@��0wR�rփ$�����K!�	@���/
�o�ӹ�^�G�	Jx1��e#��m�0��̋����2�}��I�i�9����s�,S�v�W��vH-IK��V�&�^�;�t(jyPƝQ}COF��ί,/P�w���������nk��U�ѮZ/�V�hMw����)�y@��Ŭ���ߢ�����{ˋ�V-#�͛�U��5�ݤ4��^K�1*Z���$wQ2
"�k
�WN����	i��+�1���m<u������bJ����{�k5�f\-�6M���׏	�|S���F�gw�%!��$�h�"C���^�m@ړ*� SĕX��ӓ�_�h3��s���� �����i���S�X�޿��an6����~�Z�2cp�BH�)�G &m���I�\y�(?a��/,�d�����qx��ᵍ̶�sFW  ��|�@�`�!:�q0��[�)��),���c����#t9.����?s�R�)ǁ$��)��-�\��f�ʼ��[����&�d���Z��[�z�oK�%4Emt4_5�R�^nzw�z(>�g��_D��6���?ٛ�W���s�E;��QG�)v��jy��f�dd�ެ��1R~������%�")6֫'q��\/^���6L.�A�0�5�v�J'�4�Q���R������f��s=8�݌E�ۓ�K;�B����cU��;�yu?��Uf@�%y��u�'���JM�j5 ���ۇbl�<�"�Y�^C���wd��Di�K��5uѢ~�#��x���F$#BH��~��1Fo$�_���]�l��m���r10��<&�2����q,�����I��w~N@iD��ỉ�~�S�4�0�� ���F�u�y�Ab�ji2���5��Q�j�#]i,Q9�y)��j4�^���x6G5T��4��7AԼ@����,�u訂��H��	�`Gex4n�K����7?�w*�;Ǘ��$��)�Z�;Çz8h����5c.�P��.$�Qw����w�c��sczh��j��� I
D���(u�������,�"�zE"h��P�H��R�Em�'"���8y�bcW��tu���/5�$uј��|�3UEx�0TqȱrxN(�t�
�YELy-�Qn�V�� r*v��~3�_���-N�]���1�-9��Q|��L��:�ՊI���B�O[��KU���֋��'ٖ�2�ODY�z�����\�����6//Ze��y�ZoS��V_������ �D�*4~��L�G7�j��s��؅:[2�8u{-�&_=�M%]���O<����������su�K�6��~!=ԍ����\��vb��v�����H�#�AC�I������ߴ�^�K��cM�u�	�4X���	:C�v�4�n?����@���L���^���OYA��k�;.���M��6����9\��'>�h��N��/��_LuxN?�H�z� ��K� ג�E9֖�	���榽 ��zY�������;���
���l��@���ź�'lՒ�>u����ǽ�A�d���U�����ӗ�O�eF�_�� 3��Oo�Yf,�h����R���g%T�1m(�2�7�g�
i]����Ic��f��U��tf��L�T��c��/)%�9�9-p����FcA��~�~��ݐ�h�n�^�a���a�Z5TLp��T��ҷl�\Y�@��o��vXt䭝&Z+��>�t$��+j����J벳��`��:`��������U�ҩaO�7_#k�6w>"I(-{k�SOul@�#L��K%!]�y��;?�~�FЬW��ȮHf�'$���으456b�t��g�m6�e�P=N�S��T �3yI����j��F1w�d���Ƞ�8�w�����U؆�nاrt��0�L���y��׿[sOTI�bDӵ��:�rD����OO�:���G�+�<p������
��4q�{����܈�e
�^�+s��W{Y?��])�v�f���&e޲�u���	 fX����Z�������}��p��������Ld�~�3&ѕ���%��8��ƣa
����b�b�o�+˭�ya��M�D���N�}!�hhb�&�]�3 pw=�f��[�y�d�K�ܓ�@�f���O�
o2�� b1Qk���?�e[��'!=�����ڔ|gNX�Kwc�4�y�3�tB*-�H�t_)�`�	(0^:|��a"��e�4TE��"i <H����t�=i#+_[�;%����Fl-��r��'�Ո���]wɝ�.���]��&p4������	��w��ȭe[��_;��8���Å�w,�1��ZDc�\���~�\�� y�-�d�)prIh6�x9�4-�G�ms^ke�~�(cb��P�U�`�������N5�����V[X��:�uᒺ��2C��:��h$zs���Š�?Xܒ"cw�����e��b�@�AUC!k�d"һ��mc��ņ����*�/}�;j�Lg=8��3	^�z��?���S��3F7�3����P,왒�{.���||����9o\�U^����{}pյjGg5{��h��($5$hM�».��N��
Y<���#Wdãꄸ��;AZ�Iֱ/ة^.�=7���	/���X���Ԧ�"ƺ��)A�̱3����崉���©�5;���,|ڳ��ʯ�c?xĊ<د���]���9����շ
Q24{�{�;',uf�v�TG�̷�0P}۝n�i��PѯM�9![��1��'%��nO����AO�z �;�v����e�a��Y�q�i�	�~c���_	�`���Arii�����F_6��Fj�Q(N�- �ch+��<���[X���G��5�H	=.����QL��{����6�/�Q!�hǲ�)�@J��U���Էܢ)� �ʚ�W���;?���M����AAq?n���P�SaU����*dǩڝ���/4�vH:.��uߢ���o�|����)��O��kAx�䡨���[ڎ�w��6-2�Zb�߀az}�jp,���Xf5��t��No��ؒDD��*�KNЭXD b�_2n����3�=W�W��x�\Z�mmZ:��}�U�9��oZ� g�t�@|�{݅�<36�`�V�מ�Vd`��R+�6�Fu�8�*j2�ؑf�EʾM�i�R�7c��!^Ҏ��^t�d���W�	]r�K��o0e@ �v�K9*
�rD��X#e��D~V51�Լ��)�ˈ�5.��Ii�7&/V��z���n��U�j�A_���kP�)�Ծ`���vT��Ͽ����%AY�[�i�k�ؽ����nJІ	Q�8��F9����ϗN0��T~�����2��!���5�O�-��$�5�c��&u��hA'oen/;����-�}~����p+v)�2�h��!�����2��u1>�S�(S����m�:�+��W�Ta�L����y1̞|����r�i��z�:�@(�뎩�\�|9�Jզ����a�s��Du\C�dJ��7u����	\�/Izp[��,��/���ͧ����:1�j��9K�ʺ
����Xa�*:��?.y�4mA�F\8u�����Wy�-�+����@�k��Q��s#�u6n�{�/1t0�p������*��G$&�H���e&�v������_�?�t�a�y]������㳗ڲ��Wc܇N:PN�Y͗��	]O|M������	{��T�W�5�2�߬���􅳴��}�PC��m�ϏZ�b�=ɼ(w�&����d���"c�?�=���&�;������^M��m����'gS�]��*�?u�q���$�B�<��8։����A��jm����U�v�.��k���/h[�
-0,�4���k>������Ih[i�5�"y��x	^
��m�ù o��V� 1�Fl�x�a����� ��E�Sb�\��C�E����`���}{vEV�K[*� ٕz�f��b&����}GOCa}��ۓ#��f Grޯ|�H�q'�I��9.L�2K6�`YV��Y���C`�'A���OunE��P+�R~X���zt4Km;a^�a�(V��l�i��xI���+�
b;P$s0nM'�ح���"�1{4i�ִ2�nO��}B���3\5����V)��6Q���M!G7 T���7]��aO?��I��v<���.f�.S���'t�Ff������� �7���#���������r�~�U��;B/�2��m��$�{ Z����U�A"l��]#r ��[�;;����o�Fa�#@@O�mŮfpv@�bJ�߂_�8XF�ЗP����n���Rb@�~��z#1�F3p�x+�����$��3��ѐ]ZRo\_�l�]��n{��D�v���`��8����DQ� �ٟ���x2��S��3hI���B�6�B�V��p�Q/V��:�M�C�1^S�T�J�R���H��'��-�G�+Y�i�Bsi'_��0�_�_LM��� ���ｕc2��i_� �6n��H���Bk�k��!��d�?��I���A��S�<Q,�7�l=6B�iH3�qo�e�����]*��RY�y<w#�G��<����:�����5U�C��cȤ�L���%�¶�+��-��8Q:��W]ܯ�����4���C��ˁ�E�S��Pz�ǧ���^��$��_A���o��h��j�e���1iVm�&Z��M������Ptn��$�s��zǓ�K��&�'ŀ)W�.��Z��Mdm�(\1�F�'����/UY`�d�1i5��������m�0*��٪�ǂ��eb�՝%��+��MR��
��������!i��M�cf��z �ßا-���O}.����s�d�����.4�$��O���&��S��򠵶���}P��9���C��>m�ό;X��
��ٺZ?�x�m񨣬��^,��r���dK��\�A�Ge��#E����
�X�6�E�U�	q <���S5>qO��>&�o(�p�-�i��!֑�S^�����U��6��|Sߏik����[�����(:�8.�:�7�-���@��Q��Q�P��P(N��g�Y��`�K���%X��9���z�Hdi�$껓�z��D8��	D�v�K�Z&�^+^��_P��w&mr��awj�֍�kE�8�r�~zQ�}i�ک���D�pG�ߓo��ҘX�L�i��텅������k��Tۢ���vn���@5�e�RQח$��;3l6��D1;Qe`�B&�/�|O����"�Zm�����{�hƑ�_�'D��H+��JL�f��T�pݽF�
��q��}>�=%P<P/B���bv�D��<Y�%�ۍ<ie	5>6����X�3[�����tNN0d��?��4���K;{|�"���<g��@/���ˈ��CM���G�O?F���bjS񗏩�~2�J�n�CH �Oɝw�%�����9���n�E��cq��Zۧ�жkL��{��2�x���]K�����)�?'*T����UZ/�"�򍒀���ayW�A�C�v��1��k�w'L@&'v�'��J���'���}�24�����x�S\��Ĺ���}C���ݾ��Y����c�<�3�/��UB�Qb
�悀-Ӄ�<Ȱ�mU�ǋ��fg��� �+��k�A=�X3��v�B%��[�4]�b�˛�p7A�1��H?W>�Rza��9���5�����-�:�n���`�����
�h虸KS��=hu�*����V$�MU�MZ1�l���̅�=�I�8R�Ԇ$����#z�����*�,�M l��N��=�t&vB�^��RQ����j�#�2��.��B�Zx��ƻ���Uu�oaJ>V����ÿ�DZ
W�7V����u�T������a����y����	;Ϻ���0��q�:����ݣ �0�>1ǟ���@T�>HŃ��R�l1x�G���"��œN�
���cuU����B����+�ׂ3�,��M����p#x���W��'M���J�ϐ��D�af��nlz)�^M�v{���o�m� �������t��Z��Y�X*)2w�
q��mmM�������h�
HL�U��"�Y��)G�8�,|ӻ���p�&`u�<m*�y�g�^Z�1�`=1�q�x=�뽚~����%t4 ��g����|\%��9\	���n���prN8T$\-�9��%��*��"ޥ����pι����ז�7�K�]+3�Z��߫;��b�(���A쟩�7� ���n;���� ����p�u�I���� O��+�z�����<��D$��8Ɓl�܄����(��:�ȗ��م?3�x�k�
��&������y�KE�]:Q0[o��ih��A�t�4����"xdh�$|*U0�YH�r~3E��Z�Ԛ��5�.fwz�3�sb���Pܣ�Hl1��M�@bs�����=y�`� �cS�v��rR��'K�1D.%Mu�L}Sִ�0�P,��`���]��Q��jQE��hF�ς�������lde��5@�YU�Dd3j�>��Pt��"�br��5�[.�>i�?7}�wsBM%^"#�L�@����v�R���$!��;E�ur s��%�ه��(F �o�e�;�?_f�'Wn����8^RUӰ̜�+�!20~��o����]}�(�.hl%؝Wik��o�"	��d�O��K�-ǅ�߀����|!��� �q�(�F.(��]�weD���ƾߙLI��L����E,������>����ـ��m�T������}a��{T�[�+KOy�� �*���иʊ
s]���U�OX��!�����_�?�l��XP`�m?[�хC�ʫ�)'i侈�-qD:��E������q���zO0ѳE��Q����i}*�����l�������H�]@y� � f�Hh㓳���Z[G�WX�2
�&*�1"���U���Ȼ�������Qg���oI�)1�����ޑ[2^��iK�F:�N�u��Y�?&Y���ܾ���!b��6P��Q�%�1�/��K~A�5R��������D���k�Eh�Wl�v����*UәC�恪����*��4�j�:�G!���Ai�H����̡���L�mT8�E6���+9�V��+ o�[Q��ڮ�!uښRXZ�d$3[�u4�ż��<�YS�.�.6��=$��$,���$����8(R�O��]m$����,��a#fԂ�#�[a�B��N0@J`6�b��^���H���N0G������n����*���KT<0$z��Z/���Cr���a&��*��⺣c d�E�hf��NxUm�|xUX�(�N^q��uM-��h��9�{�H�,�O�F����o���>�7�x:�O�B�Y������T�:2��%�#)��P!�1��z&m��b0+�VTŭ�pjT'WI���s΋��T�!�$���w�T��Y&�����/���߇ڱo���P�Q/�|�z�%Ŗ�n��
(k��ef�K>j��~9���vv�p�����%�Z��o���l��נ�1�z��.�_o�EҺF-�FA)�	��5�b1���ƞF�[!�w�V�����Sq�����MSsl0	!�e?���������1x׾�7���a��D�Ij��3��ߝ줫m��	Z��`�n=o#?�GjYWD,�f@��X��3T��a/��^�bs�n�F��qT�-x���PS�ќ	���t��[����0��&|K56M8�(#���e%iV�1$�M�&\GX�՞����k&�����>�����ώM&.][�6k�S}+sP�J&3+�J`sPX8h3��R���򒽅�A��/B���<E�f�-���mm1���s� �9G2��x�t-Pԧ OK�����j�ȧ�ȣ�N��NZ�h7Y���?�H�E��e�)�^w�_���G����뛒�QcV����R'�o9���Ԁ5���˝�0�ɻ6��ͱW�'�bHv�w�B4&���� A��K�"��RI�_�i%�`��׉�=d�U���"��ʵ�oA�^p>�Dxޠ@b����H��|�Cdj��|�O��sM	�Mޠ˛Ʌj���I�P$��z��祣��x��rC�����ƽx	̛a�l>�}���5/��&΂���17C�C�ܻ��^��H�/����]٭Y^kc��qgp�֠�.�[ư��W��&I����k�M��i��b�Z�gOK���K�ufs��\`�Ų�����j�Ug!+$֢���U�/��%�j�n����l�R��?���.q.� _"�.�����q��Hs}��z`��d�}��d��b���>�,����~�4\).iH��I@>Y\<�}���+�О�Y��V6�W���o}.UNn�0|B��X�=�E�C�6_O3c/���W��C�C��8A��b֨+.�R��w>Q��&�\uDx\��u}ft���3K�[�����<��/hɧ�m���N*v�aú����m9�KJ��9��JjN��4=%����n�C��@�S�A���)�o1�C,�DY�G��L�ړ'��5lӥ�ܞ��	�+V��y�	���c0Ѷ��g�*ߊ=DJ�Z�Iʴ"���`��$�L0H79(�!#�P�|@��>m�QBsHU�s�~[)�����<g���m9��~�ۍ�h�<q� G�K79AXG�U֦�~��B���Ӌ��	����Tjq�=�C�d�	��PR��n��UC�L�Va�U�Qsye��o���2�6}4+�U_C�V��X�#3}�������?߱�;.�E��\*C��0[����A��쑓� $��^3��O���  	A�@.�v�J�*��V]��ï�Wr.8Nɓ�'c>u>��kG0b�Wdb��~��,�7��o���A5��cgf�!�1}�*�u ��������lT��I-J��cN���q����"_+�J���Uh��mS��v���'DK�{�{�G!i}Sq�;�K�3{�PZB[��(c*F��һ,�J�8�7H��^V�������yɎ���y����=�f���W
ȼ#�D�g��$n�o�@��+=J�P�vN�J9ծ��d�����v��\}�گ{�o�zUsȇ>b���0��B�
�d���Q9���I���3ۙ�鮪2�=����6��܎K�沽-�!Ax�kv�E��M��L��cyxw^����dQ�9'�nuJ����y5�$Ê����}I�Q�B I�o6\�׍����,��$vz������� �'>��I͔�Y
�e�)Gc�^�A�7u�L��'A���7��(yz0"��O&q�7콘m-�# `+&��vA��߀��uU�N1H�g�Β�F����ry��#��K��W� 2��o�j�iQ~o�bhc��X7C����Ȍ�
�n�F�zVvM�Y���
Sfj��>�\�s0KE {!�n"*2��Y$�-����fwW�Lv!2;�� JӤ��\2�"�"a���vt�ɸZ��얪|���e>�?����V��A��(5��M�bJZ1�`k�y��V�P���t��S��eS��90��|�k�5_J+q���i�<G�;�$g������੻��%�h�X��χW�
T��E�� ���T�^��@@j��υ��uy���U�`����h�ǚ���e_���p���lJx��a �@/Lm����@��r:�f�m���V���ر	���#�Ċ�tKT�C�������oC|"{���g���m�@��<Y)٘���U	����)zaH�z

zdХZZjPȁ�Ǻ����=�l`<��`�7��(8�?��mFuk&�q(�S�5�-��[����4�Gd*7�ә� a�x�#� "ٰFBR:�h:��O�s�m`�w"�'��ٳ{�sYg���y����b��u͒�#��w��!��s�lF?u��,~�&�����H?�+�P�[$H�V���9�����CupE\���bdO~7iI�h�t�KC٦�Z��,�k,׺�O@H?!��7�T���>��Ȳ�-�L&ή���y�z$��� �<>���e�4�{Y��sb�;�GCβ�
K������y�)�.0�;Za�{W�hu}���ej_v;�(h'�di�N�ػ� l�H��@p�^���<�׮]iW,r��|���M��p�9񙪡7���~���ݩ�fL�kMĬ��X�[��U�K�O8�r���9��c���N����2���|��9�q>�n�n_�y��Z�]wk�
j���X2#ߠ�s(�<�UL��cp�R���)���G����\`�sxp�G]᧫�ˊ���X����
غ��M���}A
 n����"��l|��Ýyx�ws������ƣ欘�5� �=<��T�V/`OWv��^��g��o��>��2��V�P���R��*N
��;���e6L:��vh��L�ę<jVR�!m��<�~�
].��:�̔w�%�b����;*\
��m���T�N��V�H�j���{eBo��v���~B3P��[B�^H9�.��l�Ȳ[Z�,��N�^9ҍӷ�s�r7R/d��톄�������;ս�씴м�'X��@HK\6)�V��(�3O���E��� ;<~�6�xg<P�l!"��ޕ�=�B�Ha��2����� 8i|2����e���,��R������W�K=�&�'�+@N��E��vK�B�h�V�C �P6J?p������|-cA̩����^8Ӥ�L��y~�WP_y����Ș�xZ�2�e,���7�������	[�/!�VxOY*14x�5�zw�hE:�AԲ��)���+����Jft�Z��^��s���ILf��6L�=O��;.J�M��~�_(�7m�s��؃�M�!�� �yG=��Y�Ḝ�菪q�S�օ_�L��Ec�_wk����x��d͞>h4�֩sm ��Wo^���X!�/s�_�`+`�ƒ=AU���@R:�49��#%�V%���f���h�u����o�c��>�!��%���Ӣs�.t�ș�\�%����$$��3���\U���P����u�{$<�+쨎k��%<zO2���U�=z��+�JK�H8F{�ߝrث��(��ENNS�)�b����E�M�4It��6_B����^<r|����{z���4��7l�JQ<�زfMh������=5�0���3aדS�xJ�;������è�;(%��rDٳ��jkb� ��B�v��7u2�׌A�.	.���m��.@��"+D�y:_����Vu}�:7��y,���W����[;�k[��!���� #GA�~�������ݹ�k�o�h��v3x��"v���<%� �[y�"��-��_m�˪��SUD.�W�Bh�ȩ����yO5SY����]�~V() W�!X�Flh���r�uc�� U��{�������u"���bT'�n�M:+���?�W�;)ӸB�i�=ۑ�����a!�/%��qI��sx�3Ywn'C0f%��><�;�sD�tّ���(�m7��^*l���K,�v�8����y�!���T}-�.w�Alm�N�̿����z�&Oa��"}(4�M������AT��A������	�$#�j��-�����.��;RLZ�a����[1�͞����$�{�b�И@a/�������UtP'�%/?��[���_ �<aNtP�#��峃"�q�ܿ�@j\^�ӵ��^��h�Ng_��*�;�Pp��5�r �1C]=3�7�� �J�d�T�б+�/7k1.Ӆ �A�����
ݸ���=���*8S�ޅ
{�a� _�r�3a�1�v=��1 5=�h�l�n��(e��V���B�W轉�l��!@��!��ږ�-�7�˯W�g*H�)��ѦT8�us|�O���^�����,�rf��BAtTXG����:����
�_t�?m��14T�k'��z-Τ]+V���;��k4i�X]�;�z��ڂ�����߮d�ת ��Q⊗(��4��6 Z��,�������:�|Ri.
�W���qGU�F��,i�������/��(h�8LEj0�P2��E���^���J_�����{�B8p�$HZ17�2�
���@m����UOW�`�N��v�M�_�����S�S�5���g5c��ȏ��7�3��p� n65��:=��/��lcQ�N6�d�ˑQ�p���E�T"~�_����ܤ�
Z�'K�G��RiGa��.RԹ�"h�^�����I��ˡj����U��A=���Ag����:׵�!r�&,�u�ezѰǔ=����I�U�BX�o6����)�!K6�|�TO�+T�D���W�c��x��0/[��o2ӈ���6`�`R�5h��zS�c6d�9�*�\�9��·��rw�z1�PhJk���s}���x�G��(�.�\W�^Wzڐ>Y���;��|b^[�������fN�4'��6͎���Y�4��䱷QwC�o�������@Q�G g�5��~���؊騤tt�=�����OˮD�d��z�?�VL� �E���y�S2�-sn���8����9`��]"1P��j:���8嵍C�P�w��xB�d|�����P\%1��bT��Ek]K�jb9&F�8m>R�"�BNXC� 'w������A�"�x�>�u\ip���� x�y�(i4z����3�ve�{k껰��=?��������ͯ@V
J~+��I>ֈ,�AƏW�m�l~���#]�!�0Xg�Ҷl"K7[��S���-�2R�����aj�t8h#�{l'J��䡂c�� ���������4�lf�N��7"(�D�ٲX�I䭸$dp~uM<�W#�Efm�頕��nk*�c��	���nK^Mm-rL��H-ZA����������f��
p��ۜ��^��q�����K��I0��kQ��j��E�WT�E �m�DQ|b�oDI����z������Ӛ��+���|t�1���"|C�.=��Z��W/��c����Hf �g�h��#qM�@��mwe|C�
�	���HT�ԀWX��C�6ݸ�Z�D:eE�rϷC�-6�2���<�ǥ��pj1��P����)�ϋ^?;n����P�Q-�V�~�R��B�%�v�)B���}`!�%z9�^&�+�O���B9�<e��N��@�+��'6����\vt?�LH_M ��L���M���g��h��Z�"�]��lȣ�"�#hi��Gp(0��5ޞ�����0�=Lж��2��x<��߅�J�/������9^����eQ���K!��w�_�|��Ƥ�jU����h�O?;�n!��er�٥��������핓��N��Uh/��7���'��Rd�Ȧc�#�Y�ٴ^M�'(ɥ8�[��'�A	~��}�$L�헝����`B��{mby*���TU��V�j��AB]��{{�x� �ya�~����)=o��Î0�x�i�w�^D���o��W�b�䒪O��?���⢿��VIoSm9�͊AjF��f���pCM�ٱ{f���/?h�c"��D����o��V�T��ė��(��&cVa��j	Z��2Y�A�y6.���4���lBL,��	�^�&���k�������g�kQ���;0F��'}~�H�y )~!�����,f�,������x��!Mv�L�ś"rf���O�u�9�G����-�#��'ZO,�$]������R���9��{�t��w_��jM���Qt�y��#.S�_ j5û�
�Q�9wn�s��J�������ͥ��@|��:}��06� �XC�
�fE�~%�~��!�]��3͜��"��(�nc����_Z��~?s`~�j�;:�=;H�o����t��vW���ғ�O�2�p�X���unԕ ��\�49�"G)�J�/N��l<)���ڗѸ���_9��7����ӷ"t��ק��~A��p?fC�`����&	�R�H�Ί�j#��H��,>/�����V�!�e�;&��G��wD��x���e��fE4�їԛ����m�#rg8� v\e�
fa��{b9N9�b5���Ϛ��"��ڏ�\u��&�� ��;)P$��j\h�Ѯ����S$V�/�RF�N�/s��BL�B�����F�2�سW�i�~G��!�-���CKZY1gG���29_D`���A��8�����S�B��k��n�|���m29E�Ad��j����V��x��o[z�i����`qh�{�2.���^0-�]�����E�ʢ;9Q�! ��Ki�ye;̖��A�&�S���9{�Y�2���Vn��/g߬�ac����_�D���.B��	�q5�n�uB��{��Aл��~ A�Ed� �˖�q�(WpI��Tы��w��J*�Ш����&�7�N	���L�!|@�t����;�:&)L� N���$�e'�MM3Y[�Cݜ�6�~�**9"���8�>ԡh_X��H��>�U����[��5f�X6�W�`�.G�y<cF�f������3��1٢��I�3q�ȝ~t^����y���XfG���F��]q{$�㑧�%	�o�i_b��wMrYA���[mS�gW��U~>��י��Py��Ԑ�^1�@�p��ҪCe���a�t��\t?E��M��|V��0tg�B�@�<�(�z.H���K��w����)+��c�^Q{�0!f����.K����彑F����Vt;}|�bٖ�v�Β�v��d|���Ǳ�VC3����'9�����Y����,[�{g�.~b���m��K�1y$Q�N}a���U��s�)d6"J����#��W�<a'�II ��L���	F�\·�{T7:�8���V��W�b۝��j���I����f�aP���6��<����|�(lS���Xˌ�lvj���g�����	HK��+ƹ���@⻚����@dڥ�W�5��'nߪL!�.��z��1�Oa���1w$1'�H�)G��(9�)xed�C�x�E����v`n���
7fHXBc��bb&�^��7�90�6,{�t���a����~_sB�h���l ��e�4�|�OxeB�r�T
{\&��l�@���C}�n�[��v�I�D��晬Q�Z@�����������JJh$D=^=!�N�TQ�=���������V&��8sJ��QL�������_ru6��6��!&����d�-�\;���*�v�C=d�?�2�n� g�x��?2���k��^x�S�� DRB�.�0� �㪜�Z��V�l�&��d�3�'�� �¢l��/�3܃DU��"�Aߨ̱���=zi�*�h&�����-�'�+J��$���S���F��xB��-�m�t�P``�f��'��"�~���J���׼B}��Py����+��lԣre�*B;rH��{F`@Ja���0s�A|wY��^�Ԃe�[m�� n��G3(D��AC�$9��u�{���LG�}��4qx��
 �_l�2hd�x'&I����b��-=l�^�4�"��Ѥv��~���ZS}�/Ф�����]����U��h�"ց=��Oq����a����n���R�N4��Ϛ={ή�(���'z
���7u)��W_<x�m���p�.	S%"�yTz�:�u���)������K�Ch�����+�}���f��/����g�sO0O9��L��3gb�bB���_GWc/�԰���d Pi�f��Se�ԘUӦ�E��nd��ob�xj�Q̈b�TB<q�i��3l��8aU��wힾ��S||8����C�cA�CKA�z�J�n������Xj>��!ܜ�?o��' 8�T(DU�>���-��6 ��h��\���b!�gf7M��}	p�9}�E�8N"�����|G�3��7�)���)Η�s#���'�VvQ��%����,�5��Y��s� ��{�ط���d��X���T�76�PE��"�P�ꯡ��1��3�i��C�s�Q:�.�2���!�Ŗ8L��gf��ٴg����W}[*��$�V�G���ۉ�	~�~�+N���w[�N"��?�3L+��>q��a~���?�\���T\��6T&�yۖ��]
�Dd�������FU5}0�'�x���P��KN�6�T���U7����C�����˄K�k��>��WEޥW4s�8�4���A����&ԍ��Qg���
K��@?l>��6-v�w�GQ�K�q��
�T��|PU)
K���V��C����Jko���c��+jr�����+�a��I���6?y�x�
>U�8�m��+o��~j3'�?U�}�B�;/�|����Z��V�ɐ�gz�Ƞy���$G�c�~���U�%j�۳����|3�B.�1�hf�%��Uw�_����)d}1z��n�i�id��.�-+0L��ZC���Z3������.ښ3���h�2�Gn���l��N����<<�Жo��tGWEK�0:DZٻ��nN���&
�Y�3���#H�`��`O-V9��Ҡz1��	\2Z>�X�k4�L|Bx�98LlYt�.��܈�k�+��qD�o��ᙻp��ei����s�ђ؁�(�!����r./�PV>*(�]��"r�_�]���������?n�\�W��ھ��8"�ߖ�@�Mn��ZM"P��˳e�9�`�n;��!pX�_&�3����Ix��gV����"P�y�OwY��_ip�w��x��mH;���m,H�$5�c�M2��Uogr;&ؒ���ţ(�5�9����XM�������?���Ƶ����w?��Y_9\W.��s��J�Y�Dp�	�������
�����Lȼ����L6eR�ː�'3��%݊�kY,���wɫz��sC�3n	�������2�q�����P����j����W{?=v�_1������o,ͤ�!�A�W]5J<E{�N�T]��Ǯ{Z�A�8��\F�_k��@�ԳDѳq�
Ө��?�T�����g'&��~&Ac�����d�ʘ��O��>� ��־ ]��ʶ�"j;4	 �3l��$��a���z�Z0�%G����I��J�i~�/��d�DA<hb)�V���Ǒ�]scE�-rFI���n�W����o���
J���ߢ舔r���xf�إYUFU"M�v�P���}X�z���!ϋ��'��L�++���Ţg�V���Oxg���|"ʲ:)�Z/��:�;/����ɦ0�{5�+�������'�����4�_�#p��8Y�x"@i�F9M���ee�\Hnt��b��r!�A�%��^�f�	�*���3K��Ji%+��Ň|���m�2V��� Xݔ|}��$�>��K�#��/��Тu"��[����9�����R����S��|����	��ۜ�K��+gl�����F�=@];\����DU��^I��%� :�->b{�%_�BĐ��Խ4��~�40׮�/�v���>����Xd{��j�َY�vΞ�F\�M��@Uf��F�P�+1#g�!��\�)���/+S���xI�
��%�z�aɤk�"7���n������TI[����X�~���������Av{zD@��1J��|���#�^�%5I�%�$r6��&z����^|�^�*a���T��ʮY\JQܐ{��mgs�;pMbi�-b��غ�3kgZZ��5���H307��h��<�j�3#f��}=�bo�ͯ��N����#4rx����_�M6(���H�1�3W{2�i��+�r����m�v���>�zv��ش1�-��/��2��8�/شb�qo!�Z�ʵ�Y��N�"�Z�>W��NI��pLL��Y�1;���G%�SSR7��5�����qa=�I�^Z��wE*y���ket�!z�ؘ��,u���c�n܎ ���Iq&K�q��4gR������0l}',q-�ˊg2Q�ӹ��;��5�HX�wj�� �S^I�������+��q�͟�MGTYd_�G���V�IU�a<rm����i��a���
M�E��IDj��P���$Ĉ��Y�����=�3�w\;Ի�X�D>w���p�K۲Ex��O�
�� ����0�W���@�U��l��0�̈́�/ ���lG�����	k�Ԙ�N-���f���P�Q�4�[g�,AL�iI,U�=�4�`N@�*�[{�̳���8&N����j~I�zT�p��������'���C�hȅm������~�ߡ���mD~�ԣH��ԭ��Ԅ��(�� �����Q��+��@߁���
*���,t�Uq�Z��Lw޾x�]�πW���ߤF��7�
�ze����
|�d�!U;U�x!{�,oPa3JT�����8�gL�U��5� �'�~)��	���5��X�L��P��	�?߅m��'�_�5��=��Kt���ߑ���B=�t�ܧ�ߛ7x%qϦ��b@�l���@������-ϥ�Q=���꼨���d>J�hm��\�g�ry�s��M8���d3�?*�@�Or�߁�Xz�b��aex�3mN�/��Yl0�x.B�B�b�U����]-\2K��	.L�u�*`���3��T���
��>�0�ECwլ��'w�2����:��=�<�I�G5[e83�֡�7;�=�l�����%���	Cc���A\�b��V=52��s��5�9L�z����~�E;��%�u���-�M>�A�U�**'O?�&��r}Ǵ�4�r�`�6�Q&�-�ٗ|b��e
�k�`Ա��q� �L���B#@m��M��jM�e"�H�� ��|����s|I�c�8���Z�C�ə��OH��hY�$'����`����L((u���w��	��%��;�t��
.,���,KǕ|�~��v�;ϔ?~�%t�뙘|uLRMb��wh�!:6�V�`�:�������>�`cx��9T|jȺ��kOv95P���(�c���vL,�yԈ���f����J�|as��3Dvbۙ쩢�P�v�kg�`&�.�΄�z7"���j!������+���t`�xh�y�:k��f�[�����P]E���ŬvoX�.=�[�iy����ŐǎAyw�l��2�s۬++�d}@d��D莴�;�&�R�E���q	ģF	��N@j�q���;%>o
���֌m�Z�I�)�[+�U���bs���2Q�v�x�)����7��D�ZU�'q1!BEC�&��sl��?#�ޗF�c!�U�������N̹kM��gC������M���@Le|/��������C�N�~�bOC�d
�Q�#����ꑍȝ�L��}SW�ݏ��4�"?�
x�E����o�3�['w����h�NH�Q����_ۙ=̓C���q���)��5l3}x�6!��VE�<����G������q�9t�pk �����Z�(@P�1��R��5mBC#]cS���/Φ���)��3�?ʼ��V��X�g�b�
<���>�0{�����]��w�5��8�P���{���¨vک���Jcm���z�B���T�ut�d�r�X"g���Wk��>	R����2/8�Qp&��k@d���w<m='h��?��m{F��ìP �2�"�	��5y<q"���WO����ߟ����7q�����'�v?�����Z��k�L��0\�i�Z�:���
Z���V��u̔�)�u�
aHZL���ʽ�A�8%���VܛD�H�=�v��db��R���$�S0��1j�������lɑ����7_&���NJ4H��M�33f�E���&~'�F�d2�i):2�d�M��
}�D�^0+�), ���g�2�|��,�Lp� 9�iBm*�ļXy��`L+:,�޲�����l?�fY�c2@!�I:������ix���'�"J0�m��`(>!���š$7yŁ\�v�i[;hv܈�Dcڱ���e8�Gk <m(��w��0��f�O��;���oG��OpZ�7_S� ��ο�F�$�tù�����IF�>0���+�qZT݋,�z�g�}�z�A�L����F�`z��A�k 	�Ga#&>H�L���V�J$��.b~{�͐e���A\Deo&���Ŏd9�U�h"��,k�ٔJm
����V��۲����^���ۡ]xǤy(�VR�\tiE�=Ɍo5I���ԻEӏ�>a��5L�±��C�/�V��o�s�,J���Ze ��-�k��C�q���?IePx ���hGi[&�R���{��u\�~ԟ�QP��ƒsI��a��>s>}V��Q���"�`�*��>�1���*��,Nh�=�kE����n��<�TR�c���='2���p���lz�	\��AB#�4S�0�FM0�m���LBg�!r���s��xPH� �i�>Ġ(����+�!�i���
Ȗڍ7�{���i|o`;	��_�`A���:/Y���߰)��'菺�H�g�C��?C^%
�Y� ��&T/!�W#6�٨����SO��&�0�`H[XbW ��P���F=��>��nE���pzM.u_�)U�G���G����I@��5� Qn��1^�������r~'=>����ge]�X*�g���@q��m(�H)�HnP�WЮ3��ed^�����(�oa���5O��p62Q������Y�_lG��7���X���*iOHy�\�ct^�߃+X~��oc�f��V���y5�X.1n��v��Z���rv�/�g��K�������O`�3&������/8}�R%A�XI�q��د%�8�~��C����ŭA�l�<��6��Q��A��e�ߕ���3��l��%�5Z��6��A+��OX`�i.C$+m��69K\�@�;Ц�4��j�H�J�R����Ov�����x������Y���!�-׍�I��$�hژ�[
��x�"f��F%��l*q��>���\?G�,����U>��X y��J-t��}�^!�����G�َ�]ĴE�K��xe��c�#ђ̫��{o�
��'�o��ej �?����{w]��ͩLP���	��R�d	"Y��˗C-K��=�_�	e�N/����׸*k=7�/L�Q%!i�?W����2� ����?�q��Q+�E�8�u��^�&�n�(�*�|�
V��5̤���bp��so  ;b����lߥ�V~��L@JXs�T��&�BP[N�#�^#�[�*n:ٍ�G�^!���9�S_R�D��>��^��],eC�n��3Iuw�|g^����V��۬�QT���2�OdV���L\FMAc��ޣh�����w9��;<d��(�nj�8t.�z�և�c0�+�e�9���ޣ�BZ",��1%�~����ܗ@=r�KZ]�ܓ��z��Ƴ�@��p�}K��i�DA\�ؿG	MU�!#�\jW0'؝�ވ���n���(��6�)�(��$⏡i������-�R-7�Z��7�r�JG���Cz��T�6"�L��r�F��ѻ#��|}��W�˳��a8֨�~�R�����D�;Z&��B�8��l;��"Q�߯����'9C�i0��,����}������c$�̚�O�{Վ)����w6/A{H˽U���e�����������Ndy�0	�$ 5��z�P��n0[
V�(���Q}��tR79��h���q�>�iIcdt����Jz��Jm����ܮyq>ae����YS)� 5H���e��w����Z
p,�С�h���}6Cz޻J����\� =��(�Mr�+L�9#�	W�Q�iN�]�0#`:�䨪{B=/�!>��j�aɾc4b*)e���e����Gn(z#����G�Q�}��2&�Tx!>�BѢ��6Fi�� �%�{�[lV �B�QB|�]��#�Vb��wh4�?~.���8�By���W*_Kd쥭'�1+�>��l�����ȼ�f�(�ڧ�T;b� ,|i�MJze�E��"6G��+�)��CM���d��5��6���z���X
�<�8�%bkd��'7M)�g��\�Ǯ�,�@܎x<��#\�R�z^��+�I�wl��߸r��S�rIgQ\����O!�S�Վ�fS]fB�1�\D��C��{>�\�:�	Rņy���A���RLz�<���������|_������qy��0'LJ�8��U�z@�,�Z��b�����T���ֲAĖZ�Nm����ZTz��JSy[KOf���\D�;q�����p��v4m��6����>#�}'��8�8�c��
�9� R&G��8�O���b��hC]�$��)�P�G5�0�P�䊑v�/%�!�Q�<83*��Q� �z!��#���P^پ�!����w�T�N٢Q��T�%���>�	B��+�$�1%��]��n�i<H<9�y������OA�>6%����z�U=$�V�j�Ş�sN���N���r���>��uw��mBι�&�����1��[
c0����|X�� [�t������i糷��I��lղ�H�����1Z�� a0>��v�	W6��TŁ��n�L�Mػ���O�e�<r�}�)��/�0�f�����҈.���)>��X����~2�B�aap����
���}�����f�8+�8¢
�㹀5	�;\}��P���A�C�iJ�P��!��$��}�����Gwp^��_!B7�s&�=i��AEt8i# ��
�Nyv���U-I1���3V��O�#�?�m����ՠ\��!�x�/o�9�v-<�y�8�3���	�э,�V���������u��|u���=��3�"�� ����-5�F�;�(�Qk4���>-���5;#u�%a�OTne�+H�yps�Aw�\~�Ê�vF�`{d�� ���H\JM��d�i�m�~��p x@#�5�(�մ�\��j+[�#�$�{��Q>��x�f�OѧP�jZ��MiaL���z��-˗JҴʰ���ז���}�HN��'2+/������N��<��l��i�zs NY<�mXt���<����f�k�3i��(S��V?�I�W	!PxH��}�3��\2�؎u�{�h)����/6��Ҡ.� {n�7F��J���%]��K�I.��Z��J�?8�;��������K���/ȝ@���U�{���u݋ڈtF���'H��o� �w������	#,L�Z����������,��aK���:C{^��S�-�}��r9�J�Fi� ��� �Gc�>�섏�=��Q=d�^��64R��\�1�4�¯�&:���-뫏� ���Ñ]>RFB�'���������#/�<�1��0�5�� �D���&~�",��&�U��l���4I֖������Ԧ��p)��=~���N���+A����ם��!�'n�u�:#�%&��<��!@��X��"�Cķ(Z.t_���I��-�ҍ�bDj"A�����s�>�����p�˯���Ckol)9m�!cuF	3�s�=���G1��B�HՋJwwt��@�.s���?�����4#��M��n9ܰt`�*d����E��ˎ�xU���M�.��ѭ7�佸(�$�$n����X?D��*�5�ً��m�֊�`��!��l���("fŮ��?�4p��Ąi���Y�o�n��N�r=d�(�q)�#�,�������h)�aƪC.�Y4�105�TY��0��7�����������Y	�TU!�-
�����\��S�8���mU��#����N�|9m��ZF�8�D��~dSy�ne*]q�S��/�8-)޻��o����<�qDfܹ�5V�咳ܫc��s9���+p���e{&(�U�~�P�`r��W,��^����8�h��F g��:����ȿp!�*��vїj}����2�k�Op�MI^ofhH�X,-h����kJc,EB�����8�Ph�ϵp�.���h�d�@�L�*�k�E�P�g-A���`?�26�̙��"��T��_o|���zJ����B�W�,��,VАQ�x��r��s++�\��t*=+=�^p0�*~3\���ѐQ�V��%fj4ak�7�I���bԄPB �)&�%s0��<�#�'L��������AUDc�������Y�h��d%{�u-����M%'.���9(4�{�[\?|���"ǆ�	�5�N� <֫q�/�;�����W՗�#w����z�ϗO�axM�4�m2�y��(=�bR	@���]֐a]�O��GsW�ޞ ��;֨�� ;{R�"��[��ekh|�gҹ��m)
~�a˗&N������	�k�M�DQU@x`�8i�_���獹��̬���}���<(���$2�Q��n�T�< ,l����_'[RC�0�kK���R�3z�~W鴫m�tZp>�V������MlM��k�_@��G$�HU9��*@h^��e�
 �z���趷>t��C��:�Q�_kx��f��!�QO0�'��2KU����m�{.F몖,}�x�X%�YN�=����UXqv@û�,�;����C�'l���!=-	Ġ���S�����V�>Y�Ŀ���K��l-2o;d�/�2���k�ifYp�7��a��O��֯������M��v�$ 37m���/�O�3wZ����1�/�MLψ�D�c_7�ܥ0�F<�m]��0�ꌎ&`�����Jw����Q!:nf���#
��Z��V&!y�=-��*��������]s�O��AKju��"
�]'�S���J�&�p�CT�Y�Y~�/�-� ��S�f����K[�����)�t$���}Q[LxXb{�f&�n*�6� ڊ�?���D�.���iVؽ2��� �ܽz5Hv��t�ΐ�)<����D�r�?�g^���ND�d��Qɾ�ZƩĐ��H�ͯ�!�h���)�B�:4y��9�T
���$�'#:c�=�:;�A���:ӱ�	=�LQ`m2Ů%��e_����"�J��f~teDT6X_���iarV�h�+�1G8� dW�*� �-\�1q�2���\/d��\J�}�S_�=jm�魖@��jв��k�゜,��9�7� �o5�xO���X!�ߐ��b�=�¹�����_<Kj��O@�#�q ��g��N+�ʮ0�s�W��Q����Y����P��%z�&~�-b!rƼ)iZ����Iˈ�oCDe��2�c�_����$lk�$(��0���qD���FR�=y�/�4��kƋV{%<��3���W�i��`���/c.k�>On�YI��L݈���p�ަa���1}l���~�C��Ɇ^�pz{��%�\�ȷt�iek��ɨ9]���X��s̫s�Z��t���� (o��_��D� �T<�t��j���{����\B�sf�M̦A%̚�9�w��gu��B��P��ߟ� �����T��Z�P]��2���D#��6DfV�����d�ܙ`M��������,�	qN7\�D|=�b�&��ვ�5��1`L�>Vy��2	m�/��5��û>P��r̃A��-rr%��ԟ� %�/%>�>�%>M����B��<�j5� 9��~�/��9���p�gj��Fwe�X����)����!������1@ٙ���^"�OCxK�;OR��4U`����d����,���x��_��a�؃:}�~d7���!D�t�
>���[�ߞ��o��f愴�2'�s{2�;fr&?t���~h���m/A��g��[��lx�$a��3�D^�C\;��w����A����F��z`�����N)<c�4��i�P��z�+�W�?b"���cPXu��%��d��d�9��$ �,V+���3ָ��p�\���)ܝ��[-�#����*�ͫfY0y=[��,�h-�M� �6:/�> 7];��1�Ѹ�7ʨC���I�޼}��2��V<�vҵ��I� Φ�<Ae�-�<�q��|�ȩ�����m0�w� � ^7�ޡA����&�W�B�m4!3Viq�Q�z
�	���S��>���uM�-`�Ado�Y��KB@�4������غ������W�#єȐ8s
El}�[����x�,;~��n�.N@\�7d�����Fp�� �D7G3QL`4��o!	�q*~�L�'aw�4E%����^��a_&n	!{��o��T)�Mo�B¯(�٦���0g�AHw6���I��T�P� �^���4M�9t"5چ|{(����{��G˶��+��O�M��h�ˈ!��K��Q�����`�{ѿF4�"Ƈ�?�R�Ч�܀mF."�p�Gӝ����h�~�	_-�*����;Y�eqr.���Dӝ�ݏ'�š��_浰�=��mo2&���R	����\��dk�;���^����GԉwEiP�w�S�������T_�x��88�? �;�Q�*�9c�*�:c��w2g���֮@֖Q~W����^֏��ug���_�@
yI�3�C��#?�KG=!���~����,N�����3�J��;N%W2k��>Uy`�^��b��麑�Y�(V:W����@uqOMB`�1��_=��\��	|Y�{z�H�Duq3�F^S�jW�{7��K���,$9����u;g�"�s�(�F~�]M>&���~_�Ӥi�y|&�Ó�оO1%W��s��;��6�䑤��+�ިV\����9�0���Y:qwvm�hI|�8r@)4�A���6��?���/���´����0 �A�}7��G��O��ĵ6Ƭ՚���D����"e�k:y:'4�6��()���/�������#�'-��-XjXy��ʬ�5���R,k�E����x�E�י�,�V*|4��UiԃP���@"��#5�Ur\"��&܎�!uW��=1����"%7-��c�p������\m;�&��wd!`,u���ۺ��-�Q6�	�h��sTsj!�}�Xf�����V�i~G��:�1���v*T/��\�j%��J3�������%����8��<JԲފ�bh�����"K��nX$������>�>yZoY�R�A/���fuu'[*y�D~�I��7�J���!ܶ��xQ2&3���A䔷�E��̈:�t�K]�+z�2o��Ap>�!R)�SpL1�������,��3��n����-8