��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�rQ��7%gN���i��v1��(���:m�>���D'Ͷ���tur)���!^���p�NW���^��I<:�E����Gd ���
��Wï�����V������a`]�e�(� ��$�z�K��w��b���L_*�Io��󨒎$�����g�-�A/��n�\�I�z�OB�\�)~������SD8?؎:�;W
�����0�Uƨ����z~��"�qB��ཀྵ��<��1c1���;>^�j���I��ɑVs\u�(�5�I	\ڷ9t� k���Ajj�����z�g�D�_�a?�K��ؕe�h�k�k�=j�1��d����$�ʟ.q��]Ԟ��:| �ﺷ9�����\��+;���{yK�!l~-sM�C��
h+�ȓ,���͘3A�T,Q���i�&�u�%+VY�JE��r#o�}:yы@k�T�g�������0�+w|VӁ
6��֖�n+��%.T3־�Ȍ��B�U�4�B����]�OwKR,��Lm���(.}oS_|�
�@�Ao
���Zc�k_�Kk~���U�� �A~N���4sO����������m?b�-���Í;%�M�D(��	��nU.Q��\u��� ���� _�V#���Wp�ӽy|@A;$�-���]2e(]� �@,R��b����1K��6�����	�E���޵9/����s�q�&��m6�������4��9�My���[Ϯ����~`��c*#R!M����WvO.��VWS�tx�d��5��������"]TV6!�]�����x�^�u�~�_��(KxG���ӁQd~a�(8T���t�bCA9�QC/�[ө�Mg�*aT7�P��N�,�dHa	�p����Gx�#�q%7��s9{� �a2h&���-�;E������l�����*ľ����Z��4�3��0[z�Wo���\�,d#]���(���n��B �9ಳ0e�xw��3W%
���U�'Ȕ1�0˳:���-��n�G0]�����u܀O����T_aCO�q��1h�""J�+�&o�����0��a�6,n����ԣ/�b������Z|�x(�яE��z�V�� ��!o�~���\��y�� h��־��V�U�RJRJ�+�`!;�̽N�����<��YW�&�"2*��Dmi7������k�&�?h����O�0�Q#���J���2���[���
م���{�-�q�S��cj-v���%��$+V����Ձ[3��������	�i�v��^d:��~�O��u�U�u11O�ѩ	�(�2\��o���͙$�x�h����G�����P���ҋ�$�X��Xcd��ןٸ�S����/�Y�Tw����f�=�o�g>�>�m�f>�{$>�j\[��I��䦾u�*��fL�
�ι� �|��v~c3��RYbu��W�XU2��-P�������iC# 9���%�U�Gơ�A'sg[�IQDNbrp�pm#lx��/����g�� Ɵ(�S���B=�H3{����H6E�����&�vّ�}�e>�k�~�D���#��~Tĵ�	�����k�8�����h�)3W�VD�s+�$�\�,ؑ�n[�{�fI��nպ��zbyR�e��Vf��3/;�sk���T���i��*�E]�aRE�	�:�q�x[X�kN5�0��.�c����	������J��ZPr�<{���:�ZXw�^��hX��%m�Y��
��'d������b��R�I��t[�%p�,;D���'E-[�oiK� �HX�a�_.��<��U�įdMf5E��k���n�a8��7<��$]�#��,8*D6��y�"Wn�� �r�ōF��擲�&u��N�B��J����ȃɍ~�`
^������x�L-�� ~����J�B�5�c;c���kv�"R+�gE(8r�i,��ؼFG���l��[/��> �C,g.3�%��HY�kU���T���WÝ?*Y��G+>K����y�2����(���kޭ*��`�����2q��G.�ɷBV��5�n�yd��9���%:����#���"u� }iR.����l<��%�'X����,��ңr{ ��8I���Ag��
�3j�/Z��챰�y}��� ,����"�ɟǺ؏�/�7��:o��S�11�u����2����2��pP@�Lz�z� &2�3 =*ʖ3��XW7�`a�UЄk��z,���h+.�
�^4����䗮��2�P�GxAW�b���{H*Hnw�;����Ҵs9ʫު����w�m��D!���O�%�i9$ˌ���:�Q�iDfY���Zk7	=�%v���E�x|Wd������6~y�q��:����frx1�W�|Ǔ�#;��:��Cmiq���ޞѵN��3<X��|� (ֹ|-2q�k>�d)�* �	�tc��j�)�R��͚�埅�%��ea#>c��Xe��iH�0��Y�CK5�A�?lu�lr�[,������yy5yr�2a�N���X�9�)�eeߒUݛB��L��~�kR�//FKV���- '���8�U��&���wY/Ėp��P=��9Z����wZq'C������jȴh�	�۪���o�����p�jF�13LK$�g�]Nc�|��z2"�^��z�^L#�
��h��Y 9����٪(>�1l�tȟ|JׂfZ��A����V���^���g޺�j�inp�a�P���`�)�e.8a�V�a���b��r�v������cu�z�V��H�^���ҵ�"��2df�[��/����+Vи*�f���q4��#��z^�LVO�EEo��<�޽&� w��k��C2���o~���DJwҰb���w�.�#E�u��c'g�=�3�G��P�G�%�5�#�֙☿��j�h.3bu�������P�)�_��D�|i$�o�1VU�d��˗�������-���-���3�u��	'�>�ffrvަ��D����^;]/r��
߸ ��u]7�U�a-cCL��?�C�i6�l/������'�8'�$,�d�_w2���S�Y�6ఴChi�b���\�7 c䀞7q�N�bYƁ×�a�D��[u��⭎O�LV��*�W�H�EPG,e�#�1S F<Y���:���F�����`�2>��z*0F��wN���o�mg�Ұw�. �B�D��Ԫ.��ƾB���ԋ��M-�>�5v�!����5�޸�+Mp%�_��gJf���&ԝ\[kD��&%��ekU���Djk-û~�{�bl'��)�t| �#�.E��R*��x}���"�m�y2��g�F����p��UfPA�hE�ٍ��1K�Ծ_��o�'�˼�C?�-{N�,p#���1����{]QQF��s�D�ӓ+G�˕��߀t�!�F=r~��˩W��bթ�a�щ2�Ch��mr�V,j�Lf�-@�,Lr����Դ����M#X35�qgc��-o=?�~M+�l@`�$�~�[8)��DK��3�}�_��2�����i�}9����Z�H'e�ܽ\�}5�X���e�O�˩�ʍr�G��Z�7��?�cs;�F���~��Ƙ� �Y�]6a�>]>�L���/�^�n�~�Lo:_�)ߗ�/@���l"E6T;$��;�~��>�	�F>��%�#�%zr79�[[����@��u�� 8�xփ��隂㬌��E�Z����P�����X��;G�~�տ�fjnᱫ�}�g���r��5�c�7HEt5=D�?�y�[�=C&`!�Q�uڒ��KIA`���nSK�
o��ń���F�`=��u�k������.�;��n)�.%�.�-�+O@�f{zM�e�M��gᑤW���əj����|uS��Q>���I�'/��O�	�h��:=݇1m���eJ`�d95�Sm����=(0���t�Q�<��pDIj�2�\v���>��l���k�����"Ih�,υ0���=A�"'^�I�z��n�f�"�Q�(���0[��0q��ю��p�Hn>!%EWL]{2��ʠ�x����?+�P�v��D�p�aO"ي���.���U1�o����0�$2�[sJ�'d_�,��HQ�b]�΍X>Ꝕ�^�]������.'n�Ĭ�y�,3\�z5�)6�L�.�'�����)�	�d�_-������n;1b��Az�0-Y|�����ߨ�qr,�R���0�&��k��� �ci�D�K��M��Wm{�B�n����2 
�{����ę`�1�܈5@&[�eY�WHTw�Ì�\��(�#\&&�íuٚ� �8�����l{�:��t��A�i�3*�lI��t�2a��+�Ʃ���4"qM靘v���(ȷ��h�C��0��p=�rBf2�nަ*�T}V�����(�\�p��e�ﰻ�
<Aq��TC+t�p�b��P����|e^�*S��+ 4�<�:�*��n=T�3)�%�����.ǚ1����ŕ�.��� VW_[;��8��������#�t.���z�s��{�d�嘴c�c[E
X1L���:���v,3��;�,9���70(�&�x���9 �L4/�dJ����9K�@
�q��-�]��5��\\
W;����q���YV*9Q�Y/��Cg�T<Iv]�%'��xTt��[|����*���D�tM�M�7���4��+5 ��H���S�q�1	�k��Rܠ��ě���(Sӝ��r�'�;n� �����/Z�d��*�i�:1D*�v���u�L6�gup����dK��"����ͱ�(2o �ۭ�F��,B�sS�L�]���?Oސ�pW�*cM��@�^=Zh��1�/��_�
}�x=�,o�4>�ݾ6=1�n��:a+�����q��o��w�	"��ԍP��C�d�E�ʸ���q��TLxHwX~������F,��kJj���������O��T�u���I���%@��Ѳ�x*�?��s@�0���\G�6z"\�{�8���	��0��56�I�Qnx���gn��
(��! ��a/p�7�*:�h��qg嘕��x$�S�V̧�^���P��S�~�����ڍ`�JĹ��G�G�N� �=.�j�hgF����G�ף�M����6�;�Pk\��~�E�Ӆ��9uo�J���J�����qy9�y���äK�.�?�����4��K!r�`D,�Ab]� �}��N+��ak���e���q4�9�4\����p�;����hϽ�J�H�B�.a4�cuv�����.���=[X�m.�g�-�X;pz.\�.�W�K�&D����x�	������F�J$`9�en�S�������܊�B|��}���>���hvJ1{}R�|m��2�dע��Zm��I�Uӥ</�4�a@*��/:y�@aj�2x�=�D�Z�!AFS��@�B
<Bv8���k�����EN{��L�Y ��?�A�"FV�����r+���F�/N�w�5��~@̍N�j�9���M��C��G/p=�5�~���Y�����b����/x��HU ]jhv5�E�l��ؖ��� ħ�����뭥��T'�����1��b�vk'!���Q�����W��,��&���R��`��?y�@{x�@��/m�c�w$��F�����1#�4�G�!bb v8��`�aT/��\hhպ��}j�N���UA�_���r�,�<G[_-BP2,���&3�"�8O#~��e��L�o�����̕�Jc� �p�q+= t��eY���.P�u��w�*v��ښ9�g���?jJڼ-�W�'��ϳif�5^��<���3y+VθW��ߥ<_��^+�p9,���V��~��3c�ͤ�M�/O�7���nN��&.���h���7�e����
�29� ��`�AOᬧ�K3�\�jg��Qr
�����XGU���rX��O�*!�-�|1��v63�k�VW�i�/����	h��%�-h+��.����q�%ˉ+�;����~׸1�_;����/��˘]�����
�}���ԁ48}2��e����l�^�k��99�)���)�&�љ�֏51M�T�r�`�J�$�Q��]F�	`$�O��ٙ\`��`�I�Ca@����%Z�3�P���&�Z���C洈��9'�^�̏m��f$��@i�}�����|
�r?/9�q2�8��>#p�O�AV�I����u�ɢ��`�O})�ZK��K0Hs	����-� ��6c��MD�1Ϲf�S@�v�V`r'E����"���\��}H��������K:�����3��D��0��q;�b�G!7㓛�h�����N���.��
�W��AQ�����,^��p�jD���� ��F)�OwX8:�Ko�
��%��]�����l���?^j�Ύ^t3��)�}iZ�K;�-�j74�:Ϯ���j��vS��lwv�KM!�2P�xpO>Xy���ϷS�ך�o�a؎x(�)Cf��<G�c6P�J��_T1�sM� �2d�n<�������|�Ρ�(s���@SqYR��~��v%�>A򪨇�2d��1aIb��U^k�uDi�n�\.m�59�ܿ*HĠ�h�7~��O�x�����c�9�R�M���5o��,�)0Ve�G���9����Np�x4��'X�E�,[�TG#\�w�
$Lk�08OI>«�[�����Ɋ1����H~��l����7�၌�k@Ϩ��C�ዠ���e���F[�r]R��܊�����}���\E�f�d�,��ClKV��]�� �W�X���PR�0%��!^o�Q�w]%i�����ĘľAzXoRJA�\Δ�f�����:~?�Y�#`VP�,8d}�b"� ���\���T��g�㠕�G����K+�ѹ4}+m�|^�K'fl��U�Q��~��ǲ�,"-K�����d4o=�S��}�A�RF���F�c~�hRQ(2�èw�,fk�c溘���YX!,zA�&f;�]B���TnM�_�Y�,�,��UY���H@�ugsq�e-�k-��4<E�i�g������G��7Gy*||vu"����?�.�	b�S�T�J ����<�1ݍ=:����K+�|z�:^�bv��������uֵ���&JΡ��j��G��e%vɫf�m�B�0�/%��y9ףr�:|��0/�Lp�򑟼B���G��z�eY��4�d�=vu��ק�O�T�cq���L����
�����w��_�CbZJn�1�0B>���/�[���!�>J�pn�����~R8��2���8���'���:8v�C���f1'
?�����]�������3qоh[����n�Gv��'��cdx��e��4�6��Q���E��<�~��	��߂�$O�󋩃?D)d�q���P��.�n��FH�w���Glb��#�rz��\�"@�~�r@�lAZT�� 2V��$�(�|O��>jg,4+M<I��	$QA],cU����{=��K5ۘ�<��7,�Zؾ).�׮��{��d�h
�P�@�6������>cJғ����8���I�r�7��r��8C�`�9��N䞤xa9�������" ��9�k�2C�0S�+y,psF�a���ț�*��T$�b|���g����yY��ZQüۭ�z����!i�?�fcz��'���m�7� `��e`!w��� N�}$�J�}"|WjW��>��ʍda��F]��dr�&�/�ٚ�_>܎��~!7i3��8k��sF�Lf�U�AX��Il.�{9� ^�i�4}$,=*�ު�ВTo��e�rK��KzLѤX=ۗ�:����ҿ4��L�w�����KA�"~�<_}	l��S�!5�$�;ߢM�$~ug��Md�\�G����K�����lm4O�Z�c��7ސ�ߨ��%o��J��Z�"ęt��lUѳx=VDÈ_0�]k-�^
Կ���z�~
w[�	r�W�t�m�h[�Ԏע�a��P�;�~.�6G1�ˡ����W]n����f�F����w�2'�}��g��<?SL�ww�����~��ܼ���a�8o~V��UmY�k^R[��`��2�jg9<qS˺�\��[�qk��*���}ٟ��0 �݅��t&[����Z�Rsթä?��½�5��x:Ɏ$o�� ��)��0j��JxjQdR�����sU�Vu��Mc�4�0�H���#uG8`���߳/��|a�F���`ԩ&P	G}��.��l�E�!|9��6���x-v�a��T��`�)JT��(Y�?����!���ɹg�t���N�I-������G���p;U��~�zi�~J7�V5�б�u�l3>��%;9դWt �!���r��zX�=�x�g�<�g��V�d�7�߱qh�/�V�YM��9����S�"$O��G6����@l�)�Y����)[q�哽�6�js���x"��/����mg��ټ5͹��Z�����D�N̔[�}�r���xr�rL��c�
	�;\����]��,f��4$2�Y��B=U��O�z s�E8:������<��aШ5��E��	�AF�*��ȁ�!�c��F�M�W���c�>�U�?�
>͌�ͮ���� t�ZYM{h�����oO�Vh�֨)�Ki�F��22���IY�}]}v���]ԤU��RL�޾����=�ZO=�^R���>�s^��>4!���I����m�n�)ᑤ����H�c�-x�X��s�)�;��[�QGA��Y�#rjJa
s5�nGvܶ���q�&_O ���ԇ��qH�Bт�	��hy�=�cP�e�W+��P��^U�,�	!��z���s�vy�6c�c��|��+�����J����<���J��sھX��c�fb��hNm3�W��5�C��<V�pP�x!-J��!n�jVtP�����;+|�����x�\�]� ��q�-X�� ^6[W-C�$�/�m?�,��j~�v���.�����m����Ds<��Uڟ�mMZHy$H���j����ʠX�Ϩ�p���0ð?|�Nt%1J�Xߜv,fGU����/�>@ 4��R�ey���Z����Q_S�[ڒVbӘz݆�B+[9��4~�XSZ�:���\��G1;l8���D�㴈�^��'��XFH��E�w�p�`��ږ��/A�^ڔ�'ՇϿ~������ �
q�}e#�l��OLNc���aֻ���Q���Qƕ&�-a���su����ʢp�R�2z�'�]���zViF
�4�� )6��0���.B���)�	�D�����Zp:a���=�)9��J�d��KNzm%o �?އ<A-�(<�r,����e���!���,�����	o[j�@Ɍ*J���l��%]F��� �	NbʤZ�j�ڜh�{�-̂�z�qɱ��x�e�,|�_�ro %�&N�rI��h������
����Y��&�a}!����:��`�R*L:p�j�ѥ��k���)�]��
w�a��Qu�a�7$t���W'ύ�� ӷ��[�t1�����s���C�B�!ց�i��ս��<_X�%�Xc�Kn�ҕ���h�$��x��p�]EW�G���@�5Ć�p��aaa#jtz\m�-������B�:,aj�Os�q�@�ӳO�̜�7�����epٛw��m�E��TU� �jS�AF�h��sX#q���tGh���Tc^�{=�ٻՁ;�=� (�uN#�����M#��t؊ދ�Cj�|NCY�׮���Bu,l�ޱ���<	A�v��/R��L��>�(�<���"�zIY�r�Y��@%� E"mc�&L]se��J���7���,���N��8�
�����YDL������h�n�uًҹj^���Y}-p�����~�9a��=j�ڞ�઻	��m�T���d �0�k1i����K��H����c��guxB{�q0
�\PFl5���P_��R�$��t�#��?u3����m�t�Fh��%0��O"=�b 0�#��?�|��k�
�wG��O�o-�7�7��������C�,�l�q��g�_xX��:z�������^��2��1�:�B�t�W��g��`[��tZ���)#���^7<(��`=�d�s����\�7���S�A &�� �2���7����ڨ��ꅽ�-��3�}�O=��Ŭ���p1���0��ș���r�]�I~V�؛���9�r�D�u�.o��hu���|�	Y�_տ ,E߃����-��XP��r�l̈�e�>���P�$fT�9�]86*��bt��[o�%dGAs�\�S0��`��@N,?�.���#ݮ��`��A�Yb�9̆���-u����5�[���
�.�d�R��g^7R��Ԡ��P�ΌcP75�˒<6�l5�� G��P/���f����#n�鿧��l�1E"�`�ZB����(���D�`(&�&�$ѷ��������d�N�1�߲/g0G�䭕��4�JZ�%�Z�$@��Q5ӂ��dK#���$���He�j�P��/,�C�q�C�p�G��ڼ��To��Wb��v9����b瘵BW�-�Y������	����[g�����8�BzgG(��$�+{B�*!4-�/4�-O���9�7^KƜ�
|������[���Q��e���X~�%u�8�g�D��<���ѓ"��o���1� yiA[����]�XF���S�ǣM���,�Ic���Z
7B����	Xk�B�KWR" 5=��
��8{ճ4�"���u����Y�������?A����J��ږ/+W����Ƃ�>��ߥ��<�,�%fO�Y�Ă�[�j=��ZS�(��	K�}L�y+�+�%!��A�����\�sb�n�*ò���i�H����"x��Ⴍ���׼�$?��sS��1}�Sv�(	C���M��h�E^��>F��,V�2�v�G� �~�3]YX�H�-�g�����>m��"m�@�oj��ݦC�[UA�E�@[�2Q'���)`1s�~"�`�p�2�ptк� 2�0��Џ^�&�*g�Up�� �wJc���ӗ�0��n������a�dk��[�0��:\��:���%��O�yTֻ�����8�[z���p?�6fB���_��5�����J�R��b�|��{�'��O	�=��� ;:�-���m$Y��72a�E���ݢ�ߘ��A��Y�r�"f���T����XT{�^�r!o>T�y?��in�]��fDu�S A4�~A�ۢ���wu�
�ʖ�,e�6t�i��'ψ��P��~��h(�37��R�]q�zm�͸I��|d��L;O{*�.}O�><����w��JEwbQ� <V��鷈xb�D!����/�?[`�&��^�a���ﺨ�f�D3�������:oj�G%:�|��$����]�zg�aN�͊��bi��j����R? c���vW$),x�t�*���{V�2�f*�:ߥ���E�be��"X���F�Z9�� �ȋ[���$X�m 2[�n�s��D�����B���X�$�ߍ�W�uss�����w���_�O�G^.:{�r������ĴP��D_a3Ypst~J���6�r�-�e_��7���@1ڢ�hT�4����J+!����wؿ�<ԧW����6D-�_��"H(��-�k���y�_��F}  򶉅r[:�EJ~����"���w#�F?r3�]8���/V`Y�`T��uZ�~"��ֈ��Q!q�+�8<Ps[(l�����-��^�a_�o=e;�P��=>!��R_.j>%W�owӟ��;m��`�7�>K�
��v  �X��uP[��j�Ȋ�[�N��($�`s�|W�6�Q0����tk�I!hf�D�@)i )pǙ|�#0��@�r�Dn��e~�z��YF��ym�Xk� �}���Y�6��E4�S����_-݉5oC� ��+����C�ˬ�ײ\��7@Q��Y��z��w�>%V�*����$��A���ő���G�wj����2#��{������=��^�4��Z��QEֽ���iXw�.�h��"�I�N��F�M�{�v�*�I�A"8���9�+�\�ɜ�Ze�G��i�+��T9Ĵ��g,9���:�)�W{#� ��=�ե��P �R֪!D^Q�H�����J\���[�`}@4'�Lz9� /�aH�����kQ���yO��z�=�:�j*a��fQTyF�mz<�