��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]���y��/'��L�?���T��_�I-�^��A�����l���s?��X���lUol�^��9�b1��,@h�ݎ��eԑ����һ -b��;��%R��04� ��1&:`�QQ�Gd������?�����V�Q�Z�������+���=Nw�.�vxoNSڭ����������ˆ�|��LU&���Se�wIE�׾'R}PR��,6�)�݂������z߭�|�]�Q�ҏn(,o��B�}�М�z\�NP88�m#<-Q�Z�K�Ŝ� �\�2����E"��Q�m]�;. �8���U-�l=F�Y��t	=_�l�b�ҩ�����d��Wbjhwܧ���-�09��8��ה5���]ӎ�D�9�*�k�-s$c"��1;�9��d]ɖn ���Z!���'[��`7��^g%&�I ���0e�捆�g����o�픸�𓜢�A��i����^�� =e>oӨ��ξ�.U�e��5�����zK�O�^�T��6�c�l�ڳ8�A���|$��-h���Lպ<���D��X���y;X~���e�JD�!�K��k�ٷ.�&Y�w�ƿTd!5�6�������55�:��.M4���-�q�i6�- �s5�������_��ۃ�9mB��؃iƒX�pZ�b�9�d�	<~���6�;����b�+s�
.�o����!����1���n�p[�c5����p�m���\�UK�W�C?Eg_��+.y�\�BÑb�Z�V]٤PS�>%�ʚh�����:0��6�}m��mNF�x�!#�Z�S# H�[,s3̒Gxu�䡮^�4,���Ｍ6�߃M�ĺ?�}
n,ç*T��J�Lz!;����L�T�ʹ�"�0Ѥ+�AM>�w%���,���t�J�귆����KK�o�|V���1݁��׎�(!��b��:�q�eR��^k�<���s���g�J��Fw��K$P`I��a�W��I��㕆Q�'1�81�ڪ�c��6y�7o�"���Jy6p+�e��z�_f�ä�ߣ�)�H�9Qj��u|HK���5J�w�<E������D�r<Q�nI���so�=ۼM�+FjZ�x�]U����
�J�h��+.՜9=�n3?�ҝ�©�#�BBV-*��&g<,>����K��]T��/��73�����i��=�W��kl�l��Q��*�H{�a,�`�ڛζ����tZqpe��+�d;a5}I�$��	0�?|�쎦\Kn�}���z�L�5)�P�i��&����SH*ګ��ר8�Ĩ9�����AdV@N���K�ҍ�7L��1����^�In8|_l��rlb:���&u{�YQA�}o��� ��a��P`V�(H��Sh&�����(a
�K�W8KJ��\�Qb���� �y�r��9z81�n����,������xc���|����JDdg�ō�ɻ��'Z/�a�R��r��!K����D�i�2)<F���Qvג�N0�ܕ8�)'�MU��y6���X�R0U/���o�.��~�+��qd+�����X���}LSj�2�?����X�V��qЁ˟LU��r`�QI�����'{���@��H���H��H�Y�8~���;wN�K|)p�{V���]���.ǘ_���55�_#4Jî u��wn��Q-��e��>f�-%�J1���X4��`[JΤ��{�mOǱ�Y�����@���K`�fአp{���A�{'I��_k�\0�|�\����p�*����[���(s�w�3�`��kΗ*qҷ��LG��ϹfTVAA�G���s���{��z��p*��$wQ[�9�F2 ��⭱V5�g�1�7Ha,�*E����Q{d�FK"�`����0;C�2d�8���m�%2T��*~�5����	�}�G��p��7�,��抐²?y�|� w����>c��	�8 �h���!���B��%,��(Ud
`�\�(3R5<V>��o���)ν�m-����x��//�2�P����AiD������P��n�b� _;:��=�� �p!���&ёb{+�2jl�Rl[IJ���c�$Iv �.~��z�N�3��Ļ�	����A��鶎gsu���C@�v��ylO�sV29.4�&��M3X��K&�H����;����:be,�x��i��2J�W�w�&dߦ�{��;'��:�n�Q5����gg��/y��?�h�K�Z�58�ҫ��^�N{r'�hy�ug���ZU'J��9�١sj�E�O�f�K��N����ͧ�����B�K�7��/� �/o3#���q�o��\��3M2r������9mWܟ�ڼ9����i�`�������+oD�:4o��*�t�>��DX�;�ҵD.\���B��@�N/���� �Z��A& ��\�If��Ls�}N�0�I�tG�3K��G�`Mƍ�1H���k�~B%�Օř�x<�c�wE^��eJ�$;j�%P  o�(���t+����D���i�@���w�j.��x~ͦ���.5��H7ī�񄕮 k��5z����Q�AX<�I���� �^���ߠ*n�b:��⎏�ɣk6��ܫb9��_wE������J0t�f��)��雅vM:_1_��Jf]ʜ|��Rnxy�Zu���R���{ʒ�uk�g�R�s�/>�t�2ц�j�:
J_�ZRpYi ������O�%�JZ-X�xk���ԭbjf�[�C]B����m,H�d���KT�y�Z��6�2����\���ԍ�䦣҆�,��5�v� ��i�p�U��Kbc|�Cʻl�0X#fm����Cǃ��݄�WsX����Z^�a6��ﵬ��Qu"b�!���
�p�1�?�ȥ����kḮ���A��M��t�U��I��k�7B����Ǡʯ �B��*�9�B��W@({b �%��N�B�.��\|<o���(��ܥ����ļ�v~�)��Z�6"Dd�!-O�>Wr\v���Q�ܨ?V���<ݶ�̬��d�h!%Lq1:��܉G��t{�<�~g���	Gʄ�GE��C�˨O+	x�E��Ui#A��ACsy��pu<̋ehh��:�W:wK�<u��m�Bu�>i�,�-w�t��Ʒ[��/��wS}�=wd��G��mэ�;0ɒ��Wx���,��?�'i�ZC�e�Pٻc��CrOǛw��
��5+�${C�k�G	%�uL�J��0��#V%�5�ɹssO���_�i����q�S/<Ӫ��~#\>Z�I�*���i[���&���`�zI:"�hҮ��g�߳C�T�1n�>^�{���q�N��!$��n�[fI#��eݶ�6
,�衮L�5�[D��u�n�Q)C]?gʼ�5Q`p�&��m�QB��t�W��(L��) ��4�E��L;�
��|��?a����!�me,�g+ \��ryR�J7k��1�ǀ˗�Gz	(��+)i��z����1���Éޒ֤�,�g�{���΂��} ���n�]�N��h�;D�AH�%=��bϸ�jR^��n��J�X���8,�����+x��i�PM�������[\>EYZb}2�5{"�����W��Rf�o�=s)��I�����1�hUp�[����r�y���ِ�.Y�����#�G
����x��iB��ff$ӟ�D_���1�p���RCX�S����������Qܗ�Q�U�W����ϱnϰP��HFS��ʀ$��J�WA���*�\�)t_�]n]�oHA"���h+�U,�i���!�S�O���/r���Ό:����rt�`���~&%�	�5��dt?q@l��R+սr����U����\�D�R��j��y��B�	��V�9q^�"?�@�����B������2��z~ ���* `�P�c��>!�D]�(g�������N%��������'A�B`-0[2�EzD��D��&E_��k���P�}(+������=5���:����v�a�i�kʔ���M��$�r��R0�bK��Ȯ˟L�1�$� =UG{�]
�b��|����Jv�r�}$ա��U�����龓�4s�ԏJ����Ck�;���r2v�"$Dpd/b�ȣ��j�>}7h�NDS �w���R=��d�&�%�!��M�S}�S��=*�����$B��S��7	:8�- m~�K=6@�*��"�$jE/tI�~�����r[�k}�"0���(M�Ф�� Qؘ�@���v8zz���vu�������z�W�9�>�׵,���C�x��kq1e�w�M+��l��Tq$�:9��;��>㜚
�E~����c�%��C�0�x�rE/�b3�6�
����bZ�L�`B��k�{$�F���B#�j
�Tgյ��9�̢��T@on¦1��t�Aٶ�={2���h�zg3�
�-GU���� ⦆�z=�o�U潬 S���O�J�!����� �Z^S.7Nj���� X
mG���r{�u����<GP��J�L�`���4������	�5��J����������EqЭT#��������9N�"�3l��e<p�FC�l5�&A	*<Â�u2��$��{�P���%�-�M�@��2��!�q�&L�ud����[)������r֛���0�@�8�5~ܱ� ����l��:� 1PS2�����Jx4R���A1�-��%��g.����#p�X|'2Ĕ�ׅ^WV�8��������M�w��u`�.��hay����l��GI��Y��8���ag��VI�Ji�Ok��Voa���`J���L視�`�;��
��5����Leo�!N�ςZ<g�F���g���Jk<n�_'zp��%�!��]AN4Uw�e��*׌U���4�>s���4�?�J���_\�����Ú�C��ߡ�&/����4�@�-Ňx8z���]�QQ��\�[��.�`R���&�nk�R{��R����QE�/�?|�w�k�y�9bJ��|&�#����s��=T���JЩ��.����6hy�+Jm�SD�vD;��"9I�\C��ۖK�_w��n덳ꍬ����c��J��E^����;���M�K�n|��܈��j�{Ǻ����&���-�pST�^H@9��s�\F�߄T�`���{"!9����t��|��i�_&=]0�p�dd�0�NVPkS���!	6�
\GS�=���Ԯ����J�+*�.M�p�E�l8+�g���pՓ#�cT�3�,��Pe��+�I����%y)�����9w�m��-p�f�������g@�.����0*�皕R*JC]ci���ǁ���-	�!��͈�b����~S������&�P̄di�90z`�� �BL�W+���[	�ȢFֵ[�wm(���s��z�
�Qn��NVhP������S`5F�d�\��I/\xp�S�_��`#U0�~#̦��~�t���&T��-]U8̐�nMD�r�F�c�EX�w��	��m��]�����I��8��G۶���9]T�6�2�!��x�f���[�²Of��ŤH�^N�������z�/*�m�f�<�&A�:Ł�Yɞ�@���iY��#7���n�AYM��N�ƪ����<.�{o��LM��lx<��ŃXv���C,��WK�paP�rM�8��6�9$�n��K&���m�r���.��0��x�b�*E���/�*J���}���\��:�җ�+	������^[��$#?H�/�>%���'O���߆��s���'�k�_�o���$S��fH�J�f���>>��Y�eB#B�͝AͱO���/
lX-%�qխ�J\��f2��]ϻ"˜����)D��cGd�1�cV���Ab��Z��9��Ag�J��F�"�N�1��xU+�Oe��m|����g���|��P�;|�wy�.����׳����4��(����d^yU�G�ڕ,����\BZ>��GuF"K��C��	��[3�ěh��늘����P�L^U��l��)b\�\D60@�&q�8���?-P��_iG6���a�A[gaU���2��*L[ylđ�76��1p���،�!gt⭢{g��������q!�yU����Bz*-��#SLH�w=�7���%!������۬}_���j�Z�3Bm�Cxʐ��)�ӆ�y��"�&�L��ɿ�x� ��u$V�������]�e/CY�%8&x��@�9?Yz_��XH�J �|��H��e�����4,�&]��I���㧀=Pu�Y�6թĕ�������c���Q�}��#�S��r���WI��2I+��37�M��N*� �m�������f�����K�4'�+���\�x��N�w���U�Q��Oԛ�fZ�6�od�ҙ�,��R7��ۺ�\�@ej���0'��t%q1�mb���R��B���`^�)܇"%E_��O�0���g�/�Û,)f ����k�ۉ���[H��0�E��fV��;��c��&��z;���#�]`�o�"=��A����Y��$�X
;���r��](��[��$.5, ��D��H��U:r�1���M^���K-�$�5�ݮ�9	��O!�P<�s�:
	P0۝\���s�D���3ONf�����Y]����!)R����tj�&n݁�,�O[��wVLZp��Oc��0CN��d�j�x^�:�mz"$���'^!1$-qq�q܎c^�KO�mT��BJ�����'#��4�q1~��gB��X�Es�$%*���+�U���<�m#�,��:�u]�]31�kw�s�?��q88F]Y�o�P������ݱ?��4$���蠳���u K����9�f��_�${�AI� E'3�T��8����eY���*��x+��N�ϟ���K-� i�i9ד�8�Kη�y�f�����#�d�"�,�:�����KXA��u�/��*���&�1�]�W^N.�����B���1L	j\�Z�j1���
��7q�47o��A)��n�>�#���te�u#.a�M�#��0��N{�v�b��ދi ^��m^�O<�Hn�t�T�\R�櫾��E6�?�z�����[�p9r!/���xT�����O��&�4���X�4�KgE���
��!L���1��k��ꆦ��!#X��+\�r�[`˕o��!��#�&9s���t�l�ԍ��j:FH���e)?f�����	|��3ֲ�?�6b���y����FE;��ְ��P)�����JQ���_�I!�ƣ��<#�Z��=n0�f��T:v"��ܯ�9���R�4���s�
Ё��ě��n��G=�����y����b�B�a�M׈ݷ�:�.g���6�C���A,��g&J͊��C����S�7�BH��r��!{r(��;Q�PY��Huub��y[�\2�,���r���1Ǯs��O�����Yx(�گ8���JL�A.̼��{Fd��+�bC�Ov�V����CMB�x��"-+ڜh�!m#�:DЮ�����������L�[w��i�5������V��¡/ָ��KK�\𥟭����7�1����ʄ�@���״r�LK:��Q)�A���,�F8���g��F{��O�����Mu��ΰ(� ����z&p��b�{<�K�ҕbE]�%7�`����0<�(��zް#�>�֠1�q:��<�����T�oiΕ��(��P7k*�"~���!��:��g6!7jD�x�q��q5�팷>BPy�D��L �c�JqeO�� 
ƌ�s}�K:��]��`�p��\�0�9�S�(�"�U�y	�����{�;.�hsF���9����ژJbr�}��\�}HI@���Wܮ�+#���q���\�So�R�ޠ'�1�G;�5�a�Rn���g����5�I��\EF0��":�A��WsJG�;��Қ-L�w�`>M�F�vȇY\yJCe��oe{�&��0�R5���:�1L�_�h�[���������#Si����,5��2m��@*U�sN$�
5_�љ(���:HF����4��G+���9BO��t�@[�5��^UZ��t� :=f��h~�+���Ѿ�M�t�l8G��s�.�̰����o��A�C8k� y˻��-Qh�S�\P#��2+�2N\;;j��X�T�Ҽ��D���v�S���Ѐ �R�'�/(2�m��e��O�٣���<'�Ng��i`�hC26��>��nn4�փ�ۣ˭�DT�v|�ewp��^�H��ϋɃC����θ5�&����>�
m�`a{=,<��5C��mck���b�L�@pg��|G;������T@�|Hca]8�C�@�����~��-����G���mo�.Q'@��^պ����f[�lV�.�4�@�G��6�i"�шRB ����L��^�@=���:�S��`8綳�MNS?��l����%�0�rF��M�����ݦ�d��4��X��C{�<g�3��ۯ��+C�y{۟&�g��)e��$���'b�p��ߐcrg?&y��w`[��[�SD�(�5;�@�����>Qv��L��Z�zv��IC��p�$�[��saS$�w��R�{�{X�Fm8��}�]�䥋��އ��8�>ކ��D�J���RO\y��К��*��c>�'��*3,nחpZ!Z�!�#���i*��� ��^�?7��O��q{�ְv�Sh�ڵ��b��Q�f�)�1�r;�-�B���/�ꬥ��'�Ym�ɋ;������}�VG���%Th���GD�IʲC�~?a|���A9o��H�u���ʵ.�0�̐u�;�K��s�Ck���U�ch�0���o5}�%��U���6z�B����h�����;����L���\0uמ������zqU��s"v��tH�L�~?�BM|�4-Rܐ"@����"�(���`�Di�5n��D�u��La�����W9�z�u�M��5��=�"�f��Xw��ɸ���%�����d#�����(\���	=���$!�#��^o]�G{ͫ�8�?y���M����g����G�gg4p#h�d� �O����i7Y��	�I�L����5bU�FRC�K��E641�	�E�,������p�:�
�����_�p�z��`��bvi�Ncu���G���9l�2!zT��a��EHA�\p�T�5�bzu?�S����N9{������r�.����l������	C%Aw�mQ���7#�� p���e#^i⻾���H�������s�
<�պ�ir��^=�n:��-��J+B���3\幘�y_�5�k�OU�)�8����ǰ9�F��Y*uN�q����Iw0^4E��1դݠIRi�F����6m��j-f�Ko�U�ln���WǷT��f^�93���T���:�Y&(��u��<���_�@ԓ�#�~��Rn���W�9����[b�w\���9Mx`�hB���Tph�Ɉ�����T'��'��<�[��hڻ_�<�H�����DI��.:�0zsԃ+�X�z��&�jY(������/���&��ǁT��� ���z���y�P�l�=G���-�r�FrĪ�Ucb=��tEu�lH��7���M&@ڲ�YL|�ѢDb��D��0��N�8Vnx��Ǿ��~:Q�@��|@�%�7So�4�b��s���J�E����?^�q4�Z�>\��k�ʜ��b
��&R}� ���(��u����E{���3����çUε<�����!��yN�JʉZ��jj~.̚���v�
z�а(��Ǎ�/��,�9�M�A�kS�Ș���`(���T|��')_��X���J��X�4�h���;���|,V��~K�ސ5~����Ȕ�� ��NO�z�j�ޘ�<B���u�=�R��K�Y�4�����B��B�����>diە����N��YXw�e�����]�N�?�zm��S9ȑ0d=a��I/��
�����̼�o��w�|��F݇���B���D{���O���)H�ĥ,x��A�@3	u����o	V��`��=*9 �3��Q�Z�f�v�Բ^������������M������阖�Ȑ��VL���OLQ��5�Q�� ���s�qư���2+Cp�a�Ug��4fBj�c���}e�3Z��x��fD���|Z��?�*�:y	�B��?�x8��I�
S�X/th��l���:O�
P+j,� ���x�E�c7����e���|VG\��r4yx�t�!v�Sj	�X��'(&��1�դ�F{~�w����{x�,]�LH;��L"�q��[���f�~��{<�9�fE1�&��!\�7�\�3��&\�IcP؝�t��%�MV���vpR��Ֆs��Ц`�y�+�ײS��$�������J6�ϝ7 ��%J��a�V!~z9���F���BՓO�s.%��n�PfQq?U�<|~�_$�����dyMC����יI&�f�C~ʿ�$A���z�4����M��0{���U�S�"&�D�?��i��]��~/rH���||�`O�#)��Ł����ٳ�5�ЃD(�e�}_���M�t�5��:���Q������;�ݲ]2�>���w�"G��VY���I@3�ػۨ�c�3xj������3����h<,��n3*||(��,7c�'?y˹���U�N����b�!X$�kF��\�:��
7��/|KC"��=y�,�<X�p�<̕��B��c��JU-(�R�r�A�����4�y7���=QK����|H�#�d��.�P�U��0�BU��e�D:6�#q��R�����O2��F8�-UP_�0��~��0��>qF��7I��D������|p4c&���
o1��s��������.S�I��6~+W�Փ�s��2o�����16ޝ!~�Q��S�K��`���5F��xVbR�j~a�H�_���mkX�^EuÕE*B�.�S:��Y�(͞���P��l,ǰ�U5gH6������Nq33j��[�m��Ԅ�s8�BRV��P�}IO崗Ixe�\'W��!��D�ۧI��V{gM��,�p�}�f�+R��C����m�]���m��߮��48�T^�y�a�T�wz���opv�`��f=yUH��&��<6vF���eb���܊�_�E+6����Z3>��L�{Qp���4-!�[���2���O4R/q�u?���"R����4�Wd���
�O�ku�h����'��.ҳ 
H�����	�T�<�*�dI�x?Vw/O#hZ�毰��v���擣���Om����/���_縁��@B5�{[�vٗ|��&F_�Z� QJe��_�Z��t.�����J��Q�/�.�m/����)�:�W�[�	�GO��Wo_} �Q{⓰'Q���sE� �N)�&g��P�
Jq�Ik�R*�PҏB?S�zo��yԔ�$�ޢ�T�/��?�☦��f`Gk����׬�l���g���/�zO�F�)���������� DO�T��	q��I�.�0����.�$E�*��C�`D{Z���q���3�	]k�R�"T��\l��~ 潐���3i�D��Oݜ2���p�^u����n�	��h���	�;��}ò�K g�OC��k�X��ӵf`e}�P�l���E|�=�Q�B�"�H���>ƌ�o��#�_��(^6ٞj��ו��
9s?*S;8�kD*���_�Zv�@-b(���(��
�����yi[Go�	�t��3X�Cn�h�5��P���}���A�Ҡ�A�z�o�s�ﵙ����x�}'y�ʋb=�~���"߫��x�t<}������QAd'����e�m@vf��^����7yN��_��]^uMo�g�2�TI�����T�<�I�<Si�н=�'�J�	�"����:
o��ڝ���5D��aS�dﱮ�Kf<��M�^�J�
�A*��b(墽�<�-%:��j/�0M�8�U�`ǔ��:�y>&s�T�>C�-｣����.�Cǎ���z']��ރ)b-dE�R�j�(Vԅv�w�g�씋6����6hZ�R$`���d�m����h��/h�~�Q&�Η� T9M5ҙ��O#*`�I�e�6��Pm����G����Ufz��+���V ���R�_hQ�8�$Ja�j�*���n��CM�	�ڇ� �H8j?ɆЅ�ӂ[��NrԼU�z�3.e&}I�
-,[;��v)��)���O�y/�7z��Lf���h���Eټ�h�+~���4;&]v?�ɍ�����L���7PI%O��Y�B���o	���P�eST��0�c������x��"�]����Eĝ�����t�c"���L�_^N�f&��?{{����g�����`��W9nK��}��K�h+v�������7�����|�O��`��yCͪ�R�3W�x��X6�r|7�j��3K��8'�]Q��TlM� ,&#�v�A�p@��=.�>S�N\�7L �"�f���{X��F�N�2���]O�D�-2f������$1�+F*��Ơ}o�:Hh��(�DG\`0�4ܦ<Fa��Þ��e��0�>P74C�ڦ
���"�$u���JX�\�J#���Ѿ�0_0�MD��.w���;�B��2�i`���4i�:��H�Ҡ:�4후3�YP
��_�]��KWp�E�+K ��`n�\�;��-(`�y�+�Bg>mo�;�����OW��@Oc14�ŕ<vJ���R�N`��W�,�4�!-�y�A�*;������sU�&Ԙ-g=�eN7H���ăȣ�1?_dp��Y��I�$��cj(���q�>���U��0 �#�9�NLd�ȿ�:��ξ�ALˈ��A1�p+�9�05y~1��:��X`�~�0�
�Jm�2�)�@��z#������b�j�y�F�9ASx_n��XɃ�3y�	��ߓ/�M��X�e3���8�p��9a3�"޹<ᕧx��������a�H�� v�r!�b_���i�[ �Y&E���=C�?�U�۸�i����C!0v0yI����苫����7��Vh `pƹYb?�E\P8�S��\3o#�4�����IV��6}�Ҟ_ ��i�).n`H{�3h�p�\�wA~�t��M�2.J���K�f7'����a����Bf�B��M4�It;��%l�8�7��n�Ө��E��֟���B�Q�cO�D�d���`�S]��s_mӓ��e��T��<�L�� s���3o���y��H�em���W��%�,>����~M�Yʺ��Ӡ<K^�HZ�_$��ǈ�������{�;�Ԉ������Yh�#�h�r�o�B1S���T[�ek�͟�k񉕘�"����dq�n?j�B�ZK�T"��T��mV��p�Lݵߕo���<S�5�n�f�a�y{1�߸��w�)�*x;�N��ʻ���GWss$*���KuJ+������>��J���*uB=S�bEǄ����09On.S+GKn�p��U�_�ύ7�wi����ыA*|£�6�yx���E���\���B@H�8M�݇dJ�u$.Y6 �ŗZ"teϥ�ǸN?Z���*��wPg���w�^�!/i��q_���wê^~Jy?
���2�V
���� 	��k[�)/S͂)������v[VO�y�<�[��ڏ�h����{����$��oY ������+�k�o��Pm�9�{��툯��Bx���^$����(\u?c*׻���S��<�����<g��Q�S����s�6p��a�6�Z?Q��x�ŕ9~�:��� �s%X2`K�3|��g�/l{��ZQi��mXR�ë�7���Yك�#�JA�*�z��<���Ky��'
��a�Z�iGA���jcOR{��K�L+c!�`��7�>E�3�!_�����m���6ղDj:�
��W��;���4�G��~�|Ȇ^i��W Slm껮�m�vX�#csӶ��<~G����d�L��}Q��r~9����j$x��	YVz�Q6IZXHH�*p'�y7Q�]�ݤ�s�+��@4Ba[ze�EQ.뢃H�uÛ�1Y�I*����C�*��ǽ����h�]Ɋ\]�7t��G@ꐛ��v�|x���]�&{������X8ߩ����(Y�s� ���M��ڏc$�/l�S�ݡ��\������*,�m(7���[�<uڨ�KF��uL�W��~b�)��`��s$� Q#$�c�t����h>�$�?���X �S��}��E�%�nQDg����\ e]�`��}6K�?�ZRk�<��»���_Ӟ�
��\*ᵢ����kS~<z�/���F��~����欠���MG�|XS?gKC���.t�o��c��Lgt$-�>�bf��

gz�����!ۭM�:��KQ/�����js�!!ꦭ���^"��)楺��\�W�&b�\F�<i��}�WE��ɥ�	D+�p4Ř��[� �T%,Aq75a|S��ө�5�ѡ�w}:4�
�*3ρ�]���L�c�e�(��E���*sM�@؃1��$�Kج�rl@o���`gN�[��u�O&��M����<24H,(1(@�OlOLAc'� D��w���5YY��b���&�7{�}OC���� �ԹF���Jgi�H#�>��_�~ឰC�Ŕ���3�&c�tOl��ѠZ�+�%�B?���~����-Z�)�4��A\�Y��%��>���'K�=����������p
7(~�<�M�`X�ל��v[�g�;B
�7�!w��w�2���L�f6�N�w��ߧ��&Ձ�=�2=�'Ƴ����E����J^A��F��/����n[/��ڱyd�ʖ��=/|������8*�3�]R�Q�B �lώ)�o��5����ex����t��!#Y���i��g��q��=�a�DY�	5���Y�9�b�)D��R�h��=�����ؿ\�A>	����=;�SPi�����4]�T'_'�2��9�#!$��5�n����M8�����3�EY�{8��Z%Oϟ�m>�{3��͵� &�{K��$8�%4s-�Y���X��q�@d��:<hvb1�ܖl�Mzp�RO̬�N]t�����JK��
8���E������n���_0HNOp0,j_�����/�0��]�C&̅d����Jb��.���7]*l
@w)U�=!;ߓb_e�1C��5}IE���G�5)�Y/fE°�7�5?e���:�S,����8��D1Y��lO;���V�pzi�����l|�5;r�\�RTW��7��:5��h�e;ct U�/QU1��Q>�D�7oD-#�<.���������{�2޿�&�p�XD�&�>'�����}Wg�I9��,q~\a���K$��5�R,b� `I�v"rG�ϗ]���E>� ���*�3�E��ܿIQ���8ֺ�Y����mG#e�������D?2���\B�����j|�z�XM"�+�(�#v�k�㘵hn�zB9�}�s���I�=
�Ag�����l+�:9:K6!���l�PʬJjX"���bP8��LQ���d�;?�
��N����*�>Vi$I-�4H�����'h��7%�V���F��\���S��O�f{������:�"fH��>�Hl+��?��b�joDT�O�wyK'���4�f��D���Gx^dk�x�1���"��]�x=�Δ�m�d҉V�s��ղ�P��z�hQ1w�6��G7e9��_���{%^��FZ՗�8����]��oݟ�C��MǦlaP�rUpYpu�TS&��BDĝ������w_\�h�H��� &��h�����k(Xk2 �C�s2\Q�!�i���'�}T����%9�(aTG�s���)��p����m��gY�_J3\��A��GW2�Z���J��uQ= x�5�U�}������sӟ��%�����x��O�"$|}t��œ3֙�A*����%Yi���a�JkYU?>H�D�ݢ�0�t�oXD������4�٠v�_��6�ε��C�T����|�i°l�$;ݸ@�X(Q�+�0;���C����^��`��'`�?W$$fe��{��_,QO�e�	����P�b�2�|��(�kvh��<N��������GAw���~l8\���S	hC$WS���$�NU�KI�1�ԗn�
e�sN�޳�r��z]��1e����l���!��K�5���gkx��;�fHdZ�W<B���z�b{U�P�^N�~
��*�p���C*��+L@%&c�����`B;����ގ0!��ɏ�@M��hu�ꀆQ�'�X���E]������D���e��_�wp�3���zZ]�P����ױan�*��d:
����'Lx�N�j汔N���E���ڌ~q0£���͒�c�7�r�N��Ca���w�<.�=w�ה�$^Y���)�q␲-�	hV�( ���=�U3U>��`mzM����!�E=���M��#�BK}�;t�5zn1�l,v���l��ҙ ��k%�`�/՚_�u�S�JU������A(J@��|%��=}�Cwd	��1���dY��J�J�32D��f�(�!����T��o7F�O�nV���u#_s����``	�5'+��ng�A���܀�vz �Ysg{���l�j�r��G����nAo�Y� G�i���q�|��y6��NX�R0auh��S��Aوz�E�riɸ�4�IL������y�Plh]Ď�1����TŽ�e���ȹ�Փ����X�佲]w%����������p�l�4�)�]���Z�ʁ��b��l�m7����QR{�F6[���㦝`�L!AM7+4>���{�&�w���gף;�����d.;����i�Dn*��`�F�r�QKHp�@�`��%����rW��v�&h�b��@�]��1�w�
�s^�����ר�7�#�H@�}DY�@�C)���!��4d��JW��S���o E��sو��T_=N��s��,#��b��h�k'
��2��8������{����Z
�G�Fg�D�|��x���|���ĳ����-ܩ�p|�i�W���s�������͵�ı�#+B\%�w���T����D��������YZm8��];-)��%D��e���2��k�{�����NA��
����2�V]���>E
r��9�8)��o�W�
��|��j=֙v��+��ޟ���y��g<�Vq��R8�zJ�;_�z���������@�B�#Zh�AS���e�J/U�$�`ZxMd~ك��^E �BPTAȩ�씡��I%`�wN�O�`8�U"�����4?���=�l���Tq�.Gs^#ا�X�g��ct?42Lߍ������N�ˋ��Cbx�p��xo^g�6���걕p(ZJ�3&ӟA�Pj"�6�$0���+aW�y������xڎ���u�˵����t����1��8������� 2��1�y]�{�gF(���]���w��s�g#
ӻ@�
-Ą������J6�'����	���`s��&1�SG]�%Ubc��c�%*�:+�tOo+��SM��}�[�3[7��O㴐�F�~��&I:v�y����3�7�-��[�5ɮ�@!wt���G0ݕ�ɡ-dBpu�Do�C]�l�st)�;��hbVGs$rp�+�^�.��%�-O[*�aC���3�zǓ���GT��y���*�b;��lOM��s��j�{ �GGZ�QfW��Ď�N�T�Z�1�;��h�z�<�Y΂�������H����D�F�ډ��h��]tH/��6���}��}�TWB$[�fMD�X`��N�Y�#?�w�7D�]��f�	7c݀���~��Qf<��7�>҃"'� K{ES�@<�|��دa���+7�ĢG
v��N�C�̃'e��/����yQ��@OW���.���L���#�̄q
l��� #{<V�F���/v'��bh+��>Q���3�����
�Y������e�������@�!r�zw��rc-Wf1ȣ�dEd���о��p܃ɋ�t�Y�׿�>u��Ĵ\a�q�����-ќP�E�H�A*{<��b� �BMX4��j�X�ޡ�~�Jɵ��/�� n��*G�	�,w=������"J��Զ��Ryù0��߀(K����_��xj�����Y@�7�h�~���=�"<+��h��J�_I�<�
E'b�DXF��D,"$�(�I�z3�=��E2�J�-q,� `�2NGb���:��*�7·���0��v�j�s��C�l��׿*�������*�:���ǭ(����Jsl|�)>J�d0O�[��mS�x"�߬�*i�#����Lj{�~`�b���R�k�C�`  j���0�);٢R=w�yZꧤ���J���#.LmiSOZBU�5��z��� �,$gm�9����l\�����^񫙡}�M5��v�[�e���Is���r��b?Ծ�WfXg�X�EB2"�JII��Q������B�)f1`�C���߅R�y ��U
X/]�����H<F���+�o����`R0v.��?��	mXױ�|��x��q&^����
H��D��!�*�j����ݢK$psΖ6�Y
�ѱ&
�r<I�����=K׶���qQ���I�6�Ԣ�20C�Z�%��Rvk���_��0� �0��O#}��wU�O%�B5o)ISyv��L,�c���;G|ո����#RZ�f
K���+$���f_,bZ��З/a�񣺮��'��`��#MEJ���fa���]);I���6@B(=�WG�A��S�y~ծ��tc�����&����*+�M#��k�h�<�t����V�Q������SJ�{de��{�(�o��k���	���}�X�攞�׏nNʽP���?���^�E�p>z��p��IC�f��jU�zM�YX簳� ��~Jon�:�I��j,����Xŉr��\��� y_�sf�,r=�u�<�}��;n�������*ݿ;d3��P�.���Q.�x��~����ı7G�Q�מj	���[�]_��b���h�N��=/���C7h��YѤFw'nHSc�uѺ�n�vi��9Ҙ:m ���1��hg���l��`�?[>7���.k�_Q^�V��D�&c�� w�A�唷؜ߊ&2Խ�l��1����L��;2	�)|~2�4O�2�D��+�Z�>ub���-��l�|��W����!9��%��w�Yy(gV�SX|턺�Ʒ>���Y1�y���P�6Na���5B rω�3�w&I����g�/Q��.��c|ԑ4a$Ɉ����)�"W�Z�>��R{_Jx&�P|mK�ŞcX��r��Z�V����&!�}FT�_������C��:�)������R��6�c�u����JdU��'oco�Y���`tZl�w��5&�=8��Ov̵?�iX5+�����5��w��Er! <h�P���zg�w�']]�7ѓ8ǿ�`�Ow����?�鮽 ���;�R�y��
�M]vw&����G�5��
�DƠMb��O�� �m����4��(�۝�Au��*�)����uQ�!���"���Q|�,
m;lQ8#3]= ��B�U��}~e�w0��ͬ�
8��B�Z
������V�-��#��:���Q](Rz�7�]x~#�v4�����0B-J�.�s Q�wN���d��^�O�v�w���$�ŖbJ�T�Q��G�.�� �_��=Q�;}Cј/��*�������s���jjm+�Dg9)(w��-edmԩ��O���U�x,"��I Թk��m�����<��SJ�����Ң��TE8�b|�����tʥWz9Qp_�0�L1ԗu�VZ��+��Ȟ���8,��ޔ�O� U�Y�cך��g�0+|�~��zშд��S�Q��� |1�R^���V�'���+u-Hp�kE�m��.��	�����mc�����r���]Du$+X��7/��"�U��ª�C��^Zm�fq����XH剳1Ձ!`�f �&��!�v�V�?W�-N�� �,��Әy<��1]a�"������!��%�1�ǘ��G8�SUrm������7AC���^�UAPƵ�KQ-*7���S?n.��]Q��۫b����CCl��%��T�Z��|ޣ��I1�B^80f:��"�dס���*���vщT�o#t��ЎЭB���UR�e���A7s}�cN�uaK䧷R��p��{{��TR@� �	v��J�"o�xe���&��RE����W�}e&%oTs��g� }>�WF@A_v����{�霌��Yan3CԔ�ᇝ���E��2��!�Lߒ���\�6G�䱒������=&%e�/���'�Ů��-'a�lU�Pp>k�?��������
H�<�� +ڥ�H��~UL����8�£�����y������L����]Z5������Ť��QL�����2~��r9�	7�`?.�콐<(�m�C �BD%����ҏT�g$5'�E89�j.��s��$d�b�%o��Z��~�]�zJ��=��m������𱉜�E��דj�/�Xj������`��V@��|����EB@Z�o3_z��ya8y�&hlL��}+���D8�7�˺���>��1k�tD��L�<Oe�p�����9��՚V"�;�m���ަ��5]Tg(�G��r�7f
*a� H,D�Y��-lQ)*�C]SAk��e�ÿ��֦�r�.�[�ť-D'�>/Ur��H������n��\��8͸q	�q	6��yb�>�!ޮ�#�h'VBs@+���D��`�.�e�~��4@��B��۽O��'&6�?��N��.#���dR�N1;�x�f��pQs선L@�h[�+�0�;9�����N4G���g��ߦ�!?pvV�4�PߠRE�O�:4Ū��[��'��Ql���!аQ@�<0c���K+ N;���9Z$%�J�ڗޑ��g�FQ|�&낤�HXb�����{k�Ԯ���`,�3��#>�м�2wy�8�[��R���|`+M̀��w(ܝڸ���B���~:0�1�B��vr2	� u�'\�3����6�F��������������<T��a�7ti�1	�w�K9�$�0\�˘��dX ���a�l8]9��vq�Vm�o�j#:��9�r���?<b�k�����^Q��3��K�$����j	T���y�ʟ��To@x%��r�����Ҽk��A�f��	���"۫��<�&5�� �w����Bqp�C��{����(N�%�z�B�XB��>||�`"PߡܷeQ)A�������0a�^��ϊ5�������O��+��hW3���x!�"6�/�)V�OA��z)��R=��vPq52�ň��f�.�����,Z�T�̹�A��� ;���3&8�i�I�[Ê
�?�p��Ss�q.$c�Ꮔl*�#�sG۴� U��0��
=/V�!���L�p\�P�h����4���q����/��$"6��
�S��!LŤ|[gf2)iC+�� Q�U"�$�1'�
~<�@@��ڱ�e�m�@�l2���� '
�{���n�v>�g/�ò@\�E�V�&�fj�p��\�� ��_a����I��#������w$=�խno�!m����L�D�������QN�Gf�bm�T$���z����w�80jD����8�6�Œ�����f`~��էIA{r���Ģ����b��(H�H��U��h�8`�}�Cl�Ge�覆�p*P��:�C��`�]霅�TD�����R�8#�  A����������ۢ�aD�5�Ũ��� ���(RV�]����/�F��XV1�v�y{s���o2ѫ����ٟ�P�k�����b�&ǡ��4v�A}�;Y���R����P�)���4[�.��¹����.S��_Ub��e<�5�e��K�Mַ�Yb��.���K,ZKYte��tW9���է�]��Hl/��B�=�h*꨼G�g $ۂl��4N�1L��������{X���"	�99=sE��:�A�M>�;=\��HkZ�L��wMʁ4�:��
l�����3�����,��z��eMHJb�d,���
�կ՘'�+��.�bϸ��8�E���O���e�M�+���l�s���G������u�������7�N�Z�@��O!�-�k
S!�=P{���00+��A]�+A$�D��y�m�c"T�Sj�?��+x�왿��Mm�Ϋ$��9��˵�4���N��S��͈��Z�A���H��{)aaB{@��jy$�|o�hg���b��A�k������r��O}�謲)1���g ג����z�Za����T�s���M�����Xr��C�+��/�'S%F�?h���u��m�\>�x��xy��gp�l��u|���Im��*߈���GtC�d���*��ۚ �9�aXd ����`,щ����a�9��q��yHԛ�����gY�H_oN�;�|�Iq�mo�(W�#ź���;��r�m�X�E�'h����4Ce\���^hr,�E�0���3u�`-��W}wW�ߚ�;��nd���Y���!S
�k-.��qJE��A�lC�"�ܐ�^�<�޾J�Qe	�w�	�\�N��j��K.{�����u�ށ^����艥3�*Ш�q5
�������R��%}�ܹ��6���-�?��v�K����Y]$�k�l�#�ag���u4Q9k�vk��xڛ�{7����tO���H@���^T��g�����l+VK(�Sǝ�$�c��ޝ���P�v�e:@[�bay��j��1���#J��v����X4�y �;�@�FA񄃙���/A�]�Ե)��V����ɿ�#QB�*eR��Bh�'�y Q�4�0����N/{���}q��
+�%��{�'(�>^6\��&��$�K`�$(���A�9+���L��96�y�O�4nAef0?�#Ld��A�C��C���/D0��֖��])�&�?�h� �1U0�a�z�ߛ)�2��7�9���И�s���s��jp�
�CrE���i��b(��DH,+��M$����7��|X��g,�HB�|���}��e%r���٤DTCs��nC0 *��C̼&�#K?θ���2�d6x����S8��"]\���w��ݤ4	�'t��.�nd���漆�Ql����6v�j-�w�sx�)4��a�	rOw���c��n:�'*���xjfZ�x��du�k-.v�ܣRG_��Ag�g�`vrO��$|H�nR:`������Wo+���[�}9����(<$%�q	f �J��K��X�Û��V�iK���Ј��^�)R:EC�z{G��zo�n���/����H�OA6�����S�8�� ʶ��c��Y��{�bb��ص����s�~�җ�ɍ<<���� �|XM���+{Q�����h��pji�4 ��F��qLU����Q0�p�ݤ-F�0���{zR���P��c�5t�;�~��lt�޹`u��9܎���V��0�;D� M�D����0gP�Q6��S�~9��J��aE]r΃^Ѝ_X�$m�_PI�'��S����^�L�޼�������f�3��SZ��`d����'J�*ZPӧe���>����F=��ZEi���$�N��v���py��%���a��VF�Ї���?�_��3/<�I
���T�h�S�J�����k?!�Z f�i�l�C��п�P`5�wKO�2<1�;<��G�%�M�`��=�4d�B��sH0��<�V�#��N����$�3�71)� �ǳ7��H��-I�)q�s�X��d��.Pc������(s�)�́���ǲX[�8KV���Ƌ,�P0�Xs��`��i핀Hm�ӓ��1�K�eDAt��9-pu=���fpj�	��F�!\�T���DAT°I��1���N^�"Y�	2���I�;�|l�E1ݝ��T��?�n�t���q�`%�����,
��*ˎqH�k7�T���M��bJ�w��S~�τ�����V%P4��HΆGb�_��b���V���!I��ڢ��	-Ʊ8����  ���J{��Nּ��I˶��OSUW�P���iR����׵�̙��ࠅ	�˭ӿK7��L�v�=S�k�$�&)�
��=yb�I7�9z���ȝ;��i1�R��,GZ�����O���mP�OĊ|��{�dQ����NC^m�Jl`�ʓ2��W�?�M#6n�=� r��·�tړ��{2���n�hA�V�0��E�}�@M��*{��$Y{�(�LPѲ�˵I0{URp�ҹ矷�M�������\5i*b�q���G���+���R	���5�E��h��ifY�$��5�=�l���W���A\,���`�L�f�L��ʬ��#�R^^��aj��:��Q���y&-sH�v�D��2�Ӌ0��Q\;{y&Ҩ8:;&#t���6d1i��e�+rxLo�?D��Vo#����0�Y�rr����$���̩�|�zq��B����fOsT���ZȉȱH?ӿb�k��nF�x�!i�"!��LSd���G~Io\���Vl��ү����b��9�M�l`�yAL�����uO~�`�4}	?I���;�| ʀ���~TfJ����	�����Ct�����F���Ox,ȸ1a��͡��n�0{U�o���PR��B7�Q#�.�E="��uz�.rS��ga�<S�@"kdT�B�6�kX��weW����1r��a��s"(:<���h�l������㰿�uMI�	���Yj-Q���p~g7�X~�4�\���F�+����Ɯzf�&2yR<���e�*۞�9U&�����7�o���B[Lk���(�G����dp$>$�@	̏}���Kކ�F5���_ƇըB���JD�8��2W��c�uW�
�=�e3��n���S���Z	:��\���v�<	���bԖl���䇌f�������{��gVs�.�|y%�+�V�4!�	QZmԵ�<��|:3.����X7��x�a�&p�7����	7�	�y��)��d�F�\.�?��u�֯�[�K^3�;�Tp5J8��ՙ}���r������Q� �,~ ���e�/Rz���$8�#�"��+�&��m͊�ɰuW���@�Sj�u$8���,H[0$;D5��?�������0�Gz�ye�{~e�ή�g[�1�����"��I����\�����V@V��	-9vAB����H|=|Lx!ܩE`}�fQ�й���/���\p�zn����b�)}�"������R#��j$�ޛD�;��o���-��75�\ƚ2��u��JDk����}������S�c����RcDH����;�-���t.�K,H���~�Z���_Zo7�8�X��T`�gyK�D�O~G�"�b��V��U���uh|j���f�"�V��y���m��E%����l#LhK�)�!R����AkQd�(��E�l咓/���4t�:F5�A�逖?���:��Tٯ�+\)K�/}'"1G$C��$c���?bc��ԙ�|�WQ��w����v��Q=�� ^L�ֲk���'3� ��1۠�ʭ}S�TBIY�$����|x[�}���[ð���P0�Xu����`5�n�'�@?v��x&]����6���_��F��4��H�.��e7o���|����3l\7��n��Q�)7b\${�t�$��r�3=|8m�o����Z6�VΌ�� �0���=�
��U�F�|�U>�
� K�H�H���A�,�kJ]�c۠��E�)�MN �m�_k��x�C�G(r�|G���c#����[�31��5СfWc;:)@6�!<%y���H���V���w;������Y�g��pc�����ܚ-�p��\'�_C�ɋ��4|��dUg;Q�h2�J�	��0>�<��ğ;,�yH�;����4��p w|�O��;�B_��D���~����EwdO��\��#]��f1op�����}����p8���*ϰS")�8�G��ɒ��o�m�;��n�.���A��Z+�|�c��G�6��@?e�b�e+���Up*�6���(�R/{�Ř�ij���d���0�&��A���sD��̜�=�m��F}sy�&�o���UlXlݢ�%+!
Q<�^�<5�x���+�$N��?j�jX�0ׂ�j�a�y��!=�!Ȣք�]c�	���(nV��]�����}gr1{�D'Ю�%��$:��P�V�7�S�M� ��ܾ"U�`�Y�V �c v��2A8�=K^� I�M����~gnc����e/ߧ��%����O��M��Z��!��f�Q{���P+܀�%�۴n>�������O�y!�@&�T(�z�Nm51�l�d0\863��ș�O�zKTǡ���EG����қM����S�z޸~GPQ;���Li d'g�5LV'D3�L�X�E��GJ��;��]Ôf��Tz߯+��ѕOC���R���i�-I����-�'t~�!
L9-.wC)np��D�2t���BG����(V#-X������sXn�{�ϡ�.7n������v��*˕��oh��fGG@��-��8)�^�UfXP�$%�3�h0�5���mj��.�`�/��~�dTp�6��i�Z��h���M\�lS-�+ ��
�O}5m�����T-GK;��>��{n�� ��2S5�n�Ym�M2TIx�h��ԃ�-"}vU�3�<fovYO��̖w�3�;CX0�xo1Z���፳�)�#�J�@#�����Od�95��П�n�Xz	�1�U=9}_BA�e�?���zIu�A��/��������0��PgW��7��bĤnrG��G� ��:�M[�M�	�@�M��Z/e]�*|���m�v�~�_��sH�z:XcS��+_:nA���1!6�4�5<�ݾ1i�_�կ)�.0J=��}Պ��r�Lӊh�8f Yd��j��hYHE^ê�k�L������3���,L��Oj<L��� q�kUY��j|���-�v}� ��,j�<S�܌Q���0Mi��${6�U%)���K��4�}1�(��F�w��fk�^���kG���2��uP�wɋ���Z�¯�K�?�P3��Ie@ ٯp�QÝ֞]T���j�g�]�d���<jð�L''��N�ef�݊b�87��[�Z��S��J��`
��Re%Z�n�U*ώ2܃1�7�U�z�� "=}��KגL�����΄�t|�� F��t��V�B��G����^w'Ya�s��ٚ�S8-����JS;aԝRVJ�B��J\M������?K@8��:�+�ThxR,�k����}|{��]�5������e3�൓�#o<,�{������(�+	���|q��D؀�a�.�s�^��6N� 8�7b9�@��q�b���0t�m��7��G��.8�K��ߚ����arco����w0�"�I�r��D���/���IlD ���
)�, �w|��FF�N@^���S��u�Y^񷲄Ϲ,��(�49��,���~�k���&��|���(����L�n�ɯ��Cz��c�S�?w6�$�:��tx5K0�J�O�.g�FS���"=�:g�.�Dz\KΫ�K����Hޛ��}0����j��@b����a���b(�#T������D�������o�Z=;���^I�u.埐���������HU�/��S����CǨ,�|x`�=�Ў��{�l�\�QP3��lF����L���2+�R�V!���=��2d��=e�˴���O;ƘǸ����w�1�����P1�A}��G%�ۉBe�Ny����E��3�me��cݽq|���Z�s#����6�b�O�^����뙃i���ȈM��>tW��p�WT����7#��������e�b.�.���{&�ꠖL�O`����P�>�� ����}�;W�S0��6d�OE����:OO:�6>gNhJ�i^�	�%��p�2LH�us]���V�qD�T�FC�7��c��K�V�O�⫢~�N;
�z�d��ꎬnr%xQ;n��șp3Hʁy\@j8�ӠRm�7��� E,b&,GK�.�wI����R
�k�����@�u����֓�gVM�fgO�9�����q�%��f�$���O
�՟`���6�	.���l��kz1�TͨvԬjWpϯ
K�]&Ò��M֜�����l����Y	��o%��[Yʯ<F�_O?y�C�p�Aʩ�߯�j��/;�_�=����<K*��̽2Fnk����R��r�$���$�=�^�+d�X�m�J����=|�	D{�M5��=��D�����7)����w�'�H1"�7^�b
<ny�x��sk�)���N��-�����r ��=����Y�����S�w�օɂ`�osz�ux�M��qv�������0�I���c��w�����`�ȉ���� ��6ڱMiU�_:r�:�K��$q���Q�]�cH<ϸ��s}<����ץ_w���j WIEhe��^����l��
��E$�`+��h �s|�@��槀;	@�%F�"�̴g��P�;87�\�$�N�c���Օ�y�����ɾ��hދ�?����6`���3q�~kq�Nd�R{�=>�ݎG�qGR�'�b@A�;D��y��pP�i��z��涴L�1uu;�T
��^��a2_z�P����EQ��F��l��h3����ↃL��$	D㖜M//��F��"�Jt&ښ±!V�	���@�J��ǍE��@�)��"m�.����-��h���G��E���`�V0P2O���Z�1O,�?t6�m��#R�J#��E��ؽ���u��?���(�0����T�%�;ɵ�w�.N���%fhŷ�lӿW�)�*w���W��_yV�
�j��ۋ/��F�9��Z|e6�ͽLO9� x��H�ܭQk
=�=��� �!d�p�-栀n�`�S�st�1�'>����� ����e���<�]�ز1�U�������	UfK�wZQ��.C��a����8�N%�����Uif��S��
��1&����<�J`[�w�fl���C,i��	1h�o�c���O	�(����~�N����i��I�_ʶ4ʵ @���,!����E(P����" n��-�69r�)�y`��8`9K+r(~[��N j ��x�m�z��n��!+h��*cZ�-��E�	1���%$:����k@���"Gx�����,4�itG̗���s��Uy����p!�(S��I����.��B[1㘩9\L�����CD���KN_���WaW��z���i<�I��$�]�r�P�&����ҙ��O��ͺ���K����?Mf�ᑤF}/��xʒJ�h�a\*S�iV4�O�kfO��d��Kx��"I�dp����i앯����X���|�b�Q�{cU���h�¨��b�\�����������ǵ\4֌&���y��S�^��jKu��S�C���Ll�Αn�ۢ��	��m%W|l��ֲ�W�|CH�q�c��v~��^��y݁���E���A�	��@J?P ��c��N���SA����`2�[�����-���Uc�L6L�Ю�����@HùK&T��R�eF2��bÄ/���pp�AX2戭6�h�[ix.�]�j��[����qO�6���%W|mqO�4�)��6p��؝��q�mi��f1�+���o�G��M|�Ps3*���*&�'�L�9��t���*�[&+��}ܺ��ȯg���G���qX$�V>�����w�nW`8l(��'p��E��-䢸�
�9�����o�3L�mK�%��J'���7П�����J������cz�ϵ�\�s�ڴx�vj�5���?i�7�j���qs����l����/O��X�7��g��Ol�[���(�y;��sA/1��/�lN��	�6H�����Dh���+!��p@XY,V�������Y���|���ˌ�|�,�L1'�����8D�h������� �������o!�9.:�F���5�
T�$��������M���)`S�(6װ��S}��>��a|��_5x�UE�����e���@Ӵ�6?����'�:���[N�s���ki�����=��Y���6�/���a�.��UԌ|͛�*������~���zt#��;��u��qp�� �l
��j��2ˌ[�2�/�=�]��.w�����pvI������&�)f:�]�MƔ�}_�����(M�t�ד����0��M�Z�"[[�� ��P ^jͺ��ؙ��:�˄�)kE�~"-U ��4#bߨD��{z�aۅ�.�-�p���Ev����A� �BB/�9f�����c�ĲE�)�!��,���D,��w��H5^�h���t������N�w�bZ�h��W����x���h���P��'z�TR��v�}D'q��h��w�٢���=.c�F�B�	�i;��a�:���5��z6:j��	��0(�����K�ד?��ڢ���G���h܉�z�z`۵�e�~s��g��s��Ä(@*�㿐�#�m�h`�µ�B��T���Y��a�>3��D,uVh��ճx"Ԧ}~ŮGj�jAM��Я,�h�w$.�&>�#�1̒I5��� �,6U�^a��6 �>zM�&�z���d(86�4w��}A�m��\M���Ԛ��b�g=��T�,i�#��-A�#g33	2贸�ε�<Έ��w�¦�ض\���A���iR�Z@���c���CH�TI���!%-`*��ߊɘcr/A�E�`1�+A���g���,�c0<���P`���WŒ+����v�u�VɃ@��1Id�t�-AG��gn@~�iFy\My��\�͓*��M����xvC��QAܶ����`�g����-��i�JF�2���Q����;�e�s�F�6J���5}T�}�}8�i�W�\q����4cc>���'�����hͰ+?�̒|*�H���eG�j��Ý������r�j ����۟@�EBS���{��V��/gK��;��/*֭xH�:V�SVǶl0�X̂��ξ鼯Ev���!��&=yc�J�dʮ-@�Ӆ�qr����,��4W�C�7#;������ٍ��NS�>�|t�{d��D}�h?4Uy�A���WbS'���ܩ¨��M-|g��u~A����[9 �2��;����������'�\9���а���`l��m#p�̏9E�ǰ��1���5z3�������-`���{�/�2V�|��͏;�֙�N[���f{ R3����Cv8>B@/�3�b-p�13j�܉g�t��N�^�����AR���싡�(�� u��ڱf����4ŋ{�2�//��s�� ο����e.�r��d�_M)�Oڡ Uq���� }~PΜ�'��t��y��Xa_������6�m���vefj�=��ݢ~��k����3����E��y\�����I뵁�[�`~�PW<ٽL��p
��yR7E���C_^���`អ�����|��a�3C����pJ-кy�J������X��q��
������ӝ�@���q��Bf��DhP��g�'/$��Ub�:;%�0��)��/��@P�!�J��u����8Z��$\�d�wǁ�k����IȞJ���g��7)yd缒�Y�-����. ��eݥ���ʭ,������_Q�P�%�Hz��G*K?������E-��N�7��<N�������aGC���d#��m�~��ҢdX6�w8�K"|��U�0�&�S�T�Z������6ДBRJS����zuA
�JP��4p��W^����-�q�1v8���V$�!�_#��g����Gg�r��O޳c��4"e-5�f���5zW�+/��f�zzJ}����ͅ�3����
�a*�� �����s 7L.-�Pe��'�]��ྊAj�-a0es�-W��g+m�ի&(�v�$���.ƩU��,���Wz}����G�x䡶����32Y꼻l>��C�	GSD+~(4ōt�Gm�1Hx�e�P���d��Ŏ��C�td�36�UP��a'���\ԩ���B&����m� �� ��c��Kc�\Đ'�D�n����Z�<�2����d�����;΂&��Y�a6m��bE0��t��q���a�š���	�����r��B��VF�i[xT@�-h�9�upiB�����>��	(l�%s��8
�ɤ�����eiҋ��5&ʷ�D�N&PK���vp�D39 �W�)r?��r�$F�#c¡��*��[��42:���Χ��3F��f99��}l~�X���~^xQC�˼
�G���V���5��qW���Yg��mbc铜��s݋ p�͈��l�z2�M���V�M��9�yڤ�:7�U���a_GlDՉ�͚�GF������0I�~�9��=Bݳx�I���j�f/Z�%~و��\����IѪn�A�7:��$Vg���3���]o��8U���@9�B���UFiq� �f��}��Dߠt��O���s�xR��ݨ))��B�����d
_���""CW��s�	4��T+"�[�:w7�a-7ǘ0�/sSz~k�G:�p�E��@�_��q[��ì���*��)�t=��ɾV��fC�Z Tˢ)���m�nD,�f���`4��%����@{&=F���#��V�����d�Bg����`�<BQ�a�{����X�V�2�k%��N�<TA��>H�"��2�1~��w����'0�HQv��K��^�Y����Y�0$�;(^�����k�ߟd�����$�%O��'ا:�a��K?��� �l��F����uF ��Q�ܔ�o`�8���u�fL�ʥ��2#�I��-e�U]��3�8�ކ�ܩowP&լӝ8���� ��6���/m�6�T���u��R:�D����O���}˵Cl{F��_-���
:���n2����_��-�#(��1]H�XnT��<��2��-�a�^4wf�r[C�6U{-u�CY��k������[�#�܎��Z���(�sQ��ȵ:K���3n���Rt��)��-���Ғ0F"6��~��������)�h0y�/R�=��i���N�n[����XS���t��1���<����������0˞�B�`CؒӭJ�WI�Vw^��OLC֑4�n�c��'�cf�]f%��lQ��H�'P��8���B���/Y�u٪t�X8��f:���J�P���>$a��+�3����<!3X�L����[�|j@��߽�}��U#�\��q����f�}��(Te�=��r8��!֒�[ 7~G�?���"�h�A�tn�9�W�1(�(���OyxP R����t@�j��P�v/�^%'��?b�����	cM@����H�>>��oL�),q��0pt��V��k��e]	oz�KlKQ�B�X��'>�k ��d��
1�/ ĺ��+z��e=OZ2���vf�������� 9Q�9�� Z���;0:}b%OOj�%'��w�h;�k*�t�o:�d�v�������rCU �$p������v���*�9�	$��G�2��'��l�Λx���i�n(�t,C�o���b��/^�&�k�A*�Qd!O�,Q�9~�{�u��T���ȁ���̘�� i(��!�>S���k��[f�>�`�: ��yv
������(��x}����D��-��P_�F�\�� /�i��J�I�u�b�h6����a$7�<�^51ϳ:�
?g
]���_�Ja�рt�T��c+T�s�?�v�����uD8��<�9?"1�yE��s����ű^Ή|���k&E+!v�{�1������;����W���T��7��f����>9��)��ϫ�!�O�ti���td`���:4�^?�K:%�t�&5�t�v�����ȳ���쉇Zo���Ȅ� Y�P��\6J`����+FW JVE��z������V��8�����P���TN�L�ߜl�3�:��2��!����_�0|��e��s�E���hF�73�.�#x�!
1ѝ
gA�����$�Xl��1qؖ�?��8���K��wݖ� ��Sv=�n8����Y��iP;�T�_���Wm8��=����C����:�"�j�͆��9�v+$�t
~�����ܴ���pDʕ��� 0d��g|��k�z��	�W��2xk�Js�od2��v!��.ƹ>h|��u�;6|��NU�
1cLa�zL�J�qĠ�C"V������a��m{���r))n]�̨������l^		�ν/��S�� �K�6>�������C��c�M����s}��;C�ZY�sZ�<*YQ��dTG��/"?���>�?:��1&�3rI��P��%�=�Ԏb�Tlˈ���;��=&���5%hYar��a%��z���碭W�q��~���f@�������d���o:��?ca�ת��CS��C��\��j%yNw̏+�����MУ؆u�~�E�M�ȼvO��P�|W��j{t����Pɠ�}m��:���8I��vg�t�(��߶~j�#r�F��g�+Զ��=a!b�H��B��e��bP����l��b��O9B�jy:�7G[��T?A�l��ܬ��v�x:����79��͑�>�P�	�tRvp���Mv1^�"J�׻���3`�A ������Ed[���u5kM#v����'C� B�)�,���� 7��<+� ����m�8�+�f�d��@]*Og�ۣ����4<�� ���̚I�����k���޾ :�:c�^��0B�,E���jR!K�����^>�����lb҉�nC%�
��lRtPx�5D�g$m>1�*���Z��8��˨t/��w, 㷽]&�ͬy��D۝���8��gM����&��̝�p�'����%5�9g9�ض��;bE^��������6�J��c9�tP����d�GYhT~�mr������|�&��b�<��}��0,��ѝ �b�J�@��T�
3B�/����� �j+2��=����SF
��t*J~
B��K
H�ԧ��{ʻ!(�A9�bW�ev	�^�0���E{{�zf�%�{>��ǅ	�d:2P���?��*��불�h��L��n��KJۺ��qY?��ׁj���Ф�>2�Ä�����v�;�`�G�־	��d�9��94��r���Z&o�o�Е��Y�����/���a�N���\�!|�Y)k�U�F�r ̏��/�3��'�6_���'�bR��G���y-��(������ٟɂE8�͟�ڔF�@9���;S���|n���ݱ'��awUul�/!�5 jԻ}�9,3���0�� �i�?�W����x��� ���.���E6$$���{��� `3<7P�=̧LEO�IM���	f��]ׇ��A:�(�N ��I�!]��<F\�5U;�,.{��S���1�%�3��*n�@�%����[k�p���Ք�P[<�M�x\O�ie��>
�o*�1r?��U��cR��U̮��$[3R�0g�-������G�r_��7�����s�s����H�%KmE��u�������;'��a�s����*�T�O�W]\��/~���Ts��ڲo�QtF[{���>|#�	�v_3�D�'�ܨޅͣ�t���UFYK�۴���S!������<q�OHt�Qj��h�v\�`�����`��IO-����=�-���F��4A{��+B��1�����F��Ք	kb��{�P�{��؛d9�|u��vuR�Ȍ�'�$��)�hTh�h߉��ba����w��M�%�>a��,�M�P��b�t�v����:�!C�`g���)h�L�*L���"�s���w�-Os$��J ��6[u�=� �x�5
rfȠ�n��Ò�CT�=5L8�nN�8��2�R�l�|�Ip�^Y(��^��m&t�Y��c0v��-������)��Rԓ��"�Dn!��V/�e�˭\��Hf^� ���g�M���v�8qrQ~�(�����|��f��E�9
ű�J@�K�Bk�ۀ#`O�Ha��V�R��_�x��0�|@�|5�	ޓlHp��j�Y��}�4�ڊxhQ@\v՚'C�j�v[�4�Gr갈{�~��:L��h9�;D�i�Ƒj�d4��8��K�#FYh�qfѐ���ζ9����.L��}�|K��sw=�_)�y�9/���٭-����A��Y��M�b�qpp(�SsG��L�Kz]x���wX�\ A�<̙ba�<F��N ƩѕHq����#q�����k�!C�:�6�S��X������l��$�z��h%�'b}Ｈ��iv�P ]b�s�o��\Hy�{$;�@F%.����XQ!���a�Bi1�"��$pa�Y�Z�[_�)�/`k��Ie�=�!?���TK�J���2�ϭ���s��Q�X���dB�cY�)2��Cy*	���M�P�*�A�*�����]'�<*X�7�Iz]���4t�����ްy揬=���P3�L��?�Aq{��e&+)���4W��S�"��V���;_V���v �ޖK����;':xpƟm�)���e�wn����<��a\~���"(�z����m~�����xe�5�Ru~�
HR�RM���4���|�;ع�}@u���t)�&׉ �`ʷ#�p�']���9��lB�¬ h�֓<�����+czq�t@�@\��_U��U�g0<��t%:A��K�v����9~�8Q���h����>z���*��u���wϛ�g	ZDE`l������H�U Bg<k5y�Ԓ�#��>��&A�{5Ma����;	d':�N
�鴔��>��\�{h_�M�����WI�r:���=#KL�N����Q�F���ex�S�w�ܨ����R�h�?B^~�(��|.��f����C�
cDbK�'M���ݘ��Lw�2t�E"Y��N�K$Ylv#'��p�����f����ȟB����T�|�8a���ı�r]�����"��I�>I%�"�tǹ7��v��ƫ�f�4B!i����:DtP�M)��,���I>c��0��B�Ҏr�6]/���8vM��V��c�&�'
�U2������6��3GgZ �g��a�؟��<�F5�ԄT-4\,��/4a<yol�d�ʝV!Ƙ7D�+���u�йP�Z
�4�=�mS�^���;�L)�F��i����Φf};*�kR_���/v���z�Ј�fc�U-s�d���N�n�y��T�-��ϔ�c�d���N��SL휗ZN��;����X���#'��3���h��+klp9�߇�_�),�dޝU�x�#��y4�]r����Q��1<^k���Q5����Jy/ � �1����ثZ�UH��:�eu�"�u�'_��h,�<Pl4=O�d*%�)$��Ұ��3�I��j�٩�s�-��B�?� e���i
�!�g�D�������-���a�!3A83�>��v��?	��iH�U��qC.�9��P)\Ҹ�<$���}\d� �ea�GI���&[�}9�ER�u�eyc�m��|��1.A��6�@��ʪ�Dd��L�^���PI�$D�7ﴈъ�y%�S�-7�޾�5�c�|G��� ��پ3QU�G�o�;�c���53�rV?���n[bB����eS�¼�N��q���2����<�=,�%~)`�w�Z2�݆ף��{�>��\��Ԓƃ�x����K$�����0zh�H���u��W,��H��z�/��Im>yڨ�Q�^	�uu`D�_��J��G����=%�5����4��=�����e�:1 �rV�4�\�v��*aƹ�RMq��Q����lp�2|#�7�i:X9��ڏ?���{FՐk�+O�����{�
K��-"��{f�>@���yHLI�
�k��ϣF�	'&�I��	�K��|�8�.��9����)����O�I0F�{����'���1�	��!�.
�T�6�Y�Ql�A?#W4�4�R�h��bO��Y�� 8�ӳ��Y5��8��%�� ���J��'x�� ����{JC�����i�-�����ȇ2�
�{�2�js�yd���hf��G����d��������2a��w)�^m��ѷ��U:�t����ײ{0j����%�Ji�.������T������WЎ��Ѭ�4%�S�b ��X]w2}��m���[��!2fJ缝>��	N��C��UH��q2�G��������-`�3KQ��<:=x�e����l(� �}����G;ó���M�is�we6����1�]�$MAu~�˿R{˪nɥG�@DH,��<�[
w&qŚ�'��Ж@M� �Q)�>��K�"ݩ}A��rgWB�W*`4p̋g�ޏ�������,������~���N'�{'/�A��.����C�:n��a�El�8y-�1���G�ϧ딃P���-
����o�٢f}��z�]����I��L�+g2���s��%c���6h0|d����/#a�j+l(��*���G�u���j����r�TJ��ϞA�7�Q����F�j6n���I���C<��ǔk6�P�)�.�?ƫ�\�2�����6M���B/j��Nŧ!2ي7�;e��c��y�(��o��Z/���蠹��]$סF�]����Nn{	D�Q*K�x���F��OC 7�w�
��Qx�渙�.�8�;�������FlMF�ᮒ�F�����U��t�Ћ�3�^���0f���Ҳo�q6o�""ez�F�.^uD�z�Os��SȨvϴ��Z5�uR@����(�C�m�AZ���lO_ h�j΍�x�r��e�4�n��P��X���m��V���Лh�(8ض:�	4�&�Fc�i>ӏ]��Z���]��u׍WsG<�w�~�r�X��i�0��d��Zg�4eF\RXg?XϞk��`l{����#��S�]�]#����Re�����a*m0/vT|C����'��~�Rl��H�az����jn�����nXɋO��r���s��d[�!BW��6��E�Zry����L���(_ʈ�w�ZL���p���RK�,Jy���ayu{����T��at�DS͡SXrZ��
�D�,+M8:b�Q�q�nrC��N��d���C�IҚPm�C���^�_��2���X������b]��H{�P�x�{Q"�:"��G�K�O8̎V۽|Ľy!����M�i�|�U�Yν����U���|_�2��sf8w�;�t�(��$��� }�ӕl�� ��+�9�窸����EW�V���J�NE��e�S���(BC��O����(��CVݗ�W�Ia$�y��_`f�&丳���G<:�/�齒��9�����Z� ��N�����9c2�������(W�9�R�zZk:m����s�r9��!��/�e�.e��ֲ�������E=f�̅�ԗ9h�EI=��mK��*~�g��I��ۑ�{�����xQ��	�2��S�w�����҇��\T�9ߧ_\�^[�g�!;���f�Ɲ^�a6R�K�wl$�Y�uЫ,vM�;C�R�����
�#@g�F��D�q}K0OT�Lvb��v��aݝ_�x����e;���\��{܉X>0ށ/�b�>9ʷ�SB�u���_�bk�hy˔^>54U�{�p\����[ɳ �e��:�CJBG>�t}v*`9�<n}M��������jC�|�QU�a���[���D��J��K�u@#Ǵb"��"�C�J���*c��9���{��V�怣��}�9�^8f��r4��
n"����G�1�c����3���	����e�6|���D��ᜪ3$�*�j���x����*q������{ڋ��*t:k�򎠕��@u�\��#�uM�n�y5a�g�8~��QG�-&�C �À����/]^��R�����l���8�"��m��H���D��hm4�Ux
���Z�ou�=�="4�4��Pi|!Kfj	J�
��'3B2`3�nA|��}��FÅnFO�t����11�-�<��dx���q:�眏��x��Ҫ˂I).�<�x��{�X����Z�ށd'G�� ��DKC�e�9���ķ�J�_�[_924�BI6�yP9��krGi��͓M*J���Av�	į�ÝGHJ�2�wh.��U����?�����-��B4rj����#<��}���@��ǡU~�aR0*�RS!�A��X�}��Dz�,��s��i�±�#�b��"\~s\əOt�ln������/���z W�����m�jc[�'�mPY������sE��_��z7�� �EolD.6}��Ï+�V��0�\��o�|�SA[O�Oxl��5��w�'�&O{x����'5�E�}����>	��۱�l���4���T��@����-Wy4���b�駱�~ �	����:���j�]�$`�Y�[�аx8�����y�FǤt�e�k��Qz�&����U�h~���x�0k���MK�FQ5]��j�	kp�x}D���8;���.~*{�_�T�Φ_oӛ�d�j�0=��vc1���c9�yY(��[:B���Y</s̿�!:}Fڂ�Дh�B��c�061��E����7_&~ ).L9��@�i ��Nƾ�����aV��;&a&�R�N�^�rVM�2;"�ZԻ��ـ嘘M��]��|$�0�Ș������H/��^��#���=u�w��+(�	�� �Kt>���@����C�5��I#��V�>�K� ����L��@o�*f�491E�� `�� |���G�"�����vU �����3>�
>;���E�l�!d����)��U=Ù���aq��E?͝�K����-�B��׾d�/&EY��[e�ٖ ��<3a0�&(��`��pe`�r�y[@X��	��"IW�?p�S��v��J�C�V~Ep��b�}�Rh8ހ�dU`�,k�:��F��殁jf�i������Q���\	��7��80�U�]R]!jAZ��ν�5����
�Lt�Q�B�k���:�ʇ����zGC���<����%���8��������؅Snbr��r~�:�Lz��S�̯��.�A�;������s�7�҆���UGՈ�S����E�яx��_��֑�ۙ�L�漜|��ZF֟�EN��j �<������jB,�:��*JϽCq*_��K��AYh�RG�o�^P�2����f)V[G����S��L�	�d׼dW�~��Y�w�Y��/bV��{W�
�}���e��Ӧ~�on�z�	mL/	Z��F�Sl[s*3*��`�����I�G}Ӊ�Dkj;Mzpw�)1�〈�Hң�P�Z�o>j�m1Wg�1w���|�ٙ^�te9e֎B	~i���U����}��-1U��J�$�%��C�}�A�!��mc�	ݒp��h��ւ|�a^rM�(��q��¸%|Z�Q�_��Um�QD��)��%�j�cyQ~��
#�4��v�&��{��!\�u���P\�ڻ?�k[�����ט_�h%ªA5-L{�@@�x�
P�  %:٥#��D�ѫ�>V7�멞f�[B��ϼ%� �K���$���м���(p��KJ��I��I��������}%�����:�sf�E�e��� S��c��	LcŁ��G0Ǯh����.�E�!�_�O:�C�0�bRv��@2Y���)pU�C�H��c;!~���x�Z�-���]��	��f����f����akｒ��7�9ה��[�5<1��I��in?��9�f��P��萦F����෫�bC�~\!��L��w&T׾Ė�����C �|~G�#`W������*	����r,ȶt�����z�j��F�<�OT	jJ�^�LI �]����@�^F	ք�	*Y���c3��DW�G�
��X~\���;JЍ�Í%�uC�����:���_�K���#�p~�S�!��o���.���_�?4�/��F��?m��49�䰱9C1�C>����G-Oh�nU=��_T��J��	|�Rj�OPQ�#�>��t��0vB���\x���_�zk6O���2V`���:3�L	Ơ1��7֑�ܰE�(T�0�N�y	YY��*?r}�����V��)U�S۽�@�v�zt��]A4��%�}�U��-�LZ-�d���w��ny��H[q[�v���*!k����q[�#ֻ�x]���H�h���&��#�P��R��7E��X�D_�W�
�XD������N���9l��Ĭ��
�ɉZ�V(n�E��P�{w���x�X���z
�и�h*vX���r�}��9yLO�S��&<V��RC�V�a �����8�����E�����kRY�)9��2n���h؁�H �wQ�|N���Ӆ��l�Z�}��J��]vd��Z
�y��k!�.ڡu˗��u]u{MZ����l�x�4�Sl�~DX�׭:��ܱ���n��D����i}�®�z��q<�-�!~�bX��ӹ�{%Yb
���aϽ2��g�r�ܽ��V�J�n��B�|K�M,�@�9�*�j˧FO�o��
�Cx�t��l\�LO�Ҁ$�H�*�߽B=������^I��	�r:����Һ������G�,�
���8a$��|tc���(]ձ8�_e��µ,� �t\�i�+��Hܷ���3��#�����j�#�u���$}� �h��]��&��.y�������lK�,!����jݣnP�	�cF�j����W�����W����ga�A�����C�j�KX��Үr��?��_�Q�����;�qn�U�J�y3�]V����bO�v��5����Rc��T(:�>Q����_���d���W����H�߀ǲU�5�s	��_ ����a3z{�n�:��Rs<�b�����#���������]Y��ğئu����V�!0s�ڃs���`ɤ,�id��07.��������EBPN(@S�3��]���5-Н�3$ْ���Ӹ"&p _���kj�f�x��c�Qn* �AU�V
��Q2J/�r����hơ@H:$�M����M$��t���v��l�)������NJR�c? �o�t7��>ۮ?���rȐ>ɔYEd����O�0���t��p����B½���8����\9ሣF({B��}�j��h�fDQuߵc�p��} ev�
Vq��Oן
�b���L���Y��s	yH�o���~�B"�5��t�� >����sp#w���KZ�G��%�ӭx�����k�~z�n�x��t���c`D<&�1��t� �Nŕ�rR�VnA�.��а<�
�;_�Φ �o��>Ƙ�9�Â�y=Vً�����[�=5p�16_XHR�QG{#B%�ɣn�#��IL>ls���y���a�!�U�jA��,��܊���M,�۔Y
����^�:9S��E� �3��c$�	mv�An䠑�%G?�����g=XįdRl�e;s��7�g�~5��t3�<<f0����C318Grn���A<G����n���G���e�!���.#�6x�#sCü���I}��5~��tS��O�]})>�N����4�˱r���E��Ӽb�i����k�V�C|]�?ނ"n���9Vt�����H��X�����T�?-�_��e�\2�h�V\|�kuH�~c��0�V���~���	 t�>�J?0��٧7��|����i���O�cB�G� �.�g����I��oG�t��]��G*b@�}[��v�A�c</�J�gh*�����}7�C��a(b���`�$hq���R��Dhk ����@�T�AM��!��U7=`����u������Y��]I�����d���L�"���T�������*� `�_ijL�\����8�j G��ژ�?����G�y	r	�؆D�F���ʫJ�֔b*f8k�z<q< ��
��_��s����9zt����O'E`�����l��3��!��"�����R�:jP*$���]��gj	��P@��o������5�s��qȷt/4�!�zY�):���˗���n��:I�Iȓ"�c���.t��Y��f��Ӭc3m��1O{�f�.��N��)U�T(L����CK.�m��/���@t���4��7ƻ���?�v�A'��q%WW�.��;��Y0ž�*���
�@|�%�쇰�d<b�W@���C	�Qɞ��{��(���F_�5�ZG����H�����˳:$���J�e�:���h����/.k�xR�}foX��r���l0�yޡ8�N��G�*����)��;����v���R�J�� ���qu��J��So�i!�'E� 5�%_Ŷ�5;N5���c�ƾ�\U����RNq�*71�^�?"��^���tz	j�*)ۇ��1�K���3Y1�G`ݝP�Ȝ �m<μ�ҩ���6���͏�U���]�3c�Ku��4Ե�B����;��J����ITo�����)�Z���L�Cx7d����|pN0V���\��t~�o�c��)2gDn�Q��6cYW�0����SY�
\r�n�gIbTV@��$̸�!%����PViKt�yTt��J��hNdi!�M�JF�+��֙����a�oI'�(�#�9�߃�7�"cSqP�ot 2�-����G��$;Im��+�T��1�cD�R��	c��{�W���5Y"[D�a��(��Ů�x��i}��گ�K��Ef��-�`m��+��v���s��-���^��I#�չA),]f���G�rt��wZ��n������D �]JB�����j�8)��f��S�:!�������	���30G��q�>;�\n��n�uN369$6�RWw1�����.mqf^�g�j���B�̍!���E�oS&@b�����e'X�UG�qx�D�g !�\� G����JUK��(��,&r�ړ����L�cV�C�����§ݓğ�Z��$����"0�x�KÍ,�J�c8h�W`����9+ "�yza�1S�rj��d���x��"�m��^{u14:O��Q�!��_��J����u2�������rJjƦ]�� � [�ݵg�T	�B����XB4|��: �<[TC��D�G��e�On�oȚ�gޛ�1rC�T'����������^��U�﵋S��YPF"X�����~�za}~��r�K�Ƅ��[6G�G��A?��d��K��=M��N>}' �L686��M91"�w��~j ��x�� � ߍq`�7AE����w�6Ѿhxh��h��si4�Z?�D����7��y�57��?_����H����,��uc@�6�X2�A6i��`n�����z�k>�Eځ6����gN�Y�o�8�#Rrb� �@W�kƩ��}?��)�M�=U�P6��71�>��d�hw��{W8��i3�����iJE����Z?��#{�����hw5)~��V�dCD��{M�տn#'��H�jT��>` ��~I�lS^�-ROP�2���]i6�H8�N�܊'Vr�
E!c�A��Ǻ��4G��D�)u�5:�.x�)j�P�����^>�N�H��2�Eu|̗�$�C8�ܠۈ�~��
���6�� �{��V��% ��Eˍn�V��t»k��'s�`b����-�H�b!���>Y^o��-l���F1�Ml]�ܦ� �J0���=���tԢK�=E	u�<�>S��^깘���=��Y��F���9�;#��f�*ܨ�ϱ[C,ho��%���{�����H�Fm�w�Ŏ"��=5�@^����2\��5�Ŝ�؎�����FQ|(L61��i��;gmu����Pc�D�8SƔ�Ib*��T`������"!J!� �Z�f�2�Z���y��k��%�h��XN,t�k��:�fߨ��M
���	��\-����s6�!�"'0��hnd٘��y�Zc/�og��s�`���;���O�W�ˋ�S�Ɔ>�HK��
��&-6�A�1j�T��j������E�)@�m���p�JFoIuka�J��;�kz��P���:V�0�F�k����6�0�x�G��np�f��b���4k1�v���٩�qCQˀ�i#�Y���|Q�ϋ�y��M��B\1P��]�,q^ʵeyV�wv�$0|��5j�m�T|:��N6E�j���&d�{c9��`(���ijE(��O^����'ܑ��R� �7��d�Q�G+#x�غ~���� ;uL%;�7��O�:����]���(} #O��m׍�.$��l~)a+`��j]�gJ�
�r�9^���x@��[\��0)�����nF��x�����&:^n��`�,L�v$[G�� �a�V���2ۆ�*��-�I4hkN=�2v��J�K'�:\�U˿��3w�d(ͫ���f��ꠙ{W3	u��?�k��4^ wf��ɬ�}���f"�N�jĹL�EW��̼��dڄ�Z�[�ڢ�����e{A:��Hy��N���o�3���@ٮ׶J�(�bs�PVhk`8EU֏.��k��'���-c�����hЈr�5��񋂅s[��SZ�Q�QW���e�Ii�ּ
���uG�,��:�CO:5����a�Re3��s�&z��t�J��W'J���G!Jv$#Xd�D���{	�ߖ��H]u�lU���Pqd_P���(��7�$Z�t^r~t&�x����HG�"�ac�$e�q��X�ܓI�wg~9����d��-/UK���Ѳ�.���w1�"�ʰy�C͉`H��Mk�(��5󄿎;��|��-}GQ�RB�+��lW�8��|����Gv9g��	h�~yİ	�+'�&bC���O���[�Ң�C^�
�q-��Ua!at(HC���cث{�c��Tfs)H��b`�E �{1�x�|����7�s�ܪ�hwn�oa¶��.߇��Z��72:�ӎ�x�č�����7GC�BOWa�nf���1oyŐO���~2�����^���<s���`��Onim�~�bӦ�@��NY׀ie�Y���J�O��H�l�ӓf�d�v9�?(��s���j?Y	�Z�ܮ���oH0�Y����cz�U��qɐ{�``ߺ��y�/�E²���� ���@����F(SQh��h0/(M��ys�Y�[Z^�rdb�O���gP�����~�4�6G�����F8c��O?<���nr-3�l6n���>��	'�Re�\�|1�B��W(�!ζ�9���e ���-N����3�k���+��>;9<�F�u�CZA*��s�v\2��Kgf�ki��z `�K��+Gr����,�i߱���P�ɨ�:U�_����g61�M���}�ͱ�c�´(�j��HD_��g�;n2½�;��#��5^����ި�Y���@W�B\
�>h�n�a[%���n�ܡ.�Χ�+�e��YX�'��T�p?���^�Wa%�rxu�@k��y�]�vx�Ƥ��G ּPW�,�ē�����'�	wk�1�� Ⱦ��G�)���iŭ#��5��g���?�!w�����=���b���,*�j��r��h�Py����3s�}j�A��2|�T����Ḛ�7cS[%67k��V�qQ+*��W��
��z�Hٺ���`��Q��s�j����lS̏��-1���f!|�J��7ǫB!�r�!M�:$� �����k�������@�ǥ$Yu��р�I���+��xzI�˽k��1|��PLw/lYͦ���)��R`�7��9R	�{&K%�C��|��B�B92ק_���u�Th!�x����y�Ep1Z�8��T�}?w-�j��x��h��/9I�Ѷ�U�g�utZ3�S�P�7�����{lA��Dož/K2�[�
�dKrssM�������R�!"�!'�b<"���>��-��ܘ*��h�r>�2��� ��N�u��?,���U>�"��Px\���i�".����pXxm|6�8��	�
�G05	�JRa�{�Q�7N��U`\�$r��h^VΩ�K�Q �$�'F3��t�Vƈ�<��"[{��LoAe�&���`7�s\t��LΣ&x{�Ľ��� M��+��}�v�F��5	í`T�7?�!��p�+�j_b��ʙ�)���C1t��VU
$0'��a ���'�`��=��@�Ul�&��m����g�� �S�6���^�~��3��qKeG�Y4�eNc���/�:�XDi��V�Y@ֿ�}����bw���tFh�$]����H;�P�p?5l�]Cb�$G�� ��G�<O�J�"��PpR�Z�F��0TC�6�b>Z���8<�
�����};Z��e.U����� � ��\�y��_��)G����2�qJ�m��S��:����ǉ��cQ����1w@46��_ŭ� ��������o��$d4���6��T��y��&ag����
�
g��������ߚehD�%��k��@��zBj��.�n�x�h�s�X�Q��{�Z��,.�W��wQ� �Dִ
 0�ܰt4� �73(�X̈�<͠�;��V_��3����
P}�BI��t�B�C�uR�6���P,d?��kv�7���גsS*��3��a�]���\� ���/��r��*{L�x:$�V�g��k&����"��<��x����e��7	��� 8x�u�ч82z=eB7�+2�8�_����+�����,̋}���ܥe�{�MB(_�dA�)[ct,���R3@� ���D|�!�M��n��l&�J��14�5�&h��M���:b�gI]�
�q�7�Ӂ��*` CF�Դ5����nXWTj���5��KnY��|S��=����ѩ�v��X.0�^JXQh�
�څ�v�|�ߛ��OC���:�>!f��@�%Բ�k���}��B��V�|:kz��='�۔*��5��璷�ǲcGS�\�9K^hZc\�՚Wպ�x�vȽz�p�T2���Y'$�ز�LE�TLhbXB
@�oQl Tt�pzx�'�a���*e���G�"��5�3�m`LAVg��B8��^賊���]'jr/ʥg�x��-��}GY9��L���汙j�V|�23��2���L�J��t��<@�����oW䀨��N���P���܀�B�钗Z�����h�h���}B��,��>��T~�{8�S开��(/wo���ÛEA��)O��ہJ�!�����'��q"�O�)D�1��xR p�4(@���E1��}~�Z�4J���ll�"yZ+�<����lI�k���ޝ��b�K�DjH<�I�)>�4O�ꆉ��B���,P�&,W�s���:m����O6�1�
��G 9�é��+S��p�5�-}"Pl�3H�����#� �wY����L�M��~My��M�o��<�ka��Ƈ�| ^l�բ�hIT�w�gwR�ȃ���ڲJ$��X��ɶ�E��� eQUk��"ڽwJ�"&�ʩ��a��K���6�����s�^Qm]��е��:=��FZz� H1Y��5j�L(���Y�	"��q�aջ��&���A���Ivv/������ra��D�R�ġ_D�9/��J��O�|�!I%���ǀ�PD4UO��O"�ة��2���iqEn�^a��w\
�i@#�%ɂXu��˴�:��q�i��T�A�g�6%��p�,�?]��bJ车��� %>�����"; �[Z�g�����RFa�����-i{w?/}���+K���qT�X�3��9m��R����0 �TE��ѝx�3�A��Qz��x̕:I�WxAihJ�D� �������Z��=;�T����{`,P�G�/?�9��a
�L�B���a�9N�'�]/����/�d�E�]SN�tC���Z�&<��9�z[��'r1�����oYp���!=M D�h��j�_�����x%\@,=�I)S\�~�CJ���K�	v���H�q��{t���KT�l=uxP�bH^�>|�.�}4���NȊz��
��+/�-�g�H�D��qul��>�ߣǇk�d.�TN@�/��ό�M��9XlP3y:����O�+��T��=Ft�z�´L-��o�S�'X���-��F�bU���v�̲��/ BW���n���
��nC�^Tk��.s�q��<����ɪ�f+��L��F�uR�i�k�
j�U|��+�DѸ�t5Vp�.���
��v츟+^�`{�}!f_��ߧj�7��f�8mr�죣^a~�܇�,�L�k�}�2��gQ
�2�$��/��<zd��{&ъ�Ir��J�?�BA����D�|vg�j�C󴼼�i�@Z ��yz� �$�aU�|�E��N�6TW�z��u��q�0WPj�}�c�����'rj�����W�B����W��U3�o@��䶲3z
��/�8��Ⱦ�_�L��9 �ڟ&��Ǐ��?"	�.�u���e���<Y�[9�J�� �z�G��;M*�B�N����P҆��	y�\�@$�ʹJu�P�)3%mY?�X�?��s-�yx+��B��d&�N��}O�ri�R��L���$3SD� |����w�ى�T�d�J��%;T�)�&��3,K�����Em����3-M��@K�Eĵ�O��:L���Y4� �#��<���������r��Bq�V�YU��_��Z�ֆ5�͠�(����8���
�� .���EW ��-�3��ýNE)� �W,z�� �"��4���wZ��������G'�쯄֧��)�9
�dGԢ6��0�K9$I�r=��M�H��K���U�-8'��%�&X	0~���,�jjF�˘��D5�S��Z�o�+��������FQ�Jì~
lI��v6e�1��!Ǳ���8CL�8�HZs\ѥ_@�j�������1G�f�d�,LVOGu�ؙcX�̅U^��Kݢ��fs�*g8A"h�{y�$�0���t��7��!v1��;	ݜU��p��[cGc[p�5������9e��
��
)^{,�jFM+?��2��������(էPU���Y/z�c�aE�fl����iVx�+b�ҹ\�[@�-��S2N��&`��Ŭ�Sy	��T����5FJ�$�P���Uu��U�ͭ+��xָd���9@X���WӺ3:�4�W��y=ݠPs�Act+]��d-S��mz�`�^f��X~Zk���鳰�t�pv�7�2�̅G��uw�Gz�>�{�a�m CY-���Iu��"��a݊��\��L���ب�?*Q]�4c-X볽�Տ��'���~H�{٥�x$[:!�7�b���;��I��Lt������U뜰RK櫂ðt�7$����[��Er/2H�T����)�z9ZZL�p�,O���	�F����ʤ���h�Y9�]��
F�̘��]�E�-�nwx�y`�\���P�]��'=����(؃<�'�JW*pU�t	����u�����<:��tӹ�s 4 �R���ֳU�L��7̏�#9��#��R��\��!��'����c%���j
��SN�y���oW^Jڼ?}�l@���/�셮:���YgW��#ܭ�Tٸ�Y��zQP��<��Xq;}�q΃�O���/�Th��G�����w�$�h���;�-��e�՚꨾x�,�����hPcqގ����b���ܸ�;u����g����z����؍�����+����j,�y�A�3��?�>ukŇ�kw	\[
�V�0d[�4T���!�N�~�UH��j7y����C����-���w]ő� U��4y���\␵˽�3���
��Ί�~��4��/O�^���EĹ���*��Ԝ�.t��ҿ���2�s�N�������6~KA&�K�7T��n��"�Up�D�����O�,g�O�x�ܝc@�W�7���Cr��R����LC9v8�l��%cU[V➰��i���xn
��#ݓ�k���c̄({��[�A*&����]��F(3�c�%1���V�n��A���O���Z��:�,�@����ƞ�U=ՉG!�a�����}@?��6Ug�3�s���w�2	l��$m� ۭ�G�����T41�v!c&�����?�Uz_4�� '+Q��
��V��C �>��/���F�86�h��P�.`RS��@���̠8��:u<~��Ra��Ę\��:*�5�?cI�����.��_��$�(��q�5ef�2���Á5�SU��6D��I�x�H�=���U;kj6f"�/sB��ԃ}Ȝd��rO���1V��d��wo�!x�dl+�^<� f9�]�hx���ʈ�`'�d{n%t|,pk�������q�������8;���sl�^ß�����]7}5O7��4�c���;
*�\�&3�]!Sw�E��6qN-�A�s�s)�b�t��`�� ���u��cb9y|o��q�z�c�l���;�v(Evi"��(�.^�+exìJ"�L%�Jmyڎ��dȕ��r2��߰�FHxMI��s���ͨ����;�� Ұ��xu�����E.��3,$W����j�`CO��7���L��=�\����,CfQ!5�L�1�V�Mҷ�ٳ�O��,��l��'��-gV�����;�4z��TRM ��~�5�5E"KbW[&�� P`�ˑ�`��M����r�q���zy�9ѡ/����:'Wf��)8��?x݉U|��!m%N�~�鴦�4]h#ԣ�!�PVl�f��ߪ��v�� ���+���FXm;�s�7}���v�&�۹-�e.A�a��^���Y�U뿗Y	aJ��<�J�E�=�9�VJ�g̐�w�͎�8`��4�q��Ƨ�؍8��&2���9
)�{��`���sW��f%P��0 ?��/`EÂ��R�%�Z)g�F#�i!�J�����e(��9��!>Ҋ��^����K����*�jO�a�X7��JS�N�F��U9v����i��(���\N��)��x�>��i��6�^V �����Frr������<��9Ԑ�N�)		̻�F ��H���]]+�R[����t�L"pAx����/-�s�z[E#k�-�)�G��-��#�Q��x��xJ���]:�5QG4|aXp����o̪�t��
�U*�C@��zi���c ��ɼR�y�Q� ��ӗ$ώ��f3(_+�e��do��{n.�9,�~x������U����g�hx��X���~�l����|�2~�K��h~�����m<BN�ZgМ���,�J(j�Vd��A7w�x��R3pn!��I�R����E�N4�r㜘�V�[���s���kh��F!b�F������u��r	�GG)��-���Ԍ\��,�t��e�>3yd�:^k�_���6�T9sA}'0�r�Dj�����1Rbi�7����n��;�7�&���9	p?���|�~�~���®���(�*Uۢ�OITLl�J�~���qh�`x�oW&��a�a����G.6�L���x�����X ��f�H)��5sK�/���DHH^i�Yy�qf��IyOt�O�J����]�\�Q۷����<��g%1,K��F�a�x�&y��H*���
-�E�u���A��i��J�J������`�n+rZ�ɴcχ�:"��~�01 �'�t1E)d����("�64�D�N��f4'��X7�^Է�Р�+%�8�ODZm��0z�2.̼�����U���XT�1�Ǐ�UtUط�f��S�=Q7j5L~����κ�˭҇2�j,�(Tn
�ŗ������eu J9	=I ������x� �QrSxY�5�X�Ռ�~ȩ�1����#��G�9ݥ�_�V�e|� >�/3Ɲ){/� b�mB�$  �NR�0���$�y&sX�ڽL�#�B��3��^��v`n��J��:��|F��}������b���w��0���t���9�D��nha��NF8U�hm���9#U�˻����5��@���ϵ5v`{:G�O�͛���|A�W�k�X��h��P�._�1�X��\\�����|����VZ�E�Eg��>�D��4�2?����Z4ׁoh�cń�M��ܦ̈́�~�Dk�u 9�l�^�������	��
	Q,K?��v�l����;�ڂ�;�-5���*�S2���1"J�%P�}�Z��M%ɠ�L��*:2L���l]{��7I'�U�}��aԖ-�:���ib�(�iIF�����/8���^ɦ&isyHD�>Dcd���V����~x/q���?_^ݯW@	YK���DQ�u��]�[�O׳�X���m���q=����:���9���]pR# $r��_����ھC��e};����dƕX5��J���ID���(� 9'�XA<4�5��m|n%�F�̚p�E���``�0���Y�����^����,�`���`�\E�¢7���,K$P��iq�r��S��g���Q�Z⽚O���8�9 �Y�j�ݵU��#��A�_�l�J����]�$��E^W�[�>�E��Hx�lku�u�x��:�'M���u�@ �;��y��X���Ǵ.>+��	X�oni�ɼd�*-a�|�JyS`��p=w�<�!���9�	P�g���ת<ɡӈJ7�o_d�u�	���.A=�"������-�,�8��M�_a�ą�,�+����NuoӕPGUIY�c/`�a��(&�ߔ��BRH' JT�8��@W+��"TbI�)����?M�C�9O/bf�;2���td�����&�9�&x{�m�Y�D�w�;�͡2E��Z��#��+Η��d��<����c_��b�z��8���)Z�L�^�Kw<��E2jR^��j�ZŲaZ���[z��q����n���1�R��(�	k_�PYR-�鹲�C��Ǻ� +��W�*���J�m�Hg"U�ݚ��T��^����|\2w���R̞A�uz�~鹨�̻���ws�y\/F�qg�_��RI���>�ΐ�d}s��!���!�����~��|�t)��Q��D�}�1���#��F��J[~%��s_��(��wS�#�K�h8|�Ra�=�	�f�K��o_��l��E	h|<�O�u�jO�Y?(�W\(˗uD��,[�w����I�I��94� `�_].���Ǡu�o�q�>c�^m�l��!����p�x��$��Hv���˻:�mJt�W[3[�@��6%ۯs�ձ��t�����BN@U�J?��@hW���<���D#��e��$�N�9���)��2Zu��g;;�_�X޼� 7EdG��]?a3��2	���٦�C@�c:���Oө�b�T���d��<��N �݀\^�:8�����~N�i⪡��[G������?)?�Sp���z�b��kw��]%��WȔ�SZ�Yjyd\�@+��Ww�o���fu]���A�@�h��$�Aౝ��{��G\�6M�Y���wd5n�W�Y@A��l��hV�q'J���"э���Sӫ��{gx�v`F)\�$b�O��4u}wa����j�w|�?�Lz��ykK�J9E��*	Na| +n����E��q���ӣ?C�-����S��La�������v�4�P��U0S�A���ݲ)�M�����C�>�u�z�xˑ��tNT;�����6x�?i3B���ה���}�!^�_��bN0����W&k��L�T|�fT���y�se²�>酏��bZ�T��/O듥�x���`�Q�C���+�^\I�n��.�t�~��JxUfu�8��}��c�1�O��q�9<�\n����Ot�ųF�W�j�̛�1�HHz�2�TD�� f� ��.��d�4�V��1H�"I�TȤ��}�w�#���.����G��&�$�'�*��� G��*��̻�Y�q5������4S�<hG\��͙�;zIm��N֤b5���A���,k�FGծc�q{|��Gzµ���s�:م�~�D��$�@���dK��]�&u���u�����¸tlݰ/<�0^3��������+�}��S��ܩ�ڽ�;�Qk�Eͩ��������U9�:���H�����"�L6��]�26�zv#x�- T�r�27�sg�g'1���j��o�~yݠY��b$<���UP�ݥג�T�����xe�2f�GĚ���`_�4$�̊��&��wm����U�D���UO)-B�S��G$�$ݑ�S�߰ʧ.R�����p�Fx��

�Es��t��Ն<�O~o�v��gtu5�ůR5��ac�������?lݴ�i[� %�o�UX�vzX,j3�ܭ��8 v�OA�����L���;�QW����9�����QG4@�>�-AO|{��~���{%S��9p����fl���˛�������r&>�����
�dVA��4�[ޒ�B��N1dM���d�/�}��fM%!��$�6�u���i��B!E�l²��y:k��>�����ˎ�P�Jǹ�xE�O��(�n�,�#����5�"��b�$`�a��k�1�zb:9�B�3!m���wi��0��}*	����ʷ: ��+>7�����	לּiQ�@�YHw�KeX�������r�H���9>�L;OGd�����d�PDT�,Tm�7�.L5v���~)���]nHT5����t����oO�R��@��u�_���b�!�lT��zté1���A��՟ ��^%_<s���N.jW�VSЭ���%c�e
���:���:��۝K����V�:����}�ܗ�G�.UM>jg�i�U�m�N��x��Q{Q ��
���֠���Q�$fN���Jzo���K
\�R�.'7�m�,�M��BZQ	2��?4	o�� �:?U��U��g�h͟�nFD�qZ�<��,�A���dL�9e�d��u{I�Z�P1+��c�~��ȍ|
��
5hٚ�z�%">^��c�zW'4�l������Ck�ݺq&����`���ц�4`7?g�G]���sm�߀�D���z]�������x��Q��X袂����/�p�5�����9��5�+��aʋ��Y]��M�S|K^e&M��D�������⡁�yO`v�@D2S�u/C-�,�p��)?:̓zZk�u�n/X�*)������ӍoP}�@6ax�o���n�1����$��-�P�� �8_ ,���t{�#��l>�D,�b��� �<@g*�M�Iԓ���ϋ���`��X��*����ϧ���[���J?��|��(�cK����3x2�p۾G--~]�I&s]����2�긫H��,���=,���0�Sl!^p�o�M��.�1�z.� Nc1��c:�k��߃�1��#�B�%l��'Usj�4��e(��.Gr�*�{�=�����?:�џ&�q�fqc�~����8/W�N���_PW�돱���_b]�+^KB:�+D�6%/��l���,+[����&{SW�m����W?\�3>�v@��2�D��z��L	Ei����J��n���l��Mu~#-g��í�x�B��?@�3�_ ��B�v>����^V�q�}�k�
q��V�\Q���]��7#>�4B6m)��__Fc�7�I~^`��[�R��R.�ɻ:�����8�&;����ND&�L���L��8��R��f:*��T�ސ��-q�cm���yD��E3߹啁�o�u�*����;�]��3:�l��s�~&n��kX���}*���Q�4N��+��h �X{���,�|��b�	ѭ̴<�6�VJ�Aޏ2
@
m���%y��ͻ(��b�����`T���{��/��i:^̢pľ\Wh���DǦZ����!�u�U�~�-:�c#�|��j�ôo{T+:�h���^؇��z"�f�٩׷]9&ޣ�����?R;�)m?��ӛ�c�,Ť�C�7zn��+8�s���0���d�M4��`��v�nI��$��Tv֊�!����P�A����̞�|�Zn`�TG�i��]!�L��.���4I����6�����i9�?/��Ԣ����ag䭭�:΅��v���*ϖ+Ll�
S����"mq�[s�P�}����wz��>��(HIK5�GqJ��.R��bI��Uv4j�c�P%	���u�_������fo�T�N�%c4$�<bH�5������CB��^�(��a ��w���9?���bƆ�xD�Ij�+¥�-q/������"L%ő�ep44��n'��t��
@�(>��<�{��o7�Ӯ`��Q�|X�"D��6y$ʦ9�9=.�ψ�� c�m�w����KE����:��A��痏N��ijŦ�<hXW�z5JJ�|S9_�zBP��0��7��1[>��D�S��E�+� (Γ�������*���E<�o-SbC6>$Qf,�Kaci��ٍ�����r��K�k�&=T��������j�3�u@uT�d{t�֜
r���UI|���'Ǘ�rf�4lH�*?q��>�H�8WDg�[	�j���OU�����6f�kh�o�?���9WI�|�z2bn
!���~�I)y[�Em諾%���`T��{��/���m�WS�>)�whQ��:K��6� Y{i��|U��L�'��O�r�|���v��-��^���w;����̓��]��B1'I�J{~�l������v=�pf��iv�W`���E�zԾ�Q8�bq��Z�����[��c<T�jh�e������k�I��I� Ą{P`^��J Ǟ�b䳔Mu�K�Bf�ݴ,j���覢�vn �~�daA�:4����4 �����]qm�E��Zg>���3R./�[�-^Յ��5J_��=� 6�N��kHi�8�&ud��B���"Zz9�`�9F!�x�U��r�A�օ��1�Y�6h� Q;�"T�s�;݇Б��H)�7(�\B��_���s�F�C�Ŧ�5O�~keg��Y���s�_j�Y���I/�0� E������	�kқ���o�	��*J`�̕(�W7cƣ۷���U}n=`�K�=�nplm�r�hK�;rȵ��,���93�By�%=ڞ*g#��BzG����pj3���#	Zs���'^@.�8��L�1���8�>��@�;jF1,�v�_�6�a��S�v5l���g5�
TCre����.�{�9��(P���xf},�N�,�h/߼��[��":`Ub�<#=6mH� N�-�;��H��Y�AB!WN�$��w@��^-�=���-ǿZq!܎a�:�a	�\_ͽ�;�Ṁ�bC�2��= �d����f:��aǏ�`��RP{���g$]�<	�I7l�0��TeݹupU������8� �� ��C6�+�0a���P�Y���j��Z%5���Q�b�1�J����x?�����9�}"?��r(o��B�:iL��l)����~�_x�Llt�DsC��cہ]9��6lw�'ɶ���v\�Aq�ݞ!�MQ��߿Z��k�G��q��F���w��UՓ3���#%�A�T�Ǆ��l֣��6I��^Q�9ש���r"�a�����<tln�͏����l���o����������FT��Y5k���Ѐ�G�*�����$���`?f��BzBE�W�����(?w��Cc�-�����q�2�*#�TQn�
b=Xu(~WZ(���4�& �MJ@�Cpan�<#?�h�A��<-�E��&�)�,:I��E;��昍�|������ы_7c��\�|���zg/�%���J�ܠ_��i�Ъ4�!�e;�+m�����ϕL�=�:-�(���,τ�.ꗖ\g{�>v�0r�/�Ē�Jˊ$8_:�Ii���:��󉯅�2O�-���1�O��{ʏ����������j�l�w�k!.p|�|��N@�j�=�������Dt�tW��u�{�Ѯ����-����a�+EX�Cۉ��\|�5�!@��e�����=��*/����{d96��-���g[bi<W:'�(�*�ሿ���}��dMP��_���6r�����8��nu�'$���������v�}Z.���H�_��H�R?�G�&�:��
U*�쯞���,N�����)bgu��L���4�޳)��pi1��a�#7�KKfk8������ņ���ŀU_v08j1W��{)���(�A?�j��X����MPG6B1'mi�0��w#�At��9��H�O��4�Կ���,�oy��oT&	T>�h"R�m��=ac�Th��'u5��m��K)�������a]'j�Z?uhMX�[1ؖ�/@��hj�� �O���?| ��j'p�+H��V���;KU����r�jˍ̏+?,�UJ�fxZ2ʟ9eI��!)�ɣ�3�F���k�q�x]V���*�J��:�?�n{J�3Z��6NzL��̾DK� �p8(�k����ų�JTg�h\�hu�l�oԞ��hi��6��L�@.�(;a@b�V��!��h ��,��t�Et�J>�S6�S؟= ��mbp�H�h<3-��^��$g}��u��z��V��6�Юǧ&gG���� ��N�y�>�P���K~k��]L�hw�p�ꆦ*E	 %�couQL�������z��Vh[�`�z��Ԣ.X#`-"�$�\!�����#���!��Yoj�{�gwY��`�'C���.����Ĝ�c�>4��f&�s��'1}��U�[�*��$2��P��sD�A2���9I�(���_r�3ն�q���W��� ����<P�-3 ��?��ܟ�p�)�1u����g�K��A��s0-|������@����Tz�`�;�5�S�3��dQ�ӫ�?��
�����#G�[�'�I��L,���FÜ�_H�N����yn����$lw�0�t�AcM4�������ߪX��<��c���yϼ�Kg�����������NY�;>l灱��]�����d�i2-A�mL�B������5Ⱦ&�:�)�N7Ol4~�]	Y�9\c3ȹ���J�[��l`�)�8 �i�I"Z5b�5������,Ɔ�oe
�S4,�21�'��`�	T`�T����/9n�L��$���H�;��H/l 	�͂ӳ��@��فe~IBv�^ڪ�IC�::���*tZL���$k�@̾ۥ�dj�V�k��z)�Ջ=��g����8�}m�9��p���W/����ك������ 9��i��Y,�T��Y�I%)���g��q���xz��WZfx-��Y���'̖EM�:r(�1�f9ϧR?�2u��WY�+�Fj���t}�-O��h�P������ 	�
>��S[|a�K�k���b8�ݛe���L�-�:�4��I���j/v�w��u����D;� I��D�%��!�_�����Fx��V�ʤX�덇�v�wBc&#��ڮ�I�1ySI+,/ �	����XNOS��L&mrj��/��Q�p<z�r�wC��=G����]�['ػ�W
��\���҅T��ܖ�"`ш�f}��_8�|���X�+�t��lI��_ �_M6�=~�4@u�'�$+��Z�=Z��aB�B�����"4E��-�8'�27tH��K��L�2���ߦ�����<} �G��l\Jt������q4��deOTf�GI��h�PK��1_/Z�r
����ɏ*�y�({�#)�� Dc����b)$W��6��J:8Ĺ�������M�0�I��*�IP�+?�D�D�,]~_����b`Bu�1��Չ}��)���N͂�� <y��|vnF�#e9�&��Aw/�� ��ծ�`g�_2�����b'bc��a�8�{�e�&J7�j����f�2f�E���:gV�~�c]c]�r�w�Y�`�=��+:/y���l�(����o���oW*��w)�R\ȱ��o$�ӽ��h�!v8u�t��Q�	_	oRy8�d�l-@i씔E�����Pfy2T�5�&tλ_�k<hD�jMGB�t�W�Hպ�	����(�H�n���IY`�r�aA�@��n{���5J�^�7���	��d��Q�/N��=A����𿔛���|,�b�3E��:\-wm9�Ƅ��6an3'�����}ړ/"���(�!�e���"PK����8ڝ������Yl-G���[ү)*U�/p��2��T�y���b�ӗ��Qws�
(���u��o�{͕GŔ?��=�ׁ�.��	�cT���d.
�2����})�X��?��R#�7ǜ��l��Sp��ԅ�t�i3�����4>�,ag�0�{��V��������C�m�q0�4�����jΜQ J�?I-7X܇;$v�}�R�s���$���TޡN�u�<������&�i
VR2eͭ���EiR`G��awM �Řu�R��l�T{����v0\+32���b*+=w� ,��f1�`���	�l~��'FB���ա�Z��N�dP�q�9M1`7"x��V���A�c��V�g� Rgī=���Lf�����v�kw#��J�q��]CLψ9+l^�٤B��2a�M:Jr�"�Uamg!G�0�g`LeϚ,W���Ke�B�,+$�WԺ���搆���:�8\Ġ)/չx2G��2F�t��z�i�1x�%�w�ޑ�6�|�#����i��Z�q.�6�c��T��]8L���?\p<!����B�i��敱��Ѳ�F��=�VǇ� �Y��9�W}dZ��U���V�ke3��ǽ�^3y�l�� �?�G�X��ٛ��Q֜��������#Z ��rG��ˮ;2b�m���������{�~���7�!�khp�3���n�Rc�."]{6���b�U�Nnf���U�Ϊ�+÷��J��M�N�^�r�{�� V%Y��� �Y0���[O`��Y�d�=�����-%L��sX�{}71ޅ�pOM��FN������o8�ږ�
|BJ.9����ߟ�k�����7���Y�aP���S{�6�>���t7P�/a��EGVz�}�ze�4(���y�o����B]��k�B��8�r≃�~�����뭻�)�n�'�6Nq\-[XL�q���Q$�퇳�|��"н�5k�-n�s"���k� @�=�A�^�۝H�ft(�.�D�%�F��-O{�M)���9�o~2����Oen��ɲL�����L�&z�#y���P�qH��*�ԡ��T�4�eɕ|0*ɕf:Z$��[�*��*d�!X̎S&&5�(Y����V�qy5,��W�L6�̍2�@uC]Ŀ���Wl�P�h�T!�:�~�%����Q�cNI#Y�кI��2��2�s��hRNwS;��i
3xC)�������é�p��ia�r�;���_�2Rv�_�̀�r�<��2�Z�+w+V[�NH� 7[��<���	�(k%�ր�, 4�J���ϰ����5Г�����J�*�di[2'e��Xo�2�9 �� iT���8��2|�,���j�	������:�����먇�k�����̵I�\�ʢJ��|���;/�d	*;�QC�	C�i������}W4��:RyB�|;! B	G��+nzowC� 3[>�ۇ$�Ie��o�l��s�����?�-� ���g(�Ȩ���f��~����B�._O�th���u"�M�Çp'�=��
Bj!�+LZL��Bi\H��t+��+.}���C���C����(��|b�܄x�`02�+���*s5F�����ꪮ��P���ˍDK�R�UBVx�3�)ENN��z����鱅`�X3�K9j�����2���]�wzh�9���~ȃs�K����8�r�JAM�;��Q;�
$5�2۷������>n�B�g����a�hg%��%���o�#a��%�7��FC�`T��Rp�6e.X@��"��ڰG¶�3Z :�0���kr=9�
AkM�cB1�b�#��:)sQΌ�|�սQ��5�Mʆ��t5&�@Z�u=�]:|��7~;І�%�{�Fhp��+�g�8ތ�J�GV8\��EM$U��i� 
�����P$|��Un;^�^������{��+�c�Y�,�X/RF�\�=0� ��@Rػ6��s��Y�%9y�NG �~�0��r
���⪊k@I�nk=0N�N]֮ �b��v6�)%�Q3<����*b�^�����Y�}O[���G��a���
/^n�uK�Gޡ�������.�k�A�)ݘerU�f?g6�ڴ��� C[�P� t��m�~N6c��jʥ������$P',��Շ��Lk�I����M�0�%]~4'm�*�X\�t�Q#F/��*�h~	4�_����Y���g����~%'A�������U�`�`?A������ڤlr�^ ���%����U/��H��:��SP[왭o0�I�S�� 8\d���� 2o*űC�D M���(ٚvJ��h�;��An� �R�y�����6ʫ�[�ƆF1Q�c�#�nι��$��Qn�4K��� 8Hƌ��
Gf����gcw�A�t@
F�=Ԟ5�l�~Xf�����Ȁ1@E�Ahͬ	��u��yJiL����!��қX2M�������Wʟ.n��\j2�z�ˆ�Z�^�ҍU�!��Ul����g'/}T���(�ul���U��ט�sv�әkʿF(�j�9d�j-�k��ُ���dy&�m�p\�f�.:#�W�����m���A�S�8�_��}����$�R�:x��]%���E9t훫���a*p���&/�vS\�T��
���Af�q	;υܚ�)��*y��nF�bT<u��NmqE�.��胹YH`�RM����y�Ǭ��U�X[�+r���e�O(`��AJ�N��h|-/^+�':��.{��VN���&n��&��G�7(X��R�>H��S9�@�P������u�DL0�gz�v�j�#���p����{��yk�A~�2��厬j�7�aF'͜J��N�8��:�\��|Uᐕ��â�R��
̖N��ƕ�����~�*s�E��5�	�DO2�6W���">�!�}c���1ej,�Y������5��0̣* ���L�`�� �1�R#o2l̑0s*.&�Ϧ�Hdt���իZ�
�G(z��mzd9�g�u&)ԡ�1ߖ&���:_����p�]�Ԗ��)����q��B��(�ځ������/ �B:�� Z��6q�X�.>��\�r򐬥�y�w���Z=V�,��`_�����S�D���� ��VE6�=�K��0�y�b��Ú����Rϛ�/0E/�j�O�(���l�ճ?�	��6��.��~h?(#�G/���} �c�� "�D.���!&�P�����:*���K4�-�9Xd3�q�c��{�8��!�x�gߒӁOW�/dPH�(��/!8?A�f�?����J���@���h�S]6aj�tw��8�4:5�
���Yn�2�팆Y_��Cs���zQ�V?�O�s�3M��Uc����j�-X���oh�����X&FG>�Fj�)N��� ��.ŅD)x��Rt�sI��Eb@��ȯ�E�����Vl�#V�b��G`�^�|!���ϋԘw2�Y�r�(�VKg!�=

����C#0���b�S��q��|0�X�ȿ��⭎��^��ߊ��L����2�r״�U���3�D�.q!����1�fqdaw.v��D�<��U�?g���9t����׍�;?�8�=�J�M��b��6�<E�!���H-������c�	����b\L�=�]R�t4�
�L$E62�쓦�3�����3[�B��&_}���C�)Y f�þ��� �  �7�.�3����?��o�o|���x@�!�:�u.�LgZgO��ӯ��VC8&ԭ��͏)��P�c#[_%@\�{&�u+0G7���a+w�7����_����;£�>@��
�d��o��b���y"���� ��2m�*^W�E��)����ɑ�zޥϝsq�+S�*�u�"�o�h�+)�Z�x�B�qqǻU�f^l$���5��@�Hn��M���b��������8�-��e=ȵa�3̩����`���YF�:3�:�=x�R�p��,�`���#��p�[��S�LcG�}E��ly��&���.�5)F1qw�/��d�#aK!��K4�����1�T:�k�Bp��f�M���Nu'�AvClA��w����jϫ%��o�p�=�N��j��}P΀f\�:+��r(�Z�/��F�fh�t�u��ܺɋsB����c��U�[��-�o=�f���)! �!\<��_�UL-uwp����sx#8B��n�r�� �VQ�'k.�7g
��s�����_��EXn�Ts���y=D�]5�f���8�=fo��\����`^�ea��8dhJm{��>�6�-�\(�K�d�>�ϒ�ϲ���0��{�'�31��M��	�����=��P�4�g4j�r�|)�L�-�E#�����9]elk�Nj�q�*�E:(k��A?��|���˞�Es���E��P8�m�}��@�C\0Kz�����|i�v�mU�V �"���1t�	���w�Ʒ�������>��5L<�O4͗�x��'7�5�,�	����>r��; �.r}'��ͨ��}�s��%*J߬[�MT<<��?���dwD���3l���c�89�Ǎ��K���̓~~�'W|�\r lu��;�����P瀑�P6�h���F,x9?ꢾ���:�bO�Y���p����/7��cBrQ$]�Np'ob^�;���z�k���WnP�S!D�*�Ni]��+�[l�@ѷ.+�3Y��7���2^N�9
��|'���z_<P5�\qM��ŏ���\`�16o��8ׄ� ɼ.F�I�G��f���M�{����_�μ��흤��-AMذ�s�\�)ΒK��0tF/@bЃe�o��=*��N����N���o�뀳����r��A��@j	�2qe,�ޟqf(�l��Q�'�56����P�M���IA���6?�Gz� jl���#A\#G�����GX�!,
�G[ ���nҸ�	�7�C*)dR���ޏ��|A�+��ڨ����-Q�?�D�-_5�E�����^�Ovh��hx>3s$aD�vb>�ÈtÊ3����^Rax�,� <C~��M�8�6^z���>����-�%�������z��0��*���路 �`�Ȱ�R~���3e���xQ��|!:yR�",����iȃc>���*��y�+lط�u7�\<�2�tQ��;����ʂ�Fm@�f��]h0�{]7(D0�` ��u�ղr��)��H���M���j�9�\ls5�1��4櫺O[p��e&F`���aF#���e�6��:��9����c%0�m�������������]��~wr%�&O�P�[��G�!RpJ��D��և���9����)�T5a�����OzR� "Oe��1������
��
�W3x�^A���Ҥ��s����
�9-�yn�4�~Ϡc⬀��7KAD�4�r�|�ϴ0t��lC�?�dt
v�ܟnӒ��m�BrI��������8	"V�@Z���
�g�7�v7�����=���;��7������̡�}ᑛ��|�G����^��B��8O���9��Q��h�&�������Z��
���X.册���5̂.i�	�D[}�dݠR���+^~��	�*��=��?�����4^��H�=�׮���;r�j_%kw�L}�P9sG�mČ�TA������9�%����2�K;̬��Nju��w�L��'g>��a����0aOϓ�{�y��TZ��5
�J��Ș?�ɻ��P��Ui��/p�;"��ϰ6�vͩ�.f+2r�`�,�v��	 
�P�ҳ���q�o��*kW/��O�@���Z��-b�^���upu��� �:��T:+�E��*Zfg�q���C����*[�̜�1��/� �]��m�ꏚߒ��Bf�����·�:��C���I/�������%ơ����mޢ;N�~S9O�{�V\���I�@���ղ�9]ˀ"�kU3i�ˡP��L4�_�`��7S���V��������%eD�IFU�~<������OS��7VF�T���"�?�<QS��՚_!��E?�/a���`�3Y>�W�c���7F��B����,	��drPڪE�0�[6h
�n��f;�|Tu��_�e,}Qڻ����ͭŬ��x�����.,�����5sL��(w�}���{��j����J��7T�xŊiÁ��������� ��@��ET6��V�'6���lo��߶��=�u�[���0E@S7��`h�n�Ls�\�YB6��6܋�JsaLl��LӖ��ln�-F�Qz� �?�g�����늟� ��m��8�d.b��a�0��i�n���m���F*s)�d�v��/
�}{�]���Gޣ�mM��H%�X��5Pg	,I0��J�F�x��t���-�ZP�ꎪg��{q4z�|�����o����Z�^Ӭ�s��V�0;��s�.WN�b24e��!�c��e'��0�q���6��2�MY�Y�Iz�]T%>14`�̶�-z��I�<9�Y`�<���m=�>`���رg)�N��O^"�+��MpM��nJn��b�iZ��{�].�J]ſP�*Ӛ_�(��8T���=���V�m�Ԁt����/���2A�2&�A�^���T{�Q �%<�{�w�y�|�5l�XC<��Nt�o�ⳝ�g<OsFp�l<���*�@���܀7O�o���ϟ_��U��Ɉ����e�&��ߘ?^Z��3�)N�7��)�)���?dXt�&�jz#x���E+����*����xj��	��#�R��R�H��g౶�~���	
�u{�9b����ǎ�>E�P[k����	#Z墬��=�B��I\?����TP˺�����e�
���'�dp�.�V��i�`�6k\��5�:^�=�&N���|�B&���貒G�k�i�/襯7�R0h�\u���⪑���>&-G�����_WK�I�IBh��ќ�f�nK���9)n�����`դC�e|@$��k��l��k��!��vx�1�K�enO�K�ށ�Aԁ���Ɵ|7�������~n��X7\]oI>4�B�XݖW�7�4�XNə�[bG�!k|sT��ؔ,���K��제�N�0�/w^�tJ���d8�F� ���>�b�]�	��I��Т�����u��$����B`�������b�v+5G�%�!��J,w��+�D��Βu�s&9��c�"a5?����7��l���>�>d�� 3Ǯ���虦�9�K�~�&�<���W��V������-�f��2i��k���A��9���)2�̊)}�a���; �^;F�Sm�$���p�%)Ǹvc:y )�y~H�6�<)���<�f܉�]���Ĝ���8�)�G���ǌ_i/=]H1�6q����t����n��� w�4�D�fqS��Ե�t�REID����^G��`�k��S	�^U�\XA�>��e6n��uY�T�� �X�	a�M��O��:�(Ek� W�k��eE�'V�S��)��lg��^��4��|�Tq�ͼ�d�,����h�Z���c�:���g~��^�kiU��AQDxE����#ة[��jd��[y�J�
����3�1;�ћխ
�.�mf�ͩ�k��owJ��
x_���d��[�8�Hp3u@��m���4�9ZW�V��b�I �����vW�p�W~�\�\Ԑ�޵�Q�P��P����0���#�����‍�s`��c�@8<ǑF�݉��u�����ë������zhma��/��V:pEɑ��@,��
��ུ�)�IV#<����=$�
��ڜ���'8aZT��T(`R���f����}��O��ݢuTh7����Dw�<*$��G��t�*oXp<�e<\�E��(����֨	y���{����%ݰq��J�O�6�"��P��Y@�D����P*k��R��<�����Ruq�����I�'�n�&/����9�"�*�Dƪ`Xp����ԑ�[y�Q;��	 s]��]V�'�ȧ�RF�� �@!���0:��B��1��Eih�{����>�F�;����ȩ��~t�i������~��:q�1(u;j|�~7��"�������w�&{�Y������Ʊ	�ְ�Щ����q��&3�,z�rA��݀X:ȃgE�J�u�*g�(ŠM��͉a(�_D�F��~�Uo�(8f?�����|�3z7̫#=ԃ8 a.h�O�o�@����,Ƥ�MY�S(���4�2ໆ�+	C!��-��EG4 �C	Y�.bt���3�]P�'��\0�̮K�--�AdS�mի��� W�ZyF��,�n�����e�������I�N��h%����q�J\�hK�O����20����Y3��h�q[�Ӂ+��b��v���q$�i���Ω*[p`.��+��ϟ�h��"P�1��0���62l!��]�^{�^����ܿ���P:K۵@��Zv���NɅ�	��Q�	�+效��n���k��n�'J�'N��6z��{#�^�~�M~&�%�o	L�N�̴(�#�[/��B��`J|L��'4}�Fm��7��9�7v����\>�Kp�m��c� �.Ԟ�K�J��f��Ģ�@�Jae��{�2q�h�=���G�D��e��^y�
WV=5pG��7t2��t��Y�hY�Ub�Զ[V.�����*ƙGP�~�2���[��n����X���������3`�t_�&�����x<3O*{m%���>�S��	�N �3�#��n�$�׆��_w�iQ�1�,��/#Oi��Z�}%�Պ�}B��T6�<Qm)�^�kbo��C�94�r����1l,
��:mq�=F�Do�K��Ls���j1b4�YM�ԅipa��F�8&_��������TU��#<�X���� 6���	�[�% ���$H�ylR�&��#f7N����ȌY�������~���k5b���G �����UC{�=�Uҧ�v��@>SQ�s*]'�~Lw3����N�Ei	Ti���`�l�Lg�"�H���L�u��k&Ɵ�v��T# bx-\�4z�Z"@���E���2��	'��	O�̴}� ND��{A	,��|i�4�W&j�޸��
�5��m��oЎ����)���y�R`1�#޸!{�?"s�4Z�{�HxC��ی��aA&�Ϸ"D�J�I��A��,ؾ� �(v��������/h�������uy�wT�y{�4T�t�Ao`�1�s�x�����.�t�Y�	� �a���$u�2M.���J7<4���w���@�����ݕ$���T�J8QU����$�b
Z��U���z*bFx뉅���w��ai�Z�m�V�*��l��ڙ���v��HnQlwW!��)JLu���)���
E�\=�����1�������Q6^A���}�D�>�4�Ʋ�����3���c��Ħ������B����x,��F�y���\A�)j~��#i�nà�=�.���RS��*ȋ�,��mV3�V�~`-p��: A�\��&�(t���򸋠��2D�t}���\�:��Zu�Yi�<�����[����wXY>xnE������4�ҫ�K��u����¼
�7�KMBxVG�P����8V@H� T����ڧ"����җ�N}���OZ���W���=�_��&Oli�&HQwǊ���nF%���I�ei҄��B�|�8�u�����~[|��J��o��IxT�~?\�fi9��1d�($-i��z�l�O߇8PD��q�����PL�8�
���R�^āyB�6���r��O��n(C`��1@�Id�N�SX�`�U�g~�~�T�+w�l�Q�i���粁�=&�Mo��O���\S���-���hf���*��(�Co6�Lf����j���R͹�4|���D�-,\�e'�ޅ�4�gVMɉ�+Yj��}Z�$ȷ����庵r��q�M ͺ����D���;���@c�h��?Ђ���L�Z�_��
pS��o�!�j�i%�z��Kq+�8�)W���}�؆�$�2�r�8g_����Q����X�����(����u��F\T��Jc�cG1�#[؟9.��`���W�Ùw�t�^�3J�)}���b/@�(�����
���� ���9�(s��x���Zc�O4p
�*�G6%K�K��rT�/�3%P_�*�:r[-/��l�Ih��FTNb�43�\��|q]ꢗUܣ��y�C��#X0�BI����#�t�J�U�H�>/ߝV�d"5���bD��x�"tǔ���YM�z �1�hі֔hE'�0m���L`l��N_�׃;s���,WM,$�xL�Y��րi},mN���w�;�=�և�D��]���!�����oR
��p{_�Cn1�*���ճf���{�%Q�F�p�?�=�e���v�'��&������QTЭ��:x�Ti^h2��ز�x�CB���T��#�BBtSk��E}k�z5�7��Q��|�ŷ X�Di��H���jL��9q��D�c�_{3c��Lo��|6(�U�h'��~BN묫x��E�eSA�|�rם���!$i��ʿ�>�P�V�X��.p^r�v����(fZ�p�-��kUgc���ڷ���i��M���ro6�~̆+C��jHPwCR�ɝKbt:�Q\��T@�/�g���&@&�r̵y�����)}�u���$�:RP{��B�^9K6������G���c��6crV5o_�J��Jy�J���@j�T�a�"�e�s��"��,�,��!���F�u���+��j��a�E�K|�@NIH!U��_�,�r4�1ψ~�$������6�5���R+q�R��1=�𴼲!����������ն,C�<�'c&�����+����=���.�:����X:��R`5$0  ���]?�YU�On�9l�V���fʊ�¿�������@��-��#˴�of�E#����g�A�v��8}�ר�i�-�Be�ѫ{;�9�>�}_�`�Az�&u�0�<پwd��AGKJ:���o���+� �sL���LS{ޙ~~?�6XUg@J�`�G.1�<�?B/�秊B�C��3��"�E�3�o��ܷ��>��<p�'O~ۉ3�ˌ T�B���}�c�_�h��b�&��E��j������w��|�Z����?o���������C�4����oj��_�Dk��*�|O��ƆU��Q��@�~�PXyNli���-
��c��<)�v9�O��bݯ�G`�<'6��B�]�eA�9.h���T�N$�{J���y��F �Y@�Z&4�0�R�?�^�;��1B�D�*r�.d��`��"V��fӿ��hP��o�J�c=������JZ
i���g�\W�)4"�/x:O=�2��f��2����F�i��s,��p�=�g�j�(J��%�;O��{��k��.{��.��A�Dn>��F�5���)7d������c�����l������l��Iˇpd~���4��<�X7ia �7��q��!���3���R�E|��K��i��a��*~�Vp^AObe�P"!�!�qrDR��f��@C�;"x���Qa�+xUf1�U��D�h�}�*�lg@i*P	~����A��p+�D�@�6�ی��~�65�AQ�f 4���QC�B�2��QRZ���W��1�(�__9�Gp����(�����SI��]�x
�Z�6P����8�RT�-�!�1��P�y������Թ|xῘ��m��"��e3��u�}��a��N:OnSU\g�ƺ���\ G�n�TGXkYz�9�(_��l��~������+�z�����Gu������}T$+7�}?�����rW��WFx�مTUr���1j`O��f�;;N��	�{v�_p"�U�Ӗ������5Pv��\>��lˬ���=֜B��Ț�G>�������k�ہ���E��7 K�������4��5=:�4��5S����& ���2"w=%$��s���%T�F�N��Z�{�i�S\�P��%Ē�m�2#���
W#+|��w�~i?�})�F�E^���9�!6M�@&�����_xR`z�E�]#������� c|#O�{��њ��Y�|����_Y��G\�:�N��2�p�ei��j�z��d:_bėi�X4��	W��2[0���\!�I|����K\�@ �i��M�)���z�jn*��aմ9#X^��\H���y��O����TD�S�M�y��,Jr6J3i�i�=i�@���gfT��L�Q����ѣ��j�0�,�ϼ�үq Q��烳u�
�q�3o�i�yⱝ0F��yV���.iZz\���5�Н�.�x1��6�I�N�t��+n�8J��dsT�򏡟)�������\�.$@�Id�O-ϋ�|	1?�]Xx���?�6� ���08�a�	'���t'�653]4�58�ՠxSe��^펂4�Z��N��*����¼>����e_M�E�Y��rYD2y�#juk4�kr���|}k&X� ��~��L��78뱿ւ��
T_oqH�8�B%*�؜��}RHdξ����B����դ_ؓnB̬uk� �	��8�Mګ�Z�j썅����P��:��i>���Po	�,�&�pD
��a:�G�z,�A*�A�Q�v!�_Ҝџ[��:G#C?��aڜI���'!2�%��L)�L�J�'D)0�̨I��mj���7�n�*�E����0}�/f��Z3"����
��������ag������	c�$~Xz\4f���u71��Vմ��?:]D���WD}O��ݍ��j�Z�g���N��r�>;cs���+��=�HڭٰqqGD
�oR�-�mN(�$�ѱ1J�������ܻ�?#�T��+��>��,�Y[-ZMHH�lfK��'�\���a�e���s����{�͟��&oO:y��}��n�$�+p�xH(����wԌ���	r����M҇�=�����@u?~�v1��={�sz�/+�(� ��*_�	y4������<�ǿV�6�I_���V�8�9Ss��3"Q�f�4��:��f���­o���E&ajiG	���l���;ꎵ[<{�ѣ���J&��B����Et��~�VA��5�<��t޾i4���/i�d�_u&��=��|�w�&����
���V��A�(Si�~hq-1+�_A�+�ݻ6'����Yb���^�1b9����a�9�$�=~)���=�ω�I2�!�հD�	�=�.b��L͉�p���u	p�����A�X�#@��Ö�-O�`I^�<>>ދ��:�`5��:���E���c3���v�Bi�#�Bڙf ��Ҵ����壈��L��`_�"�5���7�?o����_<8�(k^S�o�g9U��{��Ag$�&=�`��#(ŧ��Wz�=�̹U,|#Q#��&F<8v��HG9�H|�����J�
�(�؟F<##�^�:g�6�<�Q���Q�@���i(�1!���Ny���u/��W6�O;�<�Q-`�l��h�5��r�.�|��[���#�x��HJSOUӽ�?;S$�=��X�/�g��(*s;�5:�݊���I�j�B3�'��F�Ī���.�H�(����u��W���#��L���	�)r�(����!d�����j�ql$�C��Kx m����(�H��0�I9k>�\%�T�\���W��`�sj�>1������aةf�[)G)��9����#k�
���A}�]����WSBG/�}�� ��1aE�>*�췋P�� m��F��7�z�`�$�̆��)#j�gh�Œ����c{E
aw9{*H���|��\X�eG��V�r
:p^���T��X+3��3�����n�/i��߷��QSddaF�7uLo��� C����-��!s��K(�������u�W��F%'G(������%V�p���ܮPo��Xd��$�7M#���;iV������_}��X��`�)������o��|��L��Q# [��'_ ����f�\0�����<)�F@��5z}��O�����%9LԹ}؍ط��i,/ۑ�G������#.���V۽d���ε6�{��L��D,��EG�P�2T1��`>i�~#�޲����3t�ԁ��79E����ʍ ��g���ȡ����������skEqT۟�`b2��_&	�~�k�F
��)i��n�G��\2�?�_�pk��ir&��Sl�ہ�2����8ю	�ܧI�f�P`}