��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��5���5dδ���KdXyݕ�2�j����B�}��AlU=w��m�C�}�S�[U ���c��6��u�������K���ֵZ$�<���?�ޒO 	��ȿk�Ƽ�o���n� �����4D�������;����l�{6d�0
�Z�^�^�2�;�D�
�UjR!�1�2>��Lb�`�D�l�W�?��9�J�ס�Y�u�kK$�ɓ�#�NA��Y�o�~8g�!'Q�Qd���1��+j�i��|Dσ:���x4����j���g��6��� n�벙s���c� v�f�GMcˎ�����0���6�R��$́r���E�^vq8g�O�jl\	��ч9ݢ���/�p-Zo;i�c�at��zb��M�պ@
�G{���CM��0Gm��w3���Q��ɛr�v�^7�<��cq��Z{ۙ��]l���gw��Eh��v|ۻ��&�xN�I��X�eъ�_�PB ��'%xRWh���e}��w��X�ə*J�Q7�j+#�1Q"���E/n3L�r�~��(>�,^�"O <r�b�?��cN2}�8��[�sA����+k2��\�8�YҐ	��~��@�D@�|��u	T�IU���|L��Ms���<��ˊ��U��F�5КkvП=5Ǩ���-�a���ow���I�@нr���\��.C��JxNV��IO�,�{�F�\��kR�[$t�c[��ܘ:^�� ߐ5��nV��m�H�p�m�:��y!o�k*y��P����P��U
���܂��BQ���,�O�/a������2B��1�f��oĜe7�拙���{� &���"�G1����E0Ja�>��񻺼�\�z�aA�=a��2Oq��VG��6�H���c�1��`^��uKr��Q�p�Fj>�ZJ.�~�:�4F�eV7�^�q��M5V�-���9�V6[Ev>��^X'��$9ҏykyerW?r�`�7Uy�$����G!�Y�M�}�J,�ރ��;2�Gm�p`s�fH�QC��b�jÇHE=yU�]��#�� pHbƛ��ӱ}�r|��B�z�=���iu��b�ͬ�A��3�G�j����Ɔ-CmR~5��5:muJGҷ캙]yx�:��g�B_Z�FT�ba�<�}�F���[������` sY62��R����b.�6}�����ͻ����D�e>?��rј��@+��2oñ������'�� ӕ�x�.�\}5j����\gA���<g�1�%#\>��T��С�I�A
zgI.{�.&��0�9��D@��5P�����	������R$tM�Bb�vd��b�ޜ����K7Ƙ�&�.�-/	v1(�r�\�G^9������ce�!���O\G��𳈎��W�@e��+��m�N�/�(�.�d����՜Y�3���R��w�2ʼ������R.��N�^@���ي )�Y���C��Tje���`B��%X��V�����i�b�3�.V¯	�w��i��O���K����u.�Ǫ)o�]-a�����R֎#R���\��'���~��hoЯoH�e�!���w����TZ� +W�O�6��%���&����$�P��2+[�ie�l�`Ni�Fz�OX�S��	D�W�����G�b�r��S�s0�{#�'��C�9�^�k�+�C)c�ߟX��2�9�-��4�/�X��z1&�t�m�P�}�]���Y[�0c�-���;�^beu�]/���mH�(́���ွgB�YY���\^�,�/���rb�|�<�*-�2��r-�/�խ�(��^���*�{>�o}&�H�����_t�r��5R��Г�"�O���^*m�"U5�yF<���
��
.���
Z�����^��Yb�ZՈ��5�î�8�o)7�!����*Ggya!�hſٗ���u�㺎��bRK�JLE(��;�O�bORNۉ��������R� �A��i�/Ky�Q�hVb�����]8��a7c��J{%�*����m���&����Z.�H+*}s��#Hd�^�>|��{��O* CG�R���a��_DΉ�)d�2�W/��S{�*���Y��q�J@$�r�v�oG�
�V.�5O�2�9���vcg�7z��ˬ1��߸��Xi�� ��3W��7�^#�K�d�W��nOP��<��PB����ʀ%�"���s��m���b��g�e�F�q�4=Q���o�(3\*�;�~�2�sP~7 i��O�f���]�OVi�호����5���T�X��R]��@�#�P�؞��F�`c�.|�g�f<��!�����\[r�-}�.���&��^t
��q�w�����<&�Μ�NE����NE W^r�Yl�}f�~\��<kēb�5!w�7d�n�C4S���,��m���.� hob�T :�*n�<����hi������)�|Ӊt�]�Y�L� z���I
]�OF��J������ߒyC��c�pm8��a�����{�	 %əw'�ߓ�e��D�)�"��#��v��fȩ �gaR�)?�@�o��_���?}+�!&3���ޏ̝S�v�N��.�F"K�cP����`>:~���K�|��I��^���z��4j��)�����8��~��p��+p\�����'��"-�pZ~�@>���K�"�4�s�����U�Fg!�r�����t�T�Ӯ���uł�Th�aXe��!N���lY�r4n�u�Y��dFsY�$;��Q��8"��Ҡ�����n�&�F>�0�Z zh�OD
��WD��Z��!�Ż�N�QֲLC_<��}P�m9����T�cT&V�!�ݰ<
��o ���&6�3ᯮ��w2�'���'��&��g�����#qz�d֭D���1B��t�x�n㊱�q�56���%7�M��^��O&L��e�OuE���Hn^?���6�� Y3��23��X
L�Gja��-2�W������P|?�2�?�򋠲�g�����U��{b-ndB�	;