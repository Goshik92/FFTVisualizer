��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ;l�Fv1�Lژ�O���3��������F����Q?���b�V����Ţ� K��Q�G�D��i�o�Yʫ�|�F�V{:�� �{��LBB���Z��^sӽy/��[����I����k���'_hx\�Ƥ�?���ƫC8�r��j���?�[�b��Gk����s��$E�C���Iv{��Ϗ.��R+!9u@Gf6�e+~�7k>�_3�T�@�@����58fW�o$�T�h,|���z.yhb+�[��>���W��Oѹ/t7y����8�A?X�Xw��J~���k.W�$�'��(��ꉑ'[J��TF�S���o�z󷬓�I�UW���{�|�M�a���@�F�J�Q�tx�tEV��Z��i��lzt����#��I ������T0�=C��'1#"V,���)�r����4p1����Ɠ��LS�d�,BbD�י��)�@/
X����0�9�C�'�8�5��I��*���ŀ�К�;R�g2�9B}������Qj����F�5#,VF5~z�wY@�g�ږ���jbY'��&W���Q��p�>��@牣@N�#���Up��]���ߏ����\c0�4i���jK�tƩ�H-c�����d�@+�FRxY�,��~F��(��y���^�)P݈�k4<�w���Z���?4���E�}��_�á��š�0ޜz/B��Ѽ��#f�݌$��3��z#G �W�fĨ��H+hnؐ�&�,�Ɍ��9�ċ1�(ֱ�{��v�RF�T5r�����F6�}6��2l����Ɯ-pw@���
�O1���3��~1��І6	��v�A���@�e!����� S-����193��n���2aD��T�=��yR�z-y(_ �>�	#~5-�_O?$b��t�;ݵH#h`�V{Y�:>Y����:����U�va.�O�M��?��(`�+���=}ӵU:M�k%.9Jn�ۇ�m� U�y�RUK{.��xf���¨��yb���2��\�;|�~й9�\�y��3��A��S[3M����S(�/ވ�=���ז�xLF�a����G�
�����W����~�xóX�p��S#)壯��E�V9�������u�&�ջ��'0�~h�E&k@o�毆2q���G��`3�14��9/l���P)�Z�$5�b!�_o�q�sw���'��,8�2".�,:(�{D��:o����5H�t���VF��Y7j�l��� ���3�Z����/��r�6%f�
�>cPri�Vr��lДD�<8� �*���*y�<���e��]�b0���8}z*/���F������Ui��J~�7\5��n��V���4�k�D���ԓ��H5�8���U�5��9/�&� �n���Hu~���94Ȭ �����Od��"W�6��s�Ȟ����ADO>*���8[�ޙ��mY�y��`�ō�а�z����iUJc�=Q����p.7��aKg�d�i��u�)8d����?H���dT'��������!���^U��<�� g��_�Z��tz�ĝtI!lA��>I�|���E��J?�sBC��!�Lr���Du���Hw	�����e1#7Kka�2
s����IʿOԆǚ��6�g���lה�>��e�h*R�Fp7����3w�[�.��aX͟s�!d�����/�|<A~��Tl+�f"ծ��0�OP�7Z �C,�mO��q=5ָ�jI��l�L�Jq{�3�A=�W(��Â�D��� c�΃}NL�ӷ�6�0-��oR˯��Ez~aG���|fI䙤������Mj.�|n��� �i;���uq�P��@��au�iY�߸��+��Ǟrc�ۘ�%/��9��_��C �d������!P��l�?Se������q�M��v��M=vk��0�������v�5ݏ��\#���Oc耵���FA4�;��q��|�+
)�%6@�E����Ԧ�2Z��J��x�EGdPρ�����ҠZau�ߟ\M�!�����CKj�k��*YM\ 5��Q:İ>k3R-5;����uH��M�ttn,�`�_�N�b��9�7�|R�	t�k�������xqb�5Q�r�]�X[�����2A6M�8���9b