��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,G��U�	�oJZ�@�z�����>*Q�p��~!}8~��m��sDmN��3\��\�A,��y��,�y'Zs9|�v�G��Z��J;����`��"��t�������UnRt��8WP�Z#+ϙ���\���~��/M���jы�IFA�΄�Mw$�c*A�ǉcS{�=I��{�Wj���O�5�����5`�^��Io��J�&�?���Z��|>�I��ߨ�
;�,��TJ�'�S܌��V�� L����6��2���3g�����D��d�kޱ�LɲюEb�^/��G�>N4g�ˋuU[W	�+!UDp��
��%$shp=^�3����]Gj��;W�\)��͍K��>�-3W��8�10t��~='%8��%*���(�Ci�����Ld��+T��tX؃��?Z�S~jZ����ތ�{����)��d������i#�S���<V�v>0y��:3��GT�	c^��@dp`G����XY���{"AL����B��Zla`�'ût�>]u%V������~rjL�Q&�	h@S%�eI���ƙԆH3z��(3����TEXIw{ !��8��N.�?��h�vB���8���}�9�y&�
�HT	x�J��Ο�o�  4}�N��,�����pY��Y�V+����WM�%,7 E$�L����ʀ$TQ� �_�2�V6x�P�w¡���B��ql��V����?���Ͳ����ȸ��h/�q�,��P�ˢ���%��d�wO��2�c5���@SE�6q3y,���ю��f�Oۃ1���"� 	'��q4��D�qsF?��=�K&�Ž�O���ȵl3ż�-O��:�z|�.�PxO�\J>����ښ�������i�6o��>er�-��&`��5��QK\�V9�&6�]�8��H�U��?v��g%��-�� V�n�P����>y}M���LEQ� p#��?ٷ���;ga.-���@Im�pi�<Ѫ/]:�ti�dH���$K���u�e��nd�چ2�-��̝|�=S��~���;Lz�/�J�l��~X������1�	��?~i'����z PjS.��T�Y���MS�h�������ȃ�9���`=�!^3�m�&�$xe���I�r%{m�rN!c�5��>���5�tI�m�e�m1�����l
<4���;�-��1h�~>-�ߩepR8�<G<�L�5c$�АE)� ��H�d��t*Z�g�]�w�i��r�Ɋ�.�r��q��(����?�^�1��U3��� G�\�����!*��g�"��b�Kw�:��
ĥ3k&I� �k�����a�OO?���9�]h��,�k���ʓ�7��"��5��������}��zH�<Q�����2�����/�Y�����x� �S1�ajt�{-��܌HD@G&�\�~��Z�ն�;�n��=��J=�z���yC�^�m��q�m�ZvV�.������~pj�"f��Y*3���Z=��/�$�`��,������ɿ�:�VnĘ �=8�U�+֚�K��&�-$k��G�����)Ԭ�4{��� N�F�*����!�=��J�C�W>�֥�8|Ɍ�Vj�Bڋ�>6�j���z��ݷݾ���KL-�D�ty�Y��=  ���y�_����X5��h�	 ��}j��?�z� n54��=�9�����)�J��c��l��Q���E������v#��V��]M����n��	��LXm���E*޷ɝ{	��lC�ν�6�_��Z/lj�X;vcT�X���tZ)�_'�\\^0�:�k��Ƚ��E#���=�����[�F<���<��:pһ���d�X�FȞ�U�tb?@o�`"��:�w�p�ۨ��"��+����dB�Ĝ8�����ѵ�GA�?���@P�kU<c{��.5��!j�X�Po�/�N�gLL�rF]�-��egXęR�������ϡ+"6�M$�t2�gD�,���0�9��N���v�����j��뷎w<["���x4l_�~��$�m��w�Q�{r�}Fsk�*�#��������e�����st��[���l�^����.W$�����ς�l�1��:�p�o}M`�``�I��
~Qr��z߮�^�5é�m��H|K{����N�.��S��yɱQV\t�u۲��l0��s�1���0f$�E|�H�|B����7�i`��Dl݌��C	���x_�IIF� 4����EkW]v��D=���̫�λ@��r��+4���O����7�i�3�?���I)�}�^���Foz���d��(8A�錒b$��#|�\��O|9�D[�}f?��r�(of��2��|�f9����;6�����ߞ��T�fv�6�>n�d%w8�M�a7-I^O��nr�n�z�,�?��j������1i�xg'"���i����ߊ��^�ƈ��x��_~�c��V�G�72��JwWX~G�`�ۢ�Ϙ�;�aתݍ���N�,=��~�O�߲LA�����C��ǅ���B��]1�!�ųi4�N�t��͗�$O� �o��b�)I<..���NjƝצ��x��bC���f�����+L�!dP�
����=D"�a��S��!�f����+e��l�sE:����Ѱe��Cs�.>{�W zp�&�z��{�������R^���f���t����c��<,�ӈ�#*� ��x:l��m)��;�v��x�6�JB`����[�x%�K-雴�Y�%�9�$*J� Z��Orc��� y����<h�8Eu����b�[�@�$}!���*�7�� Q>��M���J�Us��An�8K`*��pޭh�*���މ'Y�l.����q_B�DY�/H�R�KVD�k��a�P�;4{�>��_Ly��0^���U��}�PH��w*��m �Y�3�a3ԜX�V��k;/�cEC�l��p�MEg��_&�M�C@��"����^>�
�A�>4����P��fЁ#��X"E�:е=��&{:ʌN���6I�x�ߺ!kvm�^�Sl/c-�_�_M����1�zӈ�|��[[NZ�
N뾴��称���kT�QLF�K�li()G�CT�7��gw�xrL�So�$����v��(M^�����t!�q��p���i�-�i��pm�2�֍m��7�ʱ��pY�[�uXyd����)Ɉ�b�Uu
�zq�Z����ʐ��||�����L~d:=d�}����NR�����!�o[T">�y�T�����l��.���"�:g���_�r��K�KW�^-f7��<p�y"8�j��#E^.e�Kw�4��	�����ME��A��տ<����>+9;S״E@.Ȭ5���,�0��QDY��%M�H[�E�B�4\l��!V�tU72�[� �,�&Hx*Cr+��������M�G�)� ӓRpP}k�p�: ��|�����6�c�EWؒ�'���҄gA
���k�E4w{P���S��`�,w#Y��iI9��q��[,�D.�:����:hCE%�.{��*��׺��<������;������ڨr�'}Ğ���k�Y�~`#'�-�+fͅU���r�N�TdKf�]���e3"@퇠8�a����h�W����忊�0�c�*x�hbI9n���
�jO�3�*pykY�p����@��I�=���hU���<���G-�>��1�����R??��z�SG�3���w� ���-ܳ!k[��y>_�0��tk���st��#�<q���u�~|<��[R)����N��'G�$��ק��"�nl��3kd�=�Q�RW&{?��p�}CE�Bf���=X't�n;C�Pl�&5�O�>ův����O�����:q�̺��sl�V�}�JK�4E�!JBW����;<棼��vH���NZk���0x!�Bҽ��'q��Mp8T��,���I	3�;�^K9���1�i�@�~{o�Q$53?*���e�+v����Z�`M��۟�[�J�Z,�n��n���L�}�����3x��c��"d��l��N���l_򚾎`-w��L-_���Z�����xw��Y�5�筏��y��,!(���l=�(��a��o'CH�!Bj�fP�͙�ڼ��΅��n��f�[����m��7%���f߉�~r)�l�B�1�2#�jE�:%S��n��������BY��Ɇ����`�!ʞ�8EMcո�`�|
^�]�ݔ�>�bق�f��M����X.%�x'���T�VΡ��
�b��[U��8����T+����`_����j܊[b��`��\�m��#$��+���c:Т5&[/��uqM�e�Z��@:�6��ɒ�,E�-�l�l*8�:�������ۭq�bO�i���H!�xףe�Kcᤕ���뙅F�z��|�����RW?đ� ���4~e>������,�]����L|!ǋᰚD�Ѿ�"Ez ��CO����9��0]��
[�^��a����$:WZO���Cj���ʨ�)>m+�AOq���g�~Q֑��78s�	u"�� �0ۈP��a$���5z@T��1�=ܬ
-����F���lyc �&�yd�É��|I�P���f:4R͋���ŋ�Ց��nj�U��9Ӧf J��v�y0k:t�F\�>��Ao���Ca/��W��[�v� ���ڡ�&}>�?C�~|��(�V��J:Ӈ�S�W� ^^ND��k	�˅� �*�AQ�v2�M�ԨD�Y��'�e��.���-sx�V�8 W��^�p���)]�s:�7��(];."�����ȠԲ�m~4��Д�0
z�."ZI�1��(�x� r��Y�u4?0c�K�N��yV5��z�e�һ3���DBD�X��R�)��v��9ق�?ѓޘ�$w��7^"1��a�	M��Z�le�����O�O'w��\g�q�1��5O������ϛ���ܭZz�]���e0��ؾ�[p_{¿0���/�+|���z�%nِX�Ry����vz��m��.� C�������e]��Y ��� h>�X����%������	�B��h0F_���yM�͛����>��#���8<,)ٽdYZ,V~0n����H(΅J ��r�����G���U��Z����È���l�e>�5��؎��S
�*fn�x@:p��[Hyn�LuT�D��G	��ʛ|�P���[:h�M��P�<{�0�����)]y]�&� �f�2]ߢ'��`o����	�Up�}Z�_D�[kb�x=%3�e��i&��^�d��KZ��LS`Fɖ\��	�Pn�r9UU��I�uK7�T�+�����q���(��İ�ԋ �z�N�G[�!sԗT�f(�,;U/�1�_�bv�T�:��0�YM�w �MfrѤ5�q˔@T) G�E�d����V����j'.�y�S'Ϣl�H� ��풫�!VM� �#Y|M��L�Hs�]�<g)�Xc�hbJ���6>s��+���%Q�ͼ�$�a����ٟ�ד+?q4<�M���ЬT�z�*�|�% 9���u�JD������g<g9�k�t;�%|�R����pov�fC�q���*�+�s����Nf�\#��~�j��K�ؾ�/i��F�A3UOv��<�jU�kpLGE%�L���3z%?��g�׿~R*����l��^�EK<��c��o�g&\,~˾��п1,�}�GT1��0c��!U��n�j�u������I�{����)P
�h �]ڿn��p`ެf��Qtx��9���4�:j
���J;�q4>;��?s��,5E�iA<�q������J[�B8z1]q��^=ͦ�	<8v4�5�ڌ��\̡���J�GF�(ջw��8�$��$�Ĺu��D��:e��w�	�D��f��.Ze[��n��3m�|n',d@�ađ;^c�18J5 �kϜ��/?�WY/kˍ	�1X`�4�I�Z�wQ[i�v���	��pk�3�7p����لh�Ԡj�'Y	޾vs��Vm*��&$}�6-�	�����.�4/�Z-�dt����]֎��Jpĩ��*�Pvaƭ��W0Zl�d�]�0� U�| i�[O>�D'7�n�6�m�U%��N��B���D�a�պ�[pf1�z��qz� -w%?������o�}Ŏ!;�^�!Z��J.V$��ی;�m�������noO���H��l�y�&)��*��pP�^�y)�P��7��%{�i M$^.s���eU�������cm{�Q.���L#_/߈��`�*�@�������c"��*W�[:āri���6��x��n�C���A����d��T/�-p��ΓC�F�sVzu��؇t��N��9��>\	�9�g�V�IdK�Kv��Q"ȼ0�:Q���;lR��,/YS���sKXN|�A��g����=S��I˯-A