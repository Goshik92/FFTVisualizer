��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn반lŔޢ�H�d��qՠ��I�/{�a-�l�b�����)��!v���?tG�����#�g�/�@*�Aw:Gʭj�wuU��1��[�iu�_%�9o�*O$��9'3��=,�����pz5f	�mw���*(>d5%��GV�u��ݚ���s����9�"x�hs���-M1��Õ��=��ޣDʈBM
3�/Ŀ�iCB�|QD��{X
(9z@��`'/2����Bt
2���t#+'8�`��k+B�S2Pm^��1�����S��jk:oC�ti��[��浝pc���<�$�J ���Yq^��i:��W�@����UY�x���uL �j	����'���X'4������ �R �/N�K�c��_�ß�ϧ�{�c'���gS�p���aU���(�IR'uv�YA����{p�Pɖ�Rp�e(c_��=���BIe������P�ғ~Nun�FM  �~�
��ǋ��_�cӜ�%��s��M��W",QJ� 
�R�\�7THBs�j����q,	�6�o��`��pO'���[n
�%�������l��Si�1�GJ)����,��Frn��%�����-��?ʂ��ŝi�'/�$:P�qPH�2��L=�3�[ft�1�Gu�vB�N�j������}�U��qф�N嬓��V�
��m^��-�)��))��Z�L�x�'묔���M�O?dfN��nO�ĭ(�,bܳC�faӭ6�}�e���BŝwK�0�;i��	4�oi3T	����H����Ւ�y^W'D��%L_��M)��>�`�dq��1������}�>j�jz^�T�a�aM���EH��Ӹ_��B���h,a}+o�x���Ik	���A���b�K�]G�x&�+���5I`P�2������w��ê���;�N������%�S}���
��>���;^|	��^���]~	��C0���7���=&����7!�T��oS�5'�H�"t������~5��IE�%k;�AW"g����.�P��Up�1�ǋ\����Ga��n^��@
R��@˝"K���_��>y�i�4��.mk/�ݒ�>*�ډ�g���L�3����Q�k($G9��>J����n�˚��:�46���D�%��=U'C6���\a/�߮��c�؅�C8�f�s����V��1�1x�q��ʘ���M��I}���KI�<�5e�du�4
�a欇$�u��凬��%��N�ڒ�pD��$}�՚.U�hQ�����V�ьN��j88<�t:$]e3��͈����?���ҨN�@ʤx��g��{'��jџ.� ���4�������؍HB�!��`󱮟m�5����U��~<�L���ក�9�9��c��F�9n�\��_u��"�A����a%7&1��qDj��1-c�q�Ifj"U��@m�z�����2��M%�̝Hk���ϱIM�0�C����O�h~}��s��(?�.Ʊ} ��[�$S�
m�)~��\�t!��m�-)]�7z2/0�
��z�"^G�P7eՖ��wbG}���)���:���TFO=;�{��#��x�˓�rN3n)w�?����,F��r�߾���Q	p#�'�F��^�5:�����R���c��Q:N3�+�$��+p�SV\�'&tЬ���1�Q�^)�*��z<�Eյ#�)T�����.#vL-t����V����f������Z9��T�6����/�vYU�Az�9ѓ�<|�
%q3�aU��â"��%1l���s����wH:-��Lpu�	�5;��靊Wq8Rx��TK�ӳ����F�L'&�,)Dj<�jo�J���7��׃�ɻ������m�!k7�)���솩�t��'B��!`d��(B�`ݭ�KN�J ��udRߵ�����3&����]t�)�h�����8�b���R�C.u�r	V�!�f6-�|pˡ�!�k�-�hxA��Q呎�q�����tgs?�S�$M�j�[@����5�8c�B�+�33�Qv�0�{�V
?޷���ы)���h�+��7����P�D�g�"Jəo����
N�����#�X��Q�䠐�1�#�Ug�Vb���G(����t�֋v�e��SN�-�^��-A�0\�<��n΃Xg1���QdkZY�p���H2�na���q��TO��s�I��B�
L����Η*��,[3 5�����x}��\�ia���#��1(�Y1��������c/V�m�D��r��r(�c2�ڢP*�����3��g!n�'E�P��V�A�O%����:�J�{�0:]Ӈ�U7g�A�gF�\b��`���@�K���L��C�b0~��k��L�����;UG��MU�/&���ʚ2c�z3~RuF�d�:�ނ~3̍���ֵ�L`��m�?d^1f���x&�2������%���?�"n�??�ol-������R���Y)oIG?T쥤K�*	�4t�^t��X�)�点��g'��@�&a�Q�7��f��V��?亹aK��'<�k�&:'�q��Kn_Wtn��?Ԭ�Q|�Q��3��C�K89�D��v�ݣD��V,�`��w�z���Z�=��"+x�.����G���P8	 ��s�(dwvq�fߢ?��A�#y���a�Q�*��&��3,�Sڸ($�M�*��E'�O�_Èx C�:T��3`��k�Y�ߩ��ꍉ.g/�'x�/�:�@���2L#�G*vj�{�?>��7��ـL�3���@~��w���i��g�E��廒��4��	��U{Ix�<��%�[���"E,o�PW3�� �a�ӈ\�Ш�ǻp�&B�r%��w�Ra>�.e���N"�I�O�I^h�s����^*.ݑm"��%���� ���s$�IMC�z�H���L�
�Q9�^��]��?���a���jE��|~���,=��[/����`�����ν.�5��cו�����Y�.����B{���X:T�c��-�v�0����o�j*S��@����'B�������w,nW�G�}@��Z�X�P9l���2^9vD�m��L&�(�)ټ�%H+C����U�	)�G����%�A�,�O蜽���;Y�Gg�+pjy�`0�Pz����Q�q�I�k����l�0�!E�����H�K��������Lc��Z�$��5l2����ڙ����:F��ޥ\��^帠	Ct�J�X������[��g��:��M��BL#$�\rՒ~��Y���?�WAފ��� pra��b>��;hMk�g#�Z��	���+c�[ܱ<�&	�(�⁙j`�^8�����q���mz����,��
�B�J�^U�s�7#��d�A wa	�ouz���m(�P�"�u/ZԠ��4i*�Y�{��"	��m������n�z��$��v ܻ�/�㔡���|*��t#��.>1*�zL�ЈR�ư�ĸ�T����>>W��j£�
��j���6�H���q��l�Z�t���Ḿ90_
��}�]���Ks?{|i#)��EW�W�����EѲ�@b�Y�I#�	H�����|F]���0�2��^��� ��x��bX�a�.��
c^$.�v����Jghc>�8TF�OV �4M��{�{��b0|��%���$?�U%ݮ-p`V�x;#�,�G�&64��'?~/Y�m�B�	䧪v���Kg��Q�HؘOУ:.Y��j�(��w����N�Z�R<\%pQ{���%��\�O5���@�1J���pU�2����5J�[ �mc�f`��*SS{�� �aj[�۷�	�M�,Ӝ���ʤp5�*.<)�hAZ�3�Xm�<__�C���S|����'���9Q(���
c�g1��3v��!b�-%�R��~<����k��	)�'��cOu 2��RU&�鄁��WA�մ`;թ8Qt_��ZpZh�������n�.Z{C�L~0�GHᅇýE�C�3��K^��`�J�9�u�(?�j	�m\Ws1s]���&�CD�0��ձL1����K*�䊉�yّ<�;�k$c�4��'�*�:�y}e�oKiWU�`^�%����>˚�}�p��,����ьM�UH��V�;x�r��%��&�lZ��1P��g�PV�э�E�o������f��g��L�HW�eE�W�h��@��������S��`%Z����a�b<�k���WG��kϛ=����|��#M��P��\�N�q3���d��Q�&��7h��6�mgx������z�牆���R	�<���sl��]i0C����j�nz"���Q�/	j�HU��a<sb��>��w���9;Y,z
�T�\�9����jT,b&=��R��l�9;@�r�<��i#�y�Rb[���"Vj���R�!w��o(0�A�-�'o�sO��:k*Ŋ>�hz��-�y��X������9u3#u��X^	yv����
�2���w����t4ܞҩ��$+	���z$S�n�1�`����&���qM�.���@H��S~�k��uF����ڱ��y�(�t�ZySO�J��O�"��ڼ_�m;�@@��z��*�/YIR칵>ȶzMuH��sC�Z���O��9Ǣ��Vomp�&%�̱��n!Q?�K�U�%��*���2�K����c���Kt�Q�i�`�&�h�5V`l@���N ���+�fʄ�Bp֧W����
Uښ�Mq�4c��95���t�^�ÿ�qf���(s�3�hd�m�r��Quܨ	� a��>���]�78I�?�z�9�_y"h��>�;�%p��T������(�D
l�UY��e.�v����u��V#�3����+��=��M[����u!���eR�|�Sl���G/77�[�i�`r��:щO��B�M\��l �Q�v�+T��M��-�QG�q*��3�]̍����#0�݀Նv��綛]��՗ob�_�k�*�i����g����l�q�=)�ڟ��`2��,�H_߹'th�ѯB��b
�)@�x.:+no�(@G�x�N:�Q%����u�뾉�*JSTGx🐇k�id�k�;��W���g����iY(���Emk������O[/���}�A!'�� �'��ף����Ȥ?Rw���{�˙ֺ�{�%�j'�cs �С����NC�t����O�G$:��[\7��O��� �mM%�����I,���Γ1۲�l@�&���YW�+���.�2K��� ��.Ƙ:G3#ѹ�����o����pi6�L͕�$�Z�	VSЉ��w��G�9�X�ay��M鿀!�Oё�>�H8'�Q�S(d�쬼�a�Qm��(}0�2ym%f�J Ҁp�����;���~VX�R�������\X��L���3����U�6d+H"�D�sy��N�,����\�М(��#Õ�5v�2�Jo�	+�D0�2@쿘}��cH:�y��,F���x�8�fQ2���q�����L�&�Kg薩��\@+Cx��f�o��ن��o����%����鬻���b��R��;%Ѷ/����-��qeD��p�~G�q'��#��19;"�px�4���afw�,d��r�+�,ei>�k|����H�����I�[�-��^ʰ8R���yH�$F=��[�@;%Qǲ6�Zs@�'� uB�As���ǱƓU���C�n���hYt2��R�.�>���K��4<*p��B}ʏ�@�D��4Þ���A�+��+�>�J�}f��d_(ք:�:���	Gy1���v����� ��_�ϖP�����ь/�H?�{L]x�ky����z�� ��"��h�`	kVs��?\B�A��������X�@�4-U'�<��ҧ����H�&���k�@"���J�T� �;�z/6���}�Z��$�v��F�uU��Iz��J�ߤ<�$:���SmBI�ix^��U�#� �=]Ϣ��]cQl�����>d�	�㘷���d�
��g�����-�������*m^�z�]!Em��q���aӌڳ���,Hb�$��#�xPǇ�&e�+p(;}lꐥ�u`J�g�/O��9Ǳ�X���g���^���w{����g6�Ө	��U�Gw�Z=�b��z������b�En��]��Hown��p��K39��k������3
��-���Z|W.�0��R"�[P����󌡄���7d���@��~�&�G:���R7�tdP�%�� v�7��O�Z�Oo��?G�=b�����?��`ͫ�(z�n6��F�Hf��������%�����'��U���=7�ǥ��`3.�A(<�`�$���$���1R:[���o��Z/_F��f:�4���w��'�7I��MɊ�Ee|I�]77)�}�MI;�������/��7���3�z�] ��C���'hV��Sy���S@ـC6�8@.,�Vs9,���94q�B}�ۯ7�㗥	�0���
��QP+�Օ��r̬��4ȝ�G��GA�kU��+x� ��ԧ=x��dDk� ���,���JFA�1�9����3�Ch��=W�N�����9�B/l�$��6$+�M���a��Z�s�2�dͺ)�}?M)6S4\�P=&ї��[�1���P!����z��Yd�s��{�J��ftrv���Q�<�B;$(;��by~~Z�i`����!(��������'�"�,'�׏�`1��g�q�B\����U!!��(��[yui��}V���@�ҹ�ј��n�Ц��o8ۻF�{0�����E���:��2�v]s2��9p3���&r]�:٣���&}i�*��ځ��4�ϭF]a�`��v��	/�M�f�g�9s���"!�WN%����Ӵ�hu�\�W&�BF���Wh�u��4�a}��;'+L�ͧ�6�a��yӬ��UY�r�t*����ȥV@�}*�{�:_�>�2Q
��>����|`�y�����Bh"�g���h�� s�1T-����<�q���B4)@͜(.���|n���(!ԟK��z&E9��5��E	/��F��	%c�N�t�u<=�D�󒿌~�b����7�[u���k�7�B?��<�~}�C�e�|4�z��z��C邑���'"
���&���V+�<�%�J��y.�7N�w��u"X����f�$���0Q��ס�6
2���-��� '@�����%M�����Q����h�?#X�ZɃ�v����$R�:��a�#g�b��~E�����wW�ԆHG/�S�|
g7 � ��1Ofđ0�FÒ�I�,ɚ�y;���;�`lzOY�U�G��W(5���׌�]�u�A������]ƛ��"�����OiYj��K$��<���Y�-=�8��럌Dƻ=�Wwmi�)$ na��B�{�9�C(ۿ���Lz������b�1��I�e*��E�}� �G�fů���AU�g7�~ٞT�ϓ_���҄F3��窙!M쪮2dſX��n�2��4D�楣l��m��]��]FlU��V�ś�1��ȝ�RK��1Wqt�r!w�˝Ϥ��\]Ht��˵������;9d�Y�ej���*>�,�E4�הp�i#�t��D�m�%���Vp8S�(�9�%��|Es O�؊{tW=��]Rg]�U���=�7������0AMrl�a���S����X�^���-���as������p%�{AXG�� ����ҒN0��0oX��x�㋖�/����~��H5NH�xD���o� '0�a)
O6�ð�@n��}tu��I˅/$	��~��{�e:o�������:'R�vScX]���Ä윪�o�N�GΔYW�I�s�;;s���Ö�<���pcv�ť�	_� qÍw�c�*q9<�b�AC�!����M��d��0a��E�pt�Z�p�kBBW��'ʚ�+���u�Qb��ܡ�@=��}痙V���%��l�b.��o���7�-�z6���g|�&1�g����\�Y��ߞh"쩍��m6�֏��m�4��m�)��P�s>RUR��q*�x���$qj��!�E��ü����~t�ߧoZkC���`L�g��v{J���|o���:��[�r��m�j~rTA�f�7Ƒ*��|޸2~b����2�)�T�S�y�ew4� ��q�s8���b�}<\�"}g���.cދ�dZ�ك_�:�_���/7�
=m�	�ך�/Le�`����l�٩�1�%���d#�X�H^�J2.tO�~(��i��:�&-�`	<��3ȃ��0�k/��S��"�&��B9�(��4!�DF,I5�e��Z
>_Ҟ=茕�x�s	x��QACʕ�� ���K]w&:%���7.p0�K��@ÆR��ⷉe�v���c"b_�iQ�a��D�̓G/A
��Ut�|���,�?�ښ����5.Yݟ���VC�SP�3��V�\O��-�Ax�-��ˤ	���X�u�P�r �<��$ȋ��z�����=8��پ?J��ld��C�?V�84;N!�fޞ� ���mR�YŒq�A�Ý�2�1�KO��e����S��#ќ�w����~����%�Ȁi�n⧺�������|6����Ѭ��X �f�龱wX�ց���/or�ƃ~�{����8u�L��� ~>9B$������ޕ�'N��	N�b��"0Ӓ�}�QG�[�#��B��RλH��>ch��K�Wgº�>�f?�M<��f5;?x�NP�ޖCU���:���(�A� T6k�(th�V7��v���~�`����K��h3:Ǻ�>�LPDAS���1��k�Z�,�
pW;ۥg��n�'���d���q��;�w<2c(m�%Do��X��$��^�˧
�և��M~1+�$�5�L�Λ��(o�h����C����|5`�&�fB����'�Q�1b�c��k�݂���;W�%$�_2ك�5r����f\�A.�{��� �_�O�c��c`T�rLP�5��G��Ti�A�Qr��Jo��p�V�k��w_�"�"g�r�oҷ��L�v�ZE!����w;8�Ӷ��8��0H}|'���s�pӷ��0Z�yt�g�`.u�t�f��!i�vO;��9��K1���k �p���DUÑo�l������F�!��|���A����;�&�q�Z�7u����N2��O�)�~ב��2؆ޥ2�����`*S����T���f�I`��V�u�1d����6��J��s�%��,_���s�I��"m�g��f���!#�&�`����4�LGg|il8Y	(�a���1,j�@��7�c)�A�P�5~cP�n,ӛ�+���u<��w:J��.\�#o��V��">��� c�)�}anY�u[�����tBTo}��wQ&�<n��{� �ѲO9�<Bܒ{\􂉦W,H���X����x��S�V21u'���F�m8t����������	7-P�c�s�"�Gk�ܹ���ݚZg�5Y1&�b���.��7���'���nT2�8c�y������'��p�%���V9W4��?U��5����'��������HW=�/�]�d����}���6���8�}�V�T����݆C��!>����#C��$�xֹ��C����Q�%��?R	د�0>άF�)4��r��k&�f�?|6?� 
������&n����0!�.�{�r*�_�Q:g�����d�F8�����C�ǣ��*�9N���N�a(��з��q�Z�3G�o�mX������<�%?[XV#��q˟2"�0
R��r���ܟc�6��<�&�	E�e�}ͫ�R�D��&���s��imP��y����f��g�Ox���>*{7vx0SN�(��~rbp�%��jV��O2���������nR�Ŵu#�$@�d�-{�7�<\U!�e�UOM۴KL�N�}B1��*�0��K���.�̌����2����)�G-V��5��G�ۄQ19�I�_[vFv���Cφ���'�Qs��~%̮&*�f�	���f]S�y��D���⛀δi2h�g��s�x.8�urF�,c���Y@>M56���r�V�����e�S�<���`h5���3�]��Ч"z���
�
�?M�� ��*֡��r*��$�/�d�r�1�Bn�,j�T��NM�DJz)��̫�8��w7���ȳ�'"V=j5B�z#�C��r��T�l�e��&	<�:���n<A�����6b�
�TX&�S�M�ktd��s�qۺJ��NB��Sc�U�;b\�)#��dîYʰ��0:y�A���(�}�Ҟ⡪��N��2T;��ȃ$�����������qu�,\b���Җ\m�h/27Q���R��8�mPO��; ;�"�b�Z̺ź�Vq�Y i��S}Y4m��4��&�<CVo�k{7_�د��༢���V�vǳ��>��x�����U-p"a)[_�MhEdx/ʟ:y<�7��Z�>��e�,�糹���#aN�O���D�鷍F�8�$��^�8���9�P�]����ISb�ȱj�|bNo�~{�(+���޿���K��P#�,�g�����3���/�%���ζ�
���N�$�1sb����Z��㕅��pW��?S(�3���q�� ��I(������s=7�L�cZ�Pݾ_Ua[��*;��:���5�(CD��"��ӊ"+,���ͳ�@o���~d�)���Ǵ���[�q�j���j$������|�k�	Wh$c�����25:kVY�I�HY��ę"C4�G@Q�� $0����jAA!�zYz7rSR]+οv��J��l���#�Aa��:��{�bZ��duU�`F�eF��Sq���H��v��p���w�Ņ*�Ok�(J�#r�nN�0N�8���.���Rp{��&��%�3�;��Y���� k-'��u�^^Z�|yS	=�P�#B��l*f yd> ���	��ԉ����|�L�y=&R��I!���6J�.p�Y��r��etH�G%�c3���}���֨w@�$k�4{�4a�eby�?���nq��X���𵿼<���%�ڪ����IХX�r�]?r�Θw�o���w�(��zF�3���}^;Ê�/2��gh��@=x��A�/���i~�)s��eW�c$n~�6��h�L��tKq�#����τ1V��1��\(���k�s��-#a�Ol6ە�Ş�G�*t2���9C���n���_�"��T/��a��U�v��^�N�Xw�զ*QZ,���bi���krd!�z��;��%��m(�3�N�ak��$-��V��f5���v����!�
�X�Y��fKZ�37H��Fo�+P�#��U�+}��􃚺�G���754��@��j���p�|]�w�I�Ј[�`EA� `��Aj�?�pCMG
v�����au@�[��))������=�9�g��&֝��?-r]%:�����Ƞ���`���١�3Ex���>���
#�����NWQl�w�Fj�hto��NՈ$b��\	�](���a����H��S0Գ��ύ�~J����;u����̔R�9I�wCw\1�d��%-�6��+Le��YkL���I�F�0	�գ�]���Yr5(v�ك�%����D5f�҄Z�����B ��6�a�!��'ȱe՗H��n72	��.B�LF���r����9�&'`�%�]ٕ�j�J6b�˖�_a���aS�`{<���sc�2s��I�`�{�H��)�A�^�4�P�#O-��aޑ|�:�~J}�!�*H}/���N�\4��ֻ�������mFT� ��'��h�D������� P��#EܲS(E�a�`�UW^[����#][��m�i�V�P9����ق����]�%[r'Q�A����x뭿��^-
�g�M�����4���̼�`�/:
8I�%��'GqC\3���	�G-���L&�(��9R���g�w�c�ޱ{�V3��T<���Aڶ�����|�gu����(��
�xq��_�|b���w1L2[` ��60���k����JxR��Tz����=αk�?d�m�5vۭ����v���n��B���)[�i����Z��<4�@��6��~t��o��WVՖv$�?KJ}��#�RO{���.J�n�]Kf�G�OW��ld7w�j"x�F`(�	���PX	������aI��� �{Ѕ����,�S���f�
���}'����N$���ECܭ�)��8��JNVQ6P��!�R���_�u)��Ap�?�%�.�.�"��>'�+�P0�F"�{�,K�v�y`ւȃ�h�&�܅���ú�twӤ~�w�T��z&�hA���u�i3#
W��6F����͊ţqfr����ܚ�:	�͗,�P��\�E~Ay+~�����[a�����~��H��f�{����g�/3+ج\���k���F�`Z8X�����<���ָU��y$B@es}ق%m5��p�{��ǔj������8§��%�,����n>OU�_�%:��
S
H��fW�bA�vT��YQV5��Q�j��K�9)St�H���q���ef��A�����/l��Ba�k����{�7���7#�zN5��x���]�ue�9τ�����Ä7���hakx�k��QY�GI��5��VJ%�~��%Gf�Y� ��9��g1��)S��bA�B�6=@|I��%�c�|'D�Xg�Lf���Ħ��%�3t��������M�p7FCbe�4�*lK��G���Tb,[�) zuuFD?��\ͤ�)�}�δ�z1UF��g�]Lm����d���}ʘ��+�Oހc<����M����pĒ�.�&���	-q�B����CEu[J��65�R���{?q�$K�l��A�}�O"�V�PUԪͯ&9K(}��� !_�N�$���s%9��d���.&��K�D^��i
jkGe�T�	d�.�Aѣ�>a�1����h6\��`�6���_l�'&l�b��c�B��þѸ=D68c ߟJj+��2&e0�� �a��+
p;��`t`���8�r�����x@*�ǂ��3�̮�oU4�̗Ϫpj�R�����[TI\
d�����I4'2�P��hJ� �w�Cb�\����)RR�u��X�x� ^O"�h^E^�|Z�*!��^ͤ2�����lֽ����.���6�0辤rVһ���=�P�ȣ�%��9�
"?��ug� �� �R�I�T�n�D{���G�2_FϠ�$1 %�=V�Z H����k����]|�H��Z���iT�ٍ�B(ʠ�����sJI]��8N��'�`����,< :,�����'a�o<�n!������2���3@�`j! )y]L	 �!it���!0:�C�b��XHoKZ���ܘF�}�QG\G���ΤR�����#�PDg�������E�ꡜ�����>��Ŵ��u�����,������>9Y�@���WW����-���(�|��b�$~�D����z8X3E��L��gEBv�1�0YT��"�,����ȿ��~a� O|~gg���&��,�eCs��/���z���DL��|s#[sM��,�nL�s��&�;EY�[MX��Qn�׮E)K<�wg_�[s�اT�D��V(z�]?�:�K����R*�m���v���q|oQ�����0cK|���]#���d�]��z���Z«�r�9�>fg���CuOܷ�I]��ߋ��i�{W�{9l3�f����uH��6�ř���q�r�1�bA7#���r�!�z�EB�Aj���I"I��������ҕm�8�=]Y#�K'-����	�!~KC��kQ��S8�,2C�1a�� �[Z��X�����p���U�=�xC�ՅsͬSI�|���8� ]�
�#�e,19�V;�T)ɞU�Z��8����6z�OK�R�
��=��k�g���$�N�'���K��$<����5r�y���LyK�C��>Y��ԟ���O/�2oq%7��1���Qt �u[��p�D1���͏�?�H��T_�k�wx��c�� ��d�U���:ݸ�P�A��a��:L�E�?���c�|����I!N�����wڳ��E9��E�
[��l�0�[�j���^H�λ,��\Ic�CC������|K�f/ʙe�O�`~ќ���E�X����nmyQ����Cv���o����0���H(X;�����JB?jDe�1�`�M1f����xH��g���G8}��ZAYJPo"In��Ū1�պ�,�!]n��oxe���߶��QP��m�%��x��P����#��Uz�2�'N-I�������*^!P��K��%�0�RX�M�)gf��0��Dr7/5U6D3�̈́4gM�:vCr^��{�nlC�U��w�a�63̞��Cu�e���>~n����P����&�lŋ���Q�W�i[+h�;*I���-��mWU*|���4�<�ŏ�0�~i�`_���9<�J�˪��R�A�-q�|n����F�u��q�	���W�� ��*y�;�������G�X�VdB�DVh�r(؛Q̖j��K�� 
ٱ�W8te8+�|P�be"��;��42��w>���<ZAwv��:q�f��������yx��\w�D�i������yH�g|;p�`K�sP3Ct�ۃ������u�K��l
g� \C��vTnt:X�:�I��q�OkF�������>\|Kz���D�e�!$H^�s�����>�V�_�$O��&�;�ij\]���0!^X�]{�� 5��m�>�i4���{�̣�ī2����
���<C�P[�`��j=B�(��a�A<�x{ur����bMW͋�Xۙγ��Y�:�M�TĹ�<���C	5��HOM�i[G�T���I��y4�!kX~����BqT_��p.���c���g��NlXozIx������
�
�iY#�
M;�|b�ű���e0H��0髦;��q1�|�w������NHCeN��g������`q.�7�3*J���8-�aos�w���^ )%������.m6�E� x�ZnU��i��×�F�;ĉK��f�8"��vX������2 i2��)^�`��d���I�
m�|��hG�f{�_�=��Hy!0�E������}	�ʍ��`
�>d�G��4>wM2�ž�>�UW�Q,K�.�l}�h�rӄ��e����=P���Z!����0ފK-��o���~�f��2:����-�I1/6�0*����,V��Hf�]�;9[�C���~{�*����Q�bk��B�:~e`�P9�s>���'�X�l���-��1C+���K�U�~8'g^hⰺ{�L�Q�������SEشe=z�D^;N�B�Z̀�S�"H�j�<���eJ䏢EOE��A���XVr����n��(Y0��%�j&`n0�����6q� �zġ{��;M�S���a��d"
�e�����$�F��I1�P�\ ���[-�m��H��m�R�����ſ�5M�N-B����?�k��>ث���<�Q~��mS�Bf�;s�`�Kx(�KN�Fߘk�N���S�L�B2�������N�-ݎk����*�m�BB@� �9�4�1���P$\X�npi�Jn�.(�+ @VZ���:���#�����Ŋ�qQ
O��@R%x�:c���fÙ(�]��r���PF������C��b��R�U�������Ԫ~���D�{5_�i��g�����>u�K��������G�
�y/�35��_�"B�B@}sۂ�W����6��"6#� ����Kl���!D����f���"y]�X����0�t�<3�������ٷ��Y	&��]����� p�,��8�%���8�e��7��NM�� \9�EK���j�:]jZ!�EK���_R ;��C�tu�I	,��0F���s�oH��ɮ�I�#Y����f��g�phΊ��ysa�B����g
M_0՘�ʵYn�:�<(����P��"k���Zjk�6�-嚻 �;ܴ��QODmm�BUс�Te51zq��'�DSИ�h���_&i�W��������T�q�D�M��b%x�Qb�zˇ�&&��Yp�T���30g������?�xZˈ���)r�a��h{L��mim�DU'�;��`f���^x%��u6pv�� �
C�����C<�Jg����P�E�ă>��Jɺ�n��o>"�|s!TI���㸣���{�b佦����uݏ@�A@���z�"�6ڬ�#M�
��Z��p��a�'���z�4������e�����䘸��-�L�0�K��jmN%9�.��H��P�ؠ�N�ka�RP�:I.��a���.�Jb�����>=t�%_B
suNo'�sy5|(���\y��f��{�]y,&�ƹ��>	˖O"9��#�����-�V���rH���۲')���Y����vv�A����G�>��q/��o:�ڇKJx�u�}����眑&�0-� ��J�&����� C`��ʂ:���l;^1�^:�_�*ϢRq!5:B��ZZn|u����\��a��D�(�?�x���~1D���BᏮ�ڔc5h0�?u�N����p��8ܼ���2F@-Gl2��)�5A������v�q����51��sjQ��ضHAH�8K�l	����Q��D��d���,��TV_�q��%8=U��\s����
Qc�<Ǆ�)4�cղVl2$z��Q�06����l�A�ݦ�&[b�%��>2?8ΆNb���{�B�#���ݾ���!$����T�%��B��3��]��ҟ5p�4x"q�o�V~`#�vb�x1�;%��l-�[l���&b]�>�%+���g
��8�7�ſ��8�Ȯ���v�L��=?��G2���DH�����i�v�	�n�q�ަN.:�hS7�F'@▱0i�:��aW��X��\OS3w�O�(`ҜU �g�-9�!���3F*��n�sqe��f!�S����b�����̲�G��v���Z���u��� "��Y��U��g��EC6[�@��.yr��R�.?����n��A!Z���Z���,��!�R�K*i*C�hލ ��_$�6K`$���}Kv�"�K���� >o�/ ac����&���;��y���8��T5,��)���Q�k6{�#髗㎘J��OaeW�h�!ɤ��}c�ƞ���{ �D�9��]�/C(�%Hj��u���&��NYL�2�+��A��/���e�9���z�z3OZ	�Y��� w�eQ�
�1��r�"��R�z)d�
y�~6F���$�����)���~���T��bL J))d�_(:Z~�^s?R���E]�P�| ��y�����/�*]ľ��1}ϥ�¹�e��~����"�-@M[\��.���u�Re�?�>�$u2ⴳ��Ә%j�nfg�p�(���@��;.j���.f1(��q�;aPQ��ر?A�ߧ��4�^q�� Gd�iݿ��w{�&�]��5�m�S~���Bj��bH�p>ͨf�Mכ2[N��,�9�O��p���ͅ	��ɨ�9i�q\��~]�~ġ��c�~�y��[�A#�"���U�o�9����9�F ���yq�e�*Y)m��_)�׿�.�0cx��l�9��بaM��U��a�C��Cє�c@��1�feTN(�Yͱ�#g֭�7o��1;U�#�a��)�� �0��g�])%"U\9��j��QƵzF��/2vy�<�Y뢫R�{Sڶx�_��H���_�p�_󣒅zi<��j\w^z�$���R��f~e�r i}Y~����	�mt���J������z2"��NM(��[�3^�iI�V�j��������v��`��EJ�R����*߃��$[ľ��Gv�GS#
R��9V$e�8u4Ǚo�$�K��B�{��hmJ� �ڄ�Ρ�	tH�a='���:��ڬ~���z�mI�p�a��[�H#O�K�C9���<q� /���/^G�aPU��om�J��(��"������ �k>����@�Ӳ��f�̙v�U�������8	Ǜ�,6���#����������LӺ������˪�����>I_x�ZWV�`�ysw�V�
f/|�m84��v�M�#K�*��O�}�sI�8��`�@䵧{�O��X�-t�A�u�u!�{����'e�H�]��ģ� ��Rm�b.^	�^ݮ	+~,��^�`M���V��5�h�n\@����<�ڞ��0���(�<t��J��Po���?R��N�&�&�\�7�\�w7���l���������4f�V�Q:(Lj��}'��'�+
6�|Wv:h۠��Z{�Fd-��Zm��ům�_�h�.q)e������+?��=�a�jl�O�(@�Rol�oTk,3%�v��� ������1 W�nHWEf�A�V!W�^ P�|Uz�0��|�I���8��m�F��.���6,���28���&m�E@X gci��8�L����E�B�2H�l#��SK���_�G����r�a=H����ݞ� �5F/91X��04tXL2���ca� �]a� ��ݸ#1w� ���Za�w�a�r�zC�8��H7���0���oo�L�୦�S��/�MV�oZ�K��uJqv�O1�f7E}�r_
�(}�;Ϟ	� ���ɷ�^u{��÷�����\�F���Y.�l"$ΰT'X�Ґ�z�#B8�F���)J�z�χ���8�D[9\��b^o�^RtF���!ⴞ�Q���E[�31�W-C��_Ռ�39)-+��u��--��u�x~X�xyȖ���b��	�Ȟ���s@�H��1�<�Y'
�7�x,��.ɧ!�F�d�h��:��5�F������![�BPʝje��E����㱰�A��d;r�*6L��oh��~�h��&0PG���%h5����)q�ءl"A4�"�<��3�>�.�# X�Lr�4�r=ET� �>��.>���vf9��UW; �0��.]�'�.�l5J4mE�Pt���04,.��z��_�#��9S<~5$�QT��<�a+�4�X�XM�Y3�[�aZw�܎Q�Ҩ,���6�S.�rf�°դ1WL9ʑ���a��J��	C�M8X���{��=�����ɲ �N���V�E9)V�bv�c\�䧐}�	U��x��ێ�$���-������` A�6G*Pxw7��f�CdXa~�e��C�x�c�
�Y�md�/���b�,��U0Y.�j�1j���=|�S@�pn��g��s���C��-Y�<0b�@lc��<�6�CX�P���8�b�t���_cֺ�F��٤�Y�b�U����,�k��GM�;��{�����3���|R�t��������-1��S�W#�os�8
��3��O��K�ZK~��m3�j�.���ތ3����Dcln��iy�QC�߻����h���κ�6��9ϗ�}Lԋ3�Z���Γ&�屨������}��ﱭ�v��M�h��E�޹Wk�����c�GzF���.G'�ҾB�����a�=�Ts�W�28Kl����� w��=�<0뺕4�ш��߸Sơ'@��7]Y���U�ڀ\5uu�󘵲'��+��4bn�}�.�E�4>�4�2mC���,M��N�f� l�VDj#5�� ��e�<n&|�������d��"V��|%���;���ׁ�j�ќ��[�Ӊ�1��1�,Օt"�����x8�}���ˮm+J�Bt��H��奷���/��T����Dw���_��0
\M3�#&���}�g������K(Y.xȟ�%:������Q�w^�Q�5P `�u$ٿ�����yu��N4�}�=W���:�J#����d�ٴَ�sZ.[�a�,�q�PmX��g|)e�ܢ��t^D�E��-8ۀD�>h��k H�CT�Nr�C�nӲ�sc����`E��@���8|jwV��JU�Q�6��C=�L��@KU�����B#3�jD1�O��"`C�qn"�
Mc�Ee��H. �:0����^�rA��|W��S�:g�����b���e��^τ��Q�ҿ|�C��JU��� �IiB��Uͮ�ޢ�gѷ�؏J�B��V�H��{4W�#���t��}����J�e�0>H	-����UB`�=��V��ȇ7�<� w"9C�!�����փl]�@�]c��V,������٘�	��-��=�P0����i1���Ptd>����0p�B���˝"^e�~;�3�e���H�(�$���9����)�11����NW�A�D#�i�q�,�K��s�`B�/Y�|r��@CbHS̙�/̤�(�  �7��u{>������~ח[U��B��%�e]qz��8(���-�Z%+j�8�k��DQ� � ~�c��������i.D��*U�G�[��퇶��u�>�Mt�H{��h5��@�iS�?��&�������$�q㗽@�LP�t�ĥ^+��1��c�&1��yВҪ�Y`ѭ�	�3@-����
5^r�o��Ai�Ah5�6A�	�P�b���O��H��j�yܢ|Fޟ	�-o�_��+���e�Q��)�S
��)����3C;a���z�U}�p8�%�[��NfF#S�p���]s	�=���>�Y:���P�-~P����v�l).A�A�9����U&��R�
+Y�H���m���@��kd<V���[�-�[�����K���zS]�������u�?����������%o]�]����/\��j(��?M:�P�i#I�s�m��*+4S��{���B66NˋN���GL�t�>�����ݐ@~�T�`e'uw_��,0�.L��TW�������� �$܁��?�<P��m���]�i�^��/!|vb^O������B�X�T�~茊[�s��AH&�Za�!`����h��Ã��ڰ:�7���k�hP��]F�4k���j��e�Y�庺�d4��A#��x��W-G�O����B2�z�W\�f��b�C�%��}�1�6l㈉���Ǳ��KHsa���� �Q4VhH�c�J ���L�>�Z�hu���܏9"��M���.]��QMkr=a:S�=x�yN�h5Y��OJSu��7�������C��@���Z_����o�ѻ��j��Oҕ}���f)��7�I�ʶ8SO��!�]��?��HK��i��.�Ч�@/�j�	�<b,�͏�"%�y`���!���^H�ݿ�nHA��r[�[뇏�Y������{L�<�s+�~���me���_�G��m?��� ����H�l4��XR\�
j5�V}L�YuG2�����͑��׃�� %��/1��Xr`�xZ"e�b�{4��&���o�����-v���cG=�j�'��Do�/���e�S����<K�wP��s׆��Pz�o�%�iE��,�ϻ�WukKg�<8�&J�n|�I������pP��J������	�,�!W#��?_���Z�[���YO�[Sт��a��%}��)ؔ%��LzI�����7c�q��X�xl"g��]�R�xU���1�G�D�F�ߜ���I�3x�D�Ĝ�����F�+	ؽ�����JQ��G�	ڠ|�T|���u۳��m�Aͫ2�=����1-���U&��������[�3�t����|��¡5�M4(�U�%�Op���42y��'OvE��9;)�_�0A%���o�an����	�옼ְ-ZV���PmT8`��̸9�a̕9�me����]�RY�h"V$Ee^��.�`�/�/[	�2��L�w�&�͡�2�V��B4�΀{ l3��YL�*�!^��ۧ�Ł�C[ ��Oa֦B4�c��9�����6�|,�m�C���I����f;T�@��l�I�qr��	U�Ei.S�1�ti�}?����'>�>�+�	��0�	³I���뚯4�i�C�gC����h�BzYE����P��F�tw�3���_����͜v�:�Y��'�޳�M��g���z��˽X��̃ѥih(��i�<͏��Y/V��"!�k_�M���[MWX#��iK�_=��h���g���)��D�<�nx?|�����&-Ò:�"v�P_'
<�6�Z	�Z2 @�yp�>��Q��J�m$qD����{o���a8��� �#�N:��b����7 n<����BB�[N�3�uy��:��I����t �B[�)�x��D����Ue �x�0�h�0��qo&h� ��O�yt+�|�.�"�-HJ%�J���z=p�#���k�J�ШB�-p�=�J�e�`Oήʵ,eH�����Q(�Q�繱^〆ZA�;�����K����l.��EJ�`_��X���B�� =O':�_;���HaG+M��'��r= ��1�u�L!a�k3GЖ��2�q�ޭ4�X�)��C_�6p@\�>O"��	�0�Z�� ��urh;��ۆVeaȁg���O!����r���W{
f��>P�v���Qe]��'���^�=s��� qp*�k�����'+�FN�w�̀P�)5DԅU˝�H_�\>I27W�q�j_�RA?����6���u@���~��u��3Z{۞���_΢�����TG���04 6h�+e�e=.���}�U��2�$�K���#6�ŒCt��I��k��;���0s���v`-5�և�0���2,���������q[y��zQ�o�]�<�8k�R�+��O�Sv�BUM))������&F��(Y�O�~^ ����8g�P���������e�%~3������"
�q�0�����̽�͚��%ǿo>N�+ʔ�����
-���maZH�4��**�j��%.�[i��L�ltԿ��!8k�15���ejgM�lt~���`8h��m)C�f��o��WG ��]Q���)Dk����%���`:=I����^:rp��xP�ⳍ�9�>x_0@�ObyG����@:�5��'��sBi���a!���	��@���~�2v�J���9l/ �v?���
����:�%Q���lV9`����w�4�b�j� �2 �&in 8{2�v�:��靖����*
v_�NK����w�4a.hw�j���vJ{��qC!K��v��W���h>&�!Ҳ<I숇�jCA��]q*���mvwK������?G�>uuE��7d���r�'���/)�� ��_ۨҞ���1��.����{�iC�wi��	������
�	��_R��mS;�I�v�5�[Y\[pq_&�	no�[�����nt��S�j��1���]{zp�%Xiv�d�,A�Y���F/���]��TY6��6>jJ�U1��q���}�4���`gq����5?�@MF独��)��8C'"�C{�'�泏���\UD"b��.�M�Y�R-�A��7g��V����^��;]!cZ��0��V�t�u���/@�&����:f���J��@�'_1R=p�Q<p�������!����
J�s�2�gl"D]�6�S�s����\L�og�L�`�ɍ�u�?�+�����q]&�-W`J�."005�cLw�1��_�x@��}�l�8ђ|/�A��5�'��E�:�����p�@�i�������y�D �TN����$R���GҚM�B^� ##���P�ɬ_�����z'�z��I���D�|5��N�!�g�z��d�>R���c,�����Cl�
�S���Az�p���SrҘ��Pk�y��M�T��:N[#�\�3�i�g�t���S�?(�8o���`_ީQǢ��bH��¾��B�|;'�Y Z<�t#U��%�M[�нw\\�z>�ªm�e���ՒYA?d19� �����
Ƃ�J]	�b�:@ҋ�� �����E�i�kYΒ&�W@d���t����l��LnJB�Qi�~��S���_�m_ǂʬ�Tԡ�hW�Q�wC�9kZ�=P����2Z���ϻ�i7��igU�=p������q�+�r��P��>|؇I�4���������*���rIQS	X����6'��=Y��D�fÆl��9�Y��+҂�����E�1w"Ԁ��\ם��]��Cb5p�=�,_|[�rh>K���=�˝W�Ir�b���>�{h�x�Sl,!I�{Q�g��I��� �b�@���2�ٱT��x���|`^iie=Ё�	�a�r14��C��NlQ�\�g�~)�y�$�8�J>@��������Y3�9U�f��B���vV��`;/I2����SJ
�U�c�ͷ��@Ug��5�����gT�e,m�T��"��ɖ[W�����7E�s�":�׸��Ȱ �X��L�WK>�-|��Έe�dP���	68x�(�M˂|��ĀЧ��zy+�8t8��>06u�D�F )��S�%8��g	��i��q�n��c��(�@?)v؝�x1��;����xD_�?F4�S�G:f��ߘ�}i���ڎ6�L,c����\������6%�d��IFHy(��,��άdЯ=�{e�����T8���8@��+g�DO���&���d�h�/��P��m^Z��%f�J�Q��s(���yT�LEm�;fr/Qk1�#��,�����}��������KY�BO���X�)b�� ��tA�k65�˓����0�w�b� ��	��w�"��䖍Y
.����wE�'Θ�����>�0�WC���=�#��y1���Ca��ԛ���A�������H4j�_�C�7=^|���iG[��ι�o��
����C�e��Q����y��@�a�>��.�.��,�ږVꏲ������:�JO�[x�d�y�Y(=Ƀ���	MIv%S�sv���v����q-Kl�mC$�8����t�`sk�ZF��x�?���3?��{x���&�5�L�q��d�NA�~��
�{U�c�a��û��TT- �F�Ñ�|L�H@8�*7��^4pp�Κ��'U4��#k�P��ӱ6I��f�mY��e�o�6l��6 ׳ȼ�^S��E�7;��^b;���F�8{�Iv:��r��φХ������u�qm2s �d���3�vV٪�%���<�v��i��r�6a����4**�cxfJ;@\"v�+<�}�]Y���4�U�5+�ϫ���i�H�ׄ�]�P�!�#K�T�i�����-�nm�L��;�bp C1������e�q�Pa����(ޫul�,�����ճ��o�dک�-W@0n��Ql���_�� aAm��h�V�'��OS�6�����.	���(P��Xw{��C��0���=�N���!&*� .E��ae�@J�B@��9�wI�&�g�I�.iPF�g�ǌ�j�
���e��vK�b�ֈ�:��(�L�8�h_�Tk�`:�/�w!:F?��
�R�����0+��D\��3®m\�M�-�g��YMSa��*�T� [��DSH\p�8G�u�~���L�x�0LL�CV��)�j�5_���pim��i�Ϝ����+Ras^�"�[O��9�"3落!ܧ��X�I�-�e&{KS������qB��������x����8)��7EV����Q-���p�H�w sq�I^�xc\����C�	�����9͆��f��V��,y�:9]��F麝B�� ,m)��)m�E��K�58,��)����{�;	�c9e>�j"!�"�$4���@L������q>0j��m�`\ ��^�z��$Q:/0~4 X��x��FX6#��{=�3SI�2pD�*j���}<�➏��sRZ����>�^|&o5���!��{]�����{7�#NPK���j��������z{HL��HU�;?�̏^}՚�B��{ ��R[�mT���bM!�@>�`�>�R�<����+m#�w4󋠺�d�n�U��E?�UG�& u���ߟ(XM�x�Co�4e�>&�l��"�mn�n'�:9z5@��au�Ⱥ�P����\�$��#�=�N�;�}�־as6�PL[z�}Ԭ����H(�@��p	=���x�J
Xi���7%���eg��ߙ+9�p�j�<)�ŻF���'>����H�>���N�����D�G`9\%��H/���\Ѡ���Λ�R��Z5�@׋�\g�sȿ��9.��J7O T�͏�dlW�r��ɲiqcNR�i$y�~Vneԭ���4G��!��Y��کc/L&ӗ��(T��Y�WI%�����y�'����������!Ō&�j&W�6U����b5��8�<] ��Ӈau�z�Ua�t6��rt�� �yձV�)�#��F0�G.P`�_D���0soA2sd�UR���ַ$^vҭ(0IL�RA/x&.�>,�J�bA�l�՚�d%B��@���U�M~�u~Zl6(��EJ�%�'_�C�m��`������=���ԁ�κ2���ړ��z��C���j�Ğ�� nD=Q�8	;H����p!�(��*}��ߧ1�K�C��>�}��}^K��T�`�v;$�6<�KxRz9��:�c<��$8!��Lih����q������*n�l��G�`0�`ex˯^]�\�	d,�_������>>�1�y��H�cDJ�`���&���L�j��֋6M���L�e�X�)u!�'�v�3�R)^(n����4�1�۲�܇�l�ؼ0ey:-kaB�m�%�T�ĺ���h���1ڕjrGy�|}ջKaw�;Rr���9q�1����\:y����'���Ī�&�t�����R�06� �c1�Q�KO�)���?��rv���f��-�U���*�kOx)�ʄ����W$F��j�1�>�|��`��ͷ@�eӊ��2v�	��y3�]I�PJ���2���Z�9(��=����n>�EX*���� <��q��Q>4�1��A�������*țC���hۢC_�*�L�`ik������P����ǉN&��b��E�\����!0i��%�S�����`�T���ԓ�6�(|5Z��p��	���Ԧ7KPh9���V�:�l�2e:]0��U᫡w�Rb�)���f|�S�:9^ZF���;�ˍ%�g�23���[�7���.���mz���!ܲ�l�ޘ��]���v���L a���D��W���H'a9P"�����H�W4f9�"�y�HU6+iȧcY�>�Z��*��Ƒ;\���ǚ����B�<���s%kK�����@���~��\ek�veU�k��ln*��U\�u�`D�>F�X�s�JJ���c�����YC�џM@�������>;4��y�*|I�7L��q6�i��e���#ܓ`�����m�C�ծ/f�ޙvE�� ��#���	����j�bt-uO45CO��\l���5&`�G|z�lD^������Fk;5h�`g:��$�>�o�Zx4�Te�جe.�j8Q�g����'��{ϴ��G a�="ۼ*�b`�"}��ڊB*=�7��6Q�/�3�{��5/��C�5	�e�y-�ܞ~�� n�pL���D���Q�T%Y���tz�M�!�i�6�9_���M��� �#<ė�m���{@����s�S�Z���,͹�ƴE�gj��e�sg�hD��E��s����z>P�4 y��-+i`��y�p�>֎��C�(.%�jǏ��Ϧ��I>Ym�G9�	�M�0�<�4��3�YT��h�Z2p�QgW�LqF�ϾE�)((��a�f����l�b9��}�~��X�Q��{�-����6����p+�����8�Aa�/�;�,��t��V:L��=_-�"�ݞ��sDC��!�!9�EkP��� ��<l��/d��.I�L��=ˏ�����rBK�ޓf���5�'��s�C��v�>g�.�$"��o�u?�Di�c-fL����5���ɹ���LQ��W���1?�l���o0�YY��gן�����u��n�3s�T���A]�TpEq��5E]��(H#�u��!��I:?
Z�i��Ny���Q�����'}���@����:*t�:Mq�wE��t�3�z�\Q?���`���Tz@�ͮ+�Y��d�J9��VF軰G�IM伳�F?
מ�рԽ��ˤ�޹�)��6~�r�j�ԃY�[�
Fճ�Ĉ�a�1i7֬���b+=��[�u��D� ���{�dj�j()���ha���G�$�.ZX;��]��p��5M����-�4b؋CzN-��~��RgO�;죮�h<��@�HOZ�����WSp#LV�K��F�6�Do�0}�VF������1�?�ޔۨ%����=G� ��
�K�q� I�|qC�;�w��Q@�=CԾ�&y������u�$^�3�ݺ��z�d�k��:�Mc֭}��]t�F3�q��׌3��>0f$�@��P�o-�k@�V4S�-j�߃��2d��M�;�z��̔�����x*�L�d��/�&�JQi+��b$���`�.�qW3	��9��0�&/���ŚL)vj"��A�sF��M���cU,ꩧR����C�0�u!x�^���ExB����(��i�q�2J��B��r�܊q,˺��[��%����II�N|t�!|*���8��}E��c�j�C�����Z'�Y]Z,.����G��4�C[i�=Egȡ��;*fbp-�o�I�M�*�M&�m%��h�F�u�{�l�jf�^@������l�G�����Ei��eH��rͯ@��c�f�&&���H��A��Grc�*�'@�o��HG������=�-� =������S�#KK.�QG��(]�o��Y匡�eb�J�Ÿ�h�27��M����K\�ן�Gg��7�*g~>����m�PS��
�2��wr��'�q��h�\������?�`���(��q���WL8AimF�����g+>v�*(�[d�����ėwɷ÷*��in
3W����s�uѓH�㜘Jg��*VX�H�X�� ����e�j�Y��Ϝ��>P!"LB�)����/A^K?g�?F�*�9F�Z���	z|�<��}vA�N],Ϫ�O^�b�&�K4��p�qT���w�H��D�y��ww���	ţ���$�U����}��!�K���m�|첮|��U���j���9j����ɐ)h4 �vG��J�Ɖ��z>�SS������Hn~��o��A<�����e0���d��1�c�x=�E)#,E-u�׀�! �	?- I���jΓ dԩ?M%F��R+=�+C/S���S�UO�>kY��y�j����@1,p=�L����t�_��F�����gzp��Նc��-�=�C>�F�Mt�U����z�M�iJ�(�J���TdV�p��r �O�+�'�"^md�ا8@��c�u������-�ed��?0 ����q���[34�s-�N �ᄤ
�!->�Zv'l�՗+��\tAJՙeK5�����8#gB|���LB�9f�C�U��=]g��l������*���k�Ҩu�!�6�Z&s��'la�D-�,Ò<���� �ZS��,jT�ܱ[������/��؊�v<黧הI{�7:*"���[�z�̗��Z�����guN;�!��딽 	�]������UJ�G�޵�F8ɬYp]�
|�K?��`J�6O��PEU�3���G��H�Ë��~v����7�ˍ9�Y���ߚ�jC�9Tش���{��&yh�ކB�'�t5q�ZWg0 s�Z%��ΛE'bn��� ֒x���vo�X��y��v|��R�D\���֬�[ye�>�W������ ��d �3*�3ޓ�0�T6��j^�8���(��jg�\����M�Y��j?8�)s�Z7>BY|� ��W�_����'|H�� ~3��[�:u��$F�ŖL��jb�c_�&Cx��OV#��ǆ�T�ީ���#���bY�5x�[ߎz3�!�3"�
�̥wk�D8�����h�;8�$�T�%�L���}n�+z.�n��us
Guh�cLYш0��ڈ���e�]��d�@��������*F+���E����Sgn9]�>Lu�%��4$ :c�<��&��9��^{$-�KѸ؅�M.��f���Gۈa:{��ޖ�1����UC?��g���Kܔ"�4��&AZЃV�ٗ�T*��h�((���.� a���O߮"6����}?�N�lخ�7�6�Ig?-�p�U"�܆%=�����̗����/?�*� ����<0tf�(�6����!�~��G�����|�<r�5P]Z�
.����nS�Y�ٱ��$\�����D�n��QWXg:؛�w�C�Ut�0�-�Gd3�2P���~��&"��N���;mL!��kq�������Q�|��(@+4!�#'�
be��Ig7,�s$e�؜q"c��*� .S?�o���M\s��P����s�*F�;� �H@�~u�
�j��Si�i|������٤	u�BƝ�<`�3�	a�{gz')��2����}�@L5��!�����rI�8:���,&��k�V�r��h�����q�����rs4>T���o�V0	Яc�Oٶ$�-�K�+5�*w/G���e�5(�Js�sK�Iq�D������oA���'�ϽgivQ���G��r�b�Q�󇧤�޲�'�1�!��o+֥�I�Ϧ��w��oH�2g�|�s�hIr�/h۩�t�2��u��;t�V3(,m���Ӱ��8�}5�e8LB���|�}8�o����4�ߟl����m�Di��`j�[$;۪�#+Q_��X���l���b���ZW�	p�= �G�e��L�W�-rlpY�wj����,����/���T��V��Ծ��3kd���\�C�A%v�q]����8�_��Q��|n�|��&'�B-��?v �&��t�⑯� ,Z�!�Y�2�����`2b��H��֟�#�Zv�lʔ(w�*�q���	�l�=�4��emgh4nKR1Eg�@/f���H��܊�AK�����ӹ�IJ���'Ï:�ID��"i���}1�� �s-�s0>�H�T������^�%�=�*���^i{B�+�V�֦���]P�S��(sKV5�A��(	N���gE�Fn2L�~$(^kD�&k6ӎ�Xlʾ6`��~f����.֑��?�_$����+產fx�u`��jA��^���R��ќR���&ci��s[*IE���mc�l��(0�6Pd��C��G!y���!�9��PR�Q�\u�I0#+y��ֈz���
>Y����O��@��u9�Y�۠�H&���j/��^�l�-aAG��\�����`�7�
<��b\\��`f���,Zj=:]�5x,S�����k7�?���&Nσ"��y!���0�zI�7[��E��ڈ� %n[�UĔ��d������e]|��Rg���,�Rrů����isYx�"н	��F�̽!%~٧���4�ޭ�:M�w��9���E/p���ahY��.���,�C1h�j�O�G��̢�?6�I����&5E���Q:/�Wm���zJ�����h�7L�3F��
8�5l��m_��������y���#���(��Yն��1bth/��n��)K�O��nX����H�o�N�qJ׵�L@e�쇍uQ�|@��c��;�	�+�'���(9�3�&$��
�����{̜���7�m{����Z{/����o�T������lo>�=���-�@A����r�%���c���#���xM<4����M-?V��7�O_ֺwʩI{)��j��VFQ�A,��"8Er���п�D�be��Q�S�to���ϱLӑ���,_�=�,W��!�J�\�b%ޑ��y�>����E�M�%��ɧ����2��qR+�|�`���"c��7	���:q/G��G.فaP�p�Ϭ�V�QmVϟ�#�����1;�?<�5�|ۧ���E�"zMs0��H��}�.�t#.ҍ�$�efE��Dm5ş,�2Nm��Pe�`nK����o1��ãWƝS΁B�c�̩��m�)Me1��
��4�u4 ��G�}��ݧ�-�rCѻ�,�.q�$�%��	r|�N�S`��La�G�k}���V��]`JG�t��T�Ч�F�7��ZF�@"�v���#�=-m���+VԎ��[ٱ�s�B��Y03ap`�D��~��?$���{����V�Ndrø�u�3)Prly�|����Ac�܌	D[UK����
��d7�6�CDʞ�970�IB`�U��C�� !3�1�^�+�O�Y3���r��P2[��g�A�=��N��t������ַ��Q�C��~��\K�/x9�pt�������YL�#x���� �燒0�i�uۘZB1@̸���@����ި�$C�*H@@i>�[к���w˸fݼ>Ր��F�}G��W��>�B�vK%Ж�m� �v���0�Ч�f�sn�^�v%�����~�@����<�ɆT��Z��\�:C4vm-�6��F�J��n�Z�I���!�W�>eU�WT|;'�ނ6<�P�/z+"��t1/>�,����ٛ�̯�[d�7)=��?��u\�;�k�j&L���{��Bnǣ�<�AW4�Ŧ�����ϱ����_]""N'[Wv�@�գ�O�Ł1e�#�|o��~[;_�@�+�s$��"j�EJ��(�?C7D����h�S��\�x�H���/l{��>6��E0���w-���z��<��pXag�����u��W� i�)*�Ud%��<*'�~���|�}�*����>	n�t��Q{���<�����$�t��{2�w+��0=xT	�As���ȟŘTT�e�H"����%>ճr�w�|!�xZ��۱�6)�E�-���+G �_�+F�%�QmQ�.
�є�F�1������\;C"�^�$�U'�eՆ���(ؼ(��{�����CRg����~x�6
��6&Y��y���4K������d�&��}�"c86�&j�g2N@-�K>~G�Q#�Z4	d�l�v�� �V���ʎ{s�q�"L�34_��G�B��_-�꒯J)�� �A���+\$%W�ְF\x0��N�{��=P)$���mcOg,��I�
�	e=�\ 9^�V�dR:zeVv�[�y&;�f����2h^�\�i�M�j�ۡ�eQST��gha�!��$���1���Xܪj���r��9˟�Z����~��;I�$��4[Z��pQ�վ�.����=����̿j�j�]��g�I�3�"���i���V�K2n�BԐ�ST�u&[�Uf�a��l�(��ΆcɊ_�=��lK��|S�X��>8����mF����lM�\%+�E��m�ܒLsG:_��
�J�<�o�$1h^� �h� ��_��X0y�.�Kt�-�v'�t2H��i-�8���8���݌@b��"(s����M��":r�KFC��!��O[3��V�����y���}��mzl#|���:���hScM��F�e�������	<��ދ>|�����hG*ucDFD�gSܗ���߸�c���Ϲ��n�ܥ�ø�\�^S�AC��xDʈ*�O�h�CaPC�|��(�Yan�^��)CXu�bL��!�s�W���~��+�l\�&,���2b�A]G�)8*-�FF������5ǿ^��� ]ү��ݮ��?n8�����_#|��>�IJ�=0IX01'V�mA�XWg,D���`a�p��k��ܜ�\���{���|EN�R��?�:�%�B}�5LR���;���A���R�W�eGdeHɖ�5���Z@eΓG,���]��\ѐʚW��N�{|��'��/������(O�>б��i��?_��B0W��C�vs�l���m�Zr&��YG�Qe�#�AJZ�ᤧg�uCZ��Έ˹[���L���3E��YCѿ���k��*IyA�cqr8 �	�(��v�RS)��/w�3ԯ��_!5H(y�$���3F��$O4�y�c����t��Z���?p�[�9O&۰u�����n?;(�BS$���׫ԓ��,�:���b73��pN�92Tv��c����z�O��G������upN�NQ���*�����л�v��Α�# *NQ=��@N��h��a�(�Hh�?�|�=�LJ� _l����O����t���R�r6QH�N��7���)Kǆ�:"/~o/�;pE�O���B
F�b��4�Ou.v��ǻ1ܔz`w;��_��L�svY[Q��y]!�o����2cJSa�n�\��t�2EK_޾�~�-���r�2���0+�|lE����,K�B���k���5�I� 8�f�?nX����+�k�1��Ď7�q�̆�>�� ���QAM�m�C��L�L1ڪ�.��AN����D�ǀ��}/�a?5E������"�e��ܫ}T��(�l�}:�)��1FM�d9v��2yA�z��D?�i�/!��U3��̟��2��ֈ���"il��D���܌��,%����~A����2��#)W�!�.B5���"�	�;�c���fHa�I��"��w]}���/e[���߂WRB��6,慈4����p���� �dĶW5�EXrЫj��-��jom�K���N�ɣ�0'�����9�c]�*k�"�����m]�t,9� �8�Z�|�7�h�V��#��Y�~%���\��*�b��E�o����u@!�P(���7(M�Ҁ 
a�gD����9xyp	5����N5=��i��J��{��3��ez��2@p\�G�0{��=����Z��=,���|_��R�i��6���,1slc*1���Q��a�Q�����F�ѓ��E4_����P�]��i�����&�K��T(�xUU~���m�&��P�w����F
�� �3�n��#����h!�7�{�r�X�e5�/����j�y��l2��XZ�8<�-\E�f61�"z�<?6nXl;p~I����\i1q�%�h'�Ia7��8�h�;م�k�C^�F;)�X������� ݇*�A@u�o�¾O�6Y�=����]�p9`��>�T�ᢊ���Cs�7nS?gO��t�E/R���ȵ��;i�4���N6)e����,9�oc�d���̀ �A�ץ���I�&h,�Q��Z��NJr!�é~z$h֊��� ���#�&���[s���\���K� ��q<�� TB��7;��(�_ag���w�^�Mx!�"5.�P�E�	�H2�s�Qwxp��>�4�9���(נ"�̃C2���_i��^ �9�pѪ`m��ِ%�����;�y����,e����\����J6�iM��"� P�Ī?&Z
���X�Hu���v�b^��4��dAls��� ��s��&*�0��>����HY�ڳ� #h��ś=�z/����=���N0\�!� ǧ�=�>�tl�W
E��TN�q�������&�*jbp-���|�Ʋȑ��^H=#���۽�����=���=��qZlW�-{���	� ԍ�!XL�'g�l�z��p�Blx��S����JqM�=[1pϑ�%�O��\jނ��@ޏh��lz�n�!���Zr`8(�'�=}�U%U� �����6���3^��,��^W_���J��V������+�>��!�:���I��ݓ��p�>���l��g���'	�3Gd�%�D�OZۈK��V�Pf��p�ї+�JbK0��������;wj�<��1��E0jT�����(�weB$���KzQqu���x�e�2+g�����H\뭻�v6�]��:)�T�$�+��,3���`V.FsnI�⧨=���_=%L!
.�88k1��㳯�N�5���t�;�ؕdW}�s30@��etD�L�� �`��좬�<;a��7���(�}���T�D�sZ� �1!� �z�x(M��e{�Pf\�ǟ����Y��$cT�DFnӠޟ���������i��`?I'���4>v~�����SN|�N� 7VY8��%м�R��4iy������I�^��'*}���u�V~�������ή�MC��P���@Q�5��IЦ��f���e��j\0*U!ѹ8وxI��82ES"i�t-Ǉ{����Z�r�K�<�^�)gm������7��@� ���T�`��k��.�����J�G���T1U��)jݛ��K�Օ�} ��1���h���Y�=)x��)�VAq����ӈ��cd\Y�8�ba���l�mR�T!�=L��M�|7��
ߘ��-ntP~"7E��/�	G(�5��J񝱇�E�aX��Y-ANw1�l2��3�f���o��T�z��%/�45���H�o3�Bi1����d��W���9���'���U��3�@���4�gҮ����|[�Y0 �}���<MPOK]Nﻺ��X�LM�f�������!&f:vH[,��M�=It�x��m�9�������<�a2�~Nj�\*���ǭ��|��Z$���F�����}���.븍p��S�D�"n_��C�sЉ��/N��Ŏ�D�[���-�	��#�	�W(�B����^U�3����4�Ӻ�:��$��>��~���8��ԟ%�>�7o]e�.S�Y�؋��J�`=ߞv��q�(���ZpP�)��vǫEa�TMGc��O���5e��PF���V$FN�9d��� I:��ܒ­�0W&�GB�`�X�܇K��N��f'�pǋR�D��^�-uJ_�S0��+�Iɮ�d�
8�(� ���V��1<3��>����|�k/����x,��Գǂ�uw���>��|��,R��1L����̃M�&��$��f:�A�H4?d�jH뵆zA1D���!,ľl7Cd�
@��uz��P���2��\o�)6��	|�2me�o���=���'k?�;f�rN��T�[�JĹ�)@��>��b�W��3>�=�ML%q��R�sW7�VNt,�8�~hw��Z��4g�T22�)�Ds)Du=Q����w�r��D��e�r{<���'C����b��OO�q�ͦ���ѿ��p�{(`#,FԄ��j�r�<�}/�Q���B��+�Fy!s�u�&�3!+8�(����u�i�\�~� �)�L}TN�g6�A'M�3�]����雡�[�Ȫ����I�JBrH�ȤF���@��c~�62���H"��
����h.͝�>��{��؇��G�ި^|���]x���t�� -^�����d�?���f��[ȭ�hp>��_�:��J/�"��G��(��<��Y����V�̺�ͱ{H�L��J��4��g�!��7yc@B8�����s�~�|W���� 	�U��D���3�㢴�է�t���7#�q,����MJ�'�sbh��j���؄���t��gB.�+�!o�1Q����Th��*��TP�vX.��<��`�:��"���⫷��Ĩ��%��j�&��L\_��Y�%�H�#!a�=Z+u��/2wOe+��:�F�]FC-�� ӱ2c�▷s�o�%�o��Rd`&YU�[ɦY/���E���1���s�r�������ʻU��=�C��_ܘ�0�}r��]�<�;y�$����e�#n�6� �������(���x�H)��45� l��I\4�Y�i�*&��ikY�A���Ӹ�	[����ƾ�ė��~�̷~�k:,� �Hޓ��>�(�cM?�����J"����Hw�B�!���8}�J���7�h/��e)��W�^oH{6���Ak0����ݐ�ބ�R���_s�U����AOM��ߋ;�@>1잔�k�w�t�\%z�>�w�q����&D�(PT0D��//��Ew=ʣ&f��O6�E���"�w#�#ì�
�]�RU���ۋ�a����@�
	,S���E�)_��o3��W�e�����Y�Fz���l�wDO� S-se����~0����w��y3��[�>n�8<�Ԇ��V~^(���V��G�>���[Mdc�%��9Rsn��A�}���qkq���r��Ӌ~Γ�������z�As�nb�)G
�j_�
��(�&Ͳ��������ң��ӆ3����]3V��Z+w��$+�c���xi�3_{�@j^�U�+�S�L w#&�6�ĭr�"1~�]�t��+e#������Jta�4i~zRi�60��	 �vW��(5	�E	v���/Y�D,�?�>y��^p��+�"�59g�w��@h��5;�<ܐ����-+1��_�a:1�7[H�)��	4�b���H���D�4)B��bA�	p�]w,%N�����@B94�4s	�t7�;������
�ݥ�f�h-�i_{��ŧ.B(!X�����
9����p���k�u�xp��ebЅW����>P���AD�1Χ�:'B�B��l�
�3~s{�@����+(~���_}�	�L����iv�謧.��[���wԳVżY�	�H����ڻK�}�K]wH�j�[I�ަẒo�2>�0+�9o&��Rq��$�p���8Qx�yR���u�s�XR��6������1m�h��G��\D�rџi��t����ˑ*��g,nv��j���5"��#�j�(#t�#U����db@�4�=%��@B��(���)�L��Rۏ!���@�8NF����Jg��*���x��N�&�S��:����A���Ҡ��Dm�% ���R,�H��d~I&�h��/�+�7�>{��-?���vJ��	�!N��,�ӓ a�t4��r�ʜ*��<Ps }�c�eW���L
��L�L�ͷO��}�nX+��ԉq�A��o~�m]�P7��_�h�E���r|�9;	R�-�z��R%杳�x�{�&?��>����.����_��������Z��F�_�-�)H�M�,�p&#c�!��c�{��d8m��l���s��O���j���?�m%y��כ*���R�IO,�\KU�GV�md�ؒe9{���.k��Sdj�-0���������=��d�_�}��%�p�ҭ��:� �3�7�n�YuR�����N��f��+������)|5�ë���~��|a֬��?��8|�~'����=�V���F�8LCp&<)� �%֖�a$�w�q1K.�������s�Y��'룻ᰈ����}��^�JV��(�78owZ����#��?��Vsdp���k��dܝ���~m�%u��`�=��O��n}0�р�Z���W���C�
t�/BS}���w�Q8a�.?*ښ��;Hj�H��<�6)�bd`�!q[/xsv�iD7ٯ}�"�9�K1���!\�l�Ů�N�tV�r?H�Y��VNř���`�]�E�+��<Y�1"��ltg_�h)w�xF��@�k��.1#X\'67�x��#]4�������^���G��X�H�u�]f�@B��v�j3_����H��,��-��.��dI
����+���ڍ�P}�Zp���RTE���lh��i�G�I�o�Nq��p~w�$R�Yy��i����@:d)���@r��^7_l;�����oO�I�@":�#��H�BE���pQ��|f��dϙ�}�m�����r'��o�ɑ�b<��To�ߠ)2�����(�{}�Rz����J�J��Xh)qS�t����e�I��Af��k�^e�	�����_�t@)��(��l�pMD���ػ�z��J�YB��`e�'�!f~�s.8;/1��]�&Z����K	�U�F�v]޹!z�M`Z�3��VUe�o`31kTf�x��S!u�ɟ�"! "�]%�镄����.��Srp{���E��=4���t����u����U@[4Г|�<:!H��I�O��f��xwD�\9M����4�����D�DDKԈ^�}K+�|,C}@�j��˄Q�H�6K�ҢgX��kd!g��lJ�K�<a�|��^Q*������]�N��l\}`U	�����y�T��ܯ���f�$Ԓ�-��gs[OX��eW�;�;�$������MϪ� 5c�ƖH���>6����I$���`y����߱���̺X �� ޯ�X��Cf�C��V�'l�g�tBa��܊��=0T�f���I�y����h>MDi�����޻[������`�.�ؕv��U!��	��5���L���9�-�x��~��ײ¹���ETF�B�1)�W]"(�4�NJaF^o�E��`�f�b��seR�/������?�!|�{)ᯀ��k����	���Aq��R�N�|��WpC0��`��x���J�Y���yWZ�P�;�I7iu ��p�I�&7����G���A!x��r��3�/�%x=fu<z���*��*H<�2��#�gGxаR�x2�����|m=ˇxx�gNg���,���m|L���t�έK�j�O�t/����fN���D�+���w�Mz���ٞ���[8B��ć{����o�2�sG)$��T8��;%�������s�c�V� q# }�ߩ���F�m!#��`a0tػ0ȥ38�����"m��&rX���^t�L:�`������6]ڃ�N�H���o�g�MzQ�X�gX�
0��t��L�cY1�{Ez��'U���ZH��\3�7�h�9�| 	�d$�o����W#�*������V"+^�||��1����E{'�/|�]�Y,��Y��p��U��{}Vx(o~_�T�>2�MR�Ȁe���>�S�hQ���
	hz��Ȫ��6�-��no�ſ�6%H
a��UuD�����v�H��~��з��-�N��s��GM��ɓ�Cy>�@���oTcُ�L���\�)ٙ���^�[�t��d�0�4�Fg:&䔫tN�k�Zy0��,������I&������f&_ֈ_h`�Kw\ ��n��3��KSy*��<He�?��V �Za�ẅ́R`��I�t�*�3c#�LO� ��^Y���sw w��ד1c6U�`���~��c�3��B_�^�ŏ(l�}r"|,�(`ۗL�rQ�Eϗ��Z�K1<v���K5�Y�}Z�X�-ߍ��9���p�ݮU��� >�&��TR�D�+E؇z�U�s��2�����`[2 ��KjxQ3m�d,�����t�� �m��=Z�6�Jr��,�hh�o��z����R)Q�z��f`������m�]@
����~b1��76XQ��)�Pý x���<�ⲛ7����Q��1ü�,&$"���-�f�o��C^��f��X��h�Rا�Ǥcn��(���4�%r��Ew[N%����eH���h�̎��x7�O���G5m�%"%�ڻ��澏A��~�brI��D�wp�"���7H��p��˔kR~�X�z���6^�>F��۰�+$r���ꆓM�>ok�#N�ð�8��f�ٵ��@W��(�`���W�{ C���V��]��v�������O)�Y�eQ�4:��T���l��	�pv�X�hݑ_.fk�B"���Z�:5����y���F��'w+K%�c� gK�R<Ǹ_Z��h�P��7�큫b�^pBK��(�4�&�-��˭�=�ci������G���y��i�l�����Y��S�5%5�wpW��]�'���d$�J/�9y�y�$������m�����d��ӭ�S=����uJ�k�Z��F�ݓG]5䧏�g���.0\���:��7˒rC� <Vˏ��~�446�"���W�ӰA�`�e�'P��ⴅ�����J��a�1 �{8��$���0�&󔬻���3a+��C����kМdf\܀��\+zC	����	���B���c%Ms�mAl��.E{�
�U��=�K]�P��y�ӎni�h�r���(�O[#ߢק�*�F���$Wp�▬�~<=���[ �{���kH K!}H��-��'R�ߵ$m�ݧ6��zj�e:���,%ٹ��*`��d�̆�+s0ݮ���4=�. ����pLS����,��`�苐�[���V����u+3��t&��B�����������O���d��`��柤�<f�Ƽ�C�P���*�V4���T��E�|��d&�����r9��&	X��.�W���q�a0O[���r$����H����SX}Ta��@ڍ�L��|���Si�.�߼�?�8���r��&��i�+S���;�ߺL�>�`_zI��Jh���*G&�qZ\�	��dt����(V��s����Y����7y�ȅ�n!r�ZL�K��j��5I�͊��5�},�SX(*�V���2����K�4�ͽp��S]Z�V�"��t~���E��|�C�*��;|f����F�&g�ߍv �EԂ�� �%��;�YD�1�}�&hO�V %��owzc�F���Q,��aB�0��4&ԏ�_l�5�����#�(�DZ/kx�UwEva�����m��+�(�hڱ�~���������-��i����i�ƃ�W ��	t�5㎳�@v�V�������1n,��r��!Ό-�6���a#�ᑒI���|@��To9(��Mt�$}� K�k �2�I��Mn�[�,��/Ƶ+�o��b�Y��X�W�i+�h|�s�D�R�K��#I~N��(��������;�)�8
�G�-�4���i�|t4�wu�]����`��<�Nr�� ��h��=ר2��)��1{2���_y+M�`���(b������N�Oyy��T�F�T2e��T.��&�OLϩ�7�g�3�]8�c�G[�a�g���p���)[��A��x�jj��)V���5T���[�qæ-S��X���S%�u�tݭ,ؒ�(t|���g�ՆlD_�l2�g�}���Co��z)B�c�5���F?�D���S"�
��"m�c�����|�QN��3f�
]T8��z��bq�`��0�(?5ċ#`��f�)��Bs�8�����������I�^!��ە�^YXI֒�My%fD�}qF�rc�'���8����5��G`�%D/w��X�v��,�z�)�^��WvC��r;�����a�9�g7�c�*D��@����aF�'��YP�E~��65��O����v.�Q�)�� {L�T�-$�);��;���Ȭ/��"/�urɋl3i��:�|F g��d�cIz!�_���*�W��Z�V%4d�/p�.�3r����Vj��^�Iq"p�X��/���{hE��۬�����\M�,�	� +W��O	".:ے'e��T|OK�;[J8�q�b�:g�@�#6����a��;%�U�e�ā�����T�m���e�!�K)�>�ƍ-ld�h`E�:�D|� ���pT���6��#'i�Qo���N�6|ƉP��C�#���1+���mx��u��8H�&ù��U�4��<6��I%����,KB�����o�~x��s/<����\�Uv��
zDjǒS@�.\7ϟ�M�}e ���l(`�!ڋ�-��m�j��-�v�^X�6��H���$f�}�q�9�
�}"W:�k�Ehzb�He�����?������H+'X{;�A�������U֏q�bh��Q��"ZB&�h���A>W��4oM���CC�](��}�Ԕ�W�Ԩ���Ol�/yr�p޼��n0�Q�PRS�p�#�UEh,6W~���'ya˜�)&���Zl7���9�E��^Pѥ:�����$58�-\�V⾘i��
u���ל��mD�d��V�]tC"���wm�W{r����h�fO����̐��{`�f���@,�
k����~U�T�b#�Z��"?8��p�+w�	a�A��{���%���%�4�@�詫-a�-�Z)�z�!��z���F��P�!`�-˟@#�J@�zP0Z�����\Ψ�����Խ1"!(��>=�A�d�����G���ڳ��Q�Ϡ@�ҸI�
:X��PiEgw�Ѵ�!V�	�G�,Xtг�5�k��q؎xd �h��)_W�g2�����rP~E�H�ę�Ur-4���|�w�T͚ͭC;D��Wzr��3ͥzԵ\�O�w!���,vo~&%�{,S��Q�\]�d�!ɪ%WOi���bj����,����d�Bq�'�-ހ���7���3�O��'1-u��1�c+|��~0�.G*R�Zi�y�i'Ƈl�1rS �����
��>3ö���i#�@�R�w�G�́,�́��G:ѫ
��S)h #d� �|+)�0�O]��+�a�f����7sW�Ԏ����3�hZ�;ؤ�߷�d�%���1ĽbM#���u|�؉n|RJ(��W�5���D�8�of�$�&�n�ʦ�uv崎z�Eq��\A�eN�MG�{���s{����,�4 B<
N�>s=M0�"�m�]�ӛ!A�\?�i{A��$U��v��fnP����ċxT;`A�
�h���h����6�f�����Qs��}�o��6�=�6i��X]�;f�u��!0�刚'*�'��u>���V�a3W:d�Uf�������R��y��5�����&�N՚�A�]@�ߠ��"`_�A����z�uB?��ǫ<f<;%7�S�݉؂�چ%�����b
f����c��a�g-.�)^�l�u�J@���8Zf��QCP�4*��~"c0G�Cдy�T��[뫡��2��aӍ������㷀��a�y��N�f�/�'�ޟ�� ��2�Ӳ�t��>>%�5�^>�i����dL�#_�S���h��lqS�8��X������ �zf���1j'��2(�0/�?�7��QKR�̓Hw�Å�K��3Cȁ�f�<�rS���$�^��<�!7&e��ɔqa��L��UR󙩢߂���]�7�������%�:��[x� <K@�SXW�����-k#x��W&6�����2]`�AI�u���;SRo�<Η�'�3������
�x��&��gm_�g��nM�o6YF5��+�[���G�м���1*� �,x�e��@�+W� N����.n$Άӭ�t(=[
�w¼�!�kn�?�pA􀵇��ZY��+EN�OUW�`<�;-�����<���s�1S~�u�vr�<���+��"�{ĸ���hf��!ۑÚ;������A\c-$��Z��ѱ����N�E��^5DhV����$��F7��1=,�>Αu����w�ͱ�>�Z,�D�i�k�Xo+�,
_����`{����5U�����,ܔи�/�4'eR�:ͷ��3!!��eL�t��MD���=�v���A&s�>���q��
J����}��ƚ�n����]f���WVRF��D/�ђM�˝q@v�?�9��pD�E���S@�U�o�],�*���S��	J����v���N�#��g��'\k�0��Mz����
�FB�V{�*ʜLR2u+�
�+��xT���5���qA�E�`	��Q��St���c��@#ɸ�e�3�[�=�]�N[�fI� O�ǔ܅�+73w���܌�t����h'�\�]������[�eP׫g��s�3o�0�2������u�t���Jϭ[�,��U?W��t���cVx<.��с4���*!����r���{�IoIƉ��m�̸s�G����]Ckl徳��@�����Q�A��{�v:no߂��{R����¡����'�ʣ{���Z;Ew �]
���5F��G	�wD��Rp8��jw��d���7��Mj�j�3�)D7���?���v(��e\�`XUU@��}�@\*�i�c��A�9jY�,D�zn���MG¯㢖�˷488AeU�q�;��Hϼ?bjr�Ta0lmtU�a��./�}�2�f����N��Ổ�zDn�6Ю�H��O	TǜN�<�j,vT��a!o��sV#l~['�{�E�N��.���r��~j�z��Ƶݰ��T��"��4uҕ�n8����������X��`%�+F��MC],+�|P��6'�|�5n�.�,R��
1a���x*O�[;�z����k��rá�݃uG�����B�˾U�:˺����y4l�����:�����ڗG�V �fJr|j��?8#��o��2�*O��]Ƽ`:��tg���{���͗������c�����dï����h�\"��9�&O�L�(�nh��q9 �M�D��E$�i8�̰��V :�U��ݚ�;���|.���In���C��5��p +�`E�1{J�-�� =zw��9^x�`_ͭA��������:�<�Sp�9�Ҹ�M%����I�16o�c�/�ʱ-p��#�L�΋��ȐG�T[Hc7���|������$��?uBT��5�ٗ���)4�:J�q�Y�O/���c9�m�?�>�1/���EIW35�Ei!.:bI�gs/O�B��VR��i^�/Ã?�\/-��f��z^�i����@^�%k�N�HM��)��D�QW�d:}�	ds�9�5� M/,�	��8�8@�BЬ�_е
V��-Y��FV2x��\���� N}�G�?O�2���逺�(��0 �&Y��^೵��˾���@�0�'�<O���J�s�+[��t>ɱ0���2����9�ݟrm�[�x���35.���h���ɖ�3��Flns<ۑ45��auѿO�0�����o,Z��Ua6S��wGh�jK���;�"\��^t�e��#o""���>Iy��AsJxO����(3�m��ć�ha��]&M1a����_�x��}+��A�0>�[�m����d���?zZ^�Q��j�o�J;� V�G����[�s߀|>Z�P�H�N��?� ���ʶ��bv|m'���J��<�M�m�3�mr��g�����P}�$ �'B��^;1D#L��|�jwl�"f�۔�X! ��C��ӂ�F���_}��v{g�k!�ju���	��\���+��;�(�>[�N�������M��B�N�l*$12hB7(�ք���9J�����َL'��a�r�M�6�C����I���6�L �y�����!����q��^Jz���#`Q{	sԱQW=�G#��|�k��1AU��=(�ͣ;�I�i���u��J s�ٹ�S�E$H��1�B�s�+4�U8꣡�[�d�'���M��y������`y̖G%�?�:��I��}�uJl�v����y�6�d�dH�0O�/�1J�2duc�⌙Z���jnH��B��'7t�N�:�����U��W.�;��( ?�g�TVŎI0Da�ߣ'�'?{0�0/A��a�FX��9������u�6�jN����~sq�E�1T�`R>���U���M!ե�W��'b�k�6a�����:%�:%,8P�'*��� ���$-���m�]�;:=m*Q9�'jL�B������wa�o�zz:ҵ����i$|��;������YH^B{���olMAW;V�\b7D8�E�Y��o�PFZ�k�h�S"X��O]���[W����b�^Х�iz��K2��ֆ����u���(���.5%Qp�;�TDᒊ�n ��jg�i�^��5?��sF��P9e�.Kľ�	3)��m�ƅxh����z2�J�}�"�]7����!�N�O��66�~��	4��H��o~p� ��.N�7uutC��0T-��"F����(Q� �'��B4T:'��� X��������3����ޠ$H�Bz0`�\�b��h,@�S��O~�m�
52�����R^0q�C���`~�N�,�*�6N&�'�L3[m�C4AiƌeO��aNsD<Q��槽%��q��Q5+�Y	@��SBs����_���z�~�Ώ,\��?)k[Ʒ���C��S��h�*��F���e+,t��ptn�����mY=�aj1�cy�=|�;�AO:IaJ�z��
·�%�T�1�7��%��í��o ri�E���8��y�q����QJ�^�5ś>��~�~�Q���~</��$Ֆ$~��aC%�Ő��QWc|�ٝ9t���ߗ���^x�u�5���X��rJ2L�05�PE���U���)��z��Pc�-Nc��a*��X����3���w��X�X�[�hf3��Q���+g#�]�un��A��B����؂�H��w��s���m����Z/��:E�_�Ht�A7��mMY�!���@����db�,��̰���9�N�[\8�͵]��s�a� ��u���B#&�0LQ��r��i��VLo��ڙ�7��9��@��;�눰5n�c�#2�%�K	K��k7���:+�EB��3�V��;��Ei����Z�/�.�M{�������͑�nL򹒙9�N��]I>!�u���
WQK+ā��.�\�a�a<�,(��9G݂���Ft��NwI����q���\1����8cV4��)"C�������x�t���k�5�*�Kr~�x���}��s�1	,�	u5p,T�xC�2�r��k_p�f�"]	�*���k)N1����UF��d
�\{V�c|�wq����\�M�3%�չ����Е+�7��3��=����D�慀P��ܫ��	���1CD�d���34�]6��Y0�Gm�����ny����{��hV�ݻ�b6��Pq&�\�G�	c��GF�m����D�oc탘x_��F� ���u�	eK��(s������K.�6�����J�O뇲X��#뤩���A�/m(w��A�?�#<� �2��$6E'Y����o~P��o���	����A�ǔ&O��AM��N��1�$=�CB��1{0j?|S����XRDw��/䶮<x�e*�|������	[o�?��n���%�YnH���3�j�3��p�T����	�~��Z(��e؄��A����<��e}�]��JX��� �M�+
�"k�yמ��MvT��M�Q�Ő��6{��\��*�a�\�4�!�qӆܞ�?6�CU=���g<��7 �D�l�����Q7po���(�5�ő���!$\(�SGF�
���+xJ��:|�$_Z�WW/�)y��$�.%���6d���eBȤ43%��M=#�h<��I}"�4~�:y�z�=R�V�pNIR�X9~n,]�%=L��yt�^�2���p��]�f�B�ж��q�:��}n<����Zi�qPj�^������tRY���gT|(}�k�^�Yq�t���a�G� 4�W��}
W��BV��1M�(j���@�
7oi���	j�i�!uep>��ڤ�$�쥊�+o�%v��]�$��'T�gS�'GVG�	����0��b(��Q�{"�O(��_�)
��J�]\?]A���,�䣠c�a	�>�\>�Y����*/������̘�3�Y���?�6I>��/*eV�tI0�9y���4�"[���>�[�7�mc:U��+��"�C�6�+�u-���fbk:��¤nG�Y�.������/'�"l�,e-�蠠Ǎ�XzWKY����?��kȬ�AI���t,I+K`����"b��
�&���u�X��������S�� 
OY���tE��=�y�Z�����qR��#�t�M��������\��`s�s�b���'������Egz۬:(}}b��S�=b��q�Ia�M��݅�·g�=2�-W�j����������s�߁�RY(��lS(M%	+S���+"�RG���/	^��i�k���3~�1�&��:���^K��e!�����9�{�ǘ�jI�e�>�����kB{�h����7Ďa��n���� w@X�q��)��O�g��v�u��d�����˅R�w�>ޯ^���_<����?�o����+�9���_K<�� �Xb�,��d��BO亞��ǳ�+	Ћjӓ�g�)���o��]����3M�8��l'���R�T?o��o�3���{�I��F>�!3���P�dΟ>b��܄MΠ�4D��n�A��@�h.��9�%
��I�re�41bk�� ��e�\,��Yy��x����V�P�n� ��l��\u��j��m�A���y���i�ت$��۝�:�?�B5TO�0f5+����k�L��n7.�"~��jT�YEI���}��3�mk^�=���f���@'��H�����U,%'$�K����K�>�Uu���S������@o�i�_�1��W�?*����6�U���sK�v'Dvh͏G�6 �<-��0�Q�81N~b/�^]>a�fK`Բ4����5C����*f����]1f�VRj�N�q���b(�c�Kd�ǜ���Q���:�036��6�$f�W���)�`$��u���^�P�!;vOD�MS�������`�c�"�����%�i���B�<5{|Z�T��C�B���P� ��D�n������"�]ߜ;k��P���R?ѩ�x�sQ��mCu����"a��&L|ʈY"�G�-h���g��F��o��&�"(E�T����Z�d�ۭC�z�D��Ѐ��-.���U!Sհ�]��6A�.�6%̟��T�����.�B}���ȅ���i�O�~ռ��R�f���0�h�X�LUF�Gi�x�5��@>MUf���.�� ������)���ދ3\�~��D��%�R�J�$�����5ߖ��ߵ�s�e��ԃ��c���6:��uɥ֖�e$z��a�*}��I�iӲ��L=T3�D>�Gyl���\�
�9�FA�u�4��>�̃c����)� ���SXL�3)��R�t�FC�܈ �5]4�Q���t����
ֽq	�?�f��V崟�|����,1�A��Q�l�Hք�U��5���t#�%3v:����˺]�ܒ�]�c���{��;"v>�}�|��y	Q7�Q��,^��SC��&�����ۓ���a�3���0�'Ia��&Q��v|(9^`jY�Yֿ����q�x���w%[ĿwIp�����Ab�����b̉�9��F��kד+�oPҘ��"����Y� ��^S�Xyǎ����mٞ��\��m�a]c\��I,k�1�a;ͦ�B�%H2�<�����X5���b.[՜��B!	�����$OU��X�������c7ݼ��)�ȆO�� X��v#�]��������� ^ ��k}��$�$���>t���xRk��Hݣ͵r�����Hy�	V�FV�H)�R"J�y�x�G�S��]h\Q^��1�K�nC�`���j#3+2�R��h������~R-'���=_�T�n����_�O�6����-Ja��t𝆒��_u��m������ ��ǡ21x�Ӻh�#�RX�����j�U�Onq���GH�g�:p���L��Ή��(�M1�9����>b�A��B)�lP���S�u�����	[|QlՁ{�A-���m�k�D��;e"��k���*��޿AD�kN�t�Z�����3�o\J{=S#��B��e�d�2���x��㞴�ƅU�ܞ���8a�ˠSCN{�IU�E3�ա�r5`g��)�^�,N��3c��Z�_�\M��c��ƅ�P�q $��f�;yx&��_�?�gZ��6�bx�pg�(�$��z3�&��� 6�-�+h�G�sz��nl�,� V��Zż�o/'`p�f�K?\�ߏLW���O� �T��ņ��7�AҒ}��-����A �ܢ�ev�-�<��́�6Aʞ;U���ʿ��0jt��YI�����9�nL�	"Cj�H�#A_Ƥb�i����s�[N;���Am3i�:'+�gy����"�%��[�ӏ��_�;=&'�X�yQ)��y:��k��}Ҋ�3hw�7�|.���)hԇu8"�]Ÿ��ml3񓠭`���ևa��@�h]�q����� #�j����2vwG���[�`�I��WU�r���t�����l)ܕ�E��e�(4c/۹߹�^xe��9L�`ꈧ�.�.��m��
��9�ވ�:��&�m����!o �e���.1�CJ|:���ӻ_fv���!m�a"A��؅�!ك����`���\{��~N#���XY�P�Yma���6���G&7��=馗�hm<����@�T� b)eO~kR�'����J�Y'i�}\�:���]"uڞ����R2����iBC�X���F?5Z�U�X���O�?-Y�
�ђ2��s���BMu��b��7�d�����5d#D�K�m�|{-}.p6�R�E�^Na��ݵjD�Q��[���T���|(7��PݤZ��9�5��ϕٌb:�!Aw�
-I5~���.�G�L�ͮԧ��䆭���R���8|񯱑�rL��%�&�E4?��Tv��ƍ�Q�v�ӄx���
����Ɂ�ǵ3��U���f�O�DxZm�u<b�>4L>�N�!/���p��着y;�X7�=P����d~��(�b<]6��f;�c�sұ���'�;��+Ƃ�"��7��E�`���Q]^sr�+�V��Y�����Ū=�5S�_�҆��f��I�3�wD��TQuh��&�#���A�>I��T[��\gln�y���]sv_W�I�7�c�h�|�����-�6�W^�u�`�6����Ǫ�������^�m�Z��~�t�L-��%������Dt�����"H�ӻD5��3�we=�����H�b��b�[;$D�j�g�|���*�.x�f�@�B��W4��,�����u��[��i����~��ê��/��`��_y`�8X�	-�����@��Ah�cFa�a���� �*4T:��v1*�� xD_�~�c��c��U-X��^�F�4M��jբ�>ZEm��>��+�N��^��	�'���[�X!�sP�\4� p(@��.E>�9\  �s`�����ԍ�T�\���0���_r��0�4�a�v���y)���3����V�m���?���EE�i�!g��C�ϫ������w���� UY�R;�W����O����4f����j�]0����o��,g����O�&�2VF3'�"���#%��.��h|�M��}H�/ok�H�(���gBg�}��}ћ��IFa�cl�$�;�����whR�D���$�?[���H����8��|��c;����Kf��3T��n՘� �����&��Im��9�v�O��T�����+��e���fjڪ��7�:yᰂd�g��J+���ll{Pu�tQ��jd�(�kgS�XJi3+��2��N:�\�E	?+��,�G����{��p|�(f�,"EUf���ahkj�B1�Ժ��6l�},n�T��M��kKK����n(s=˅�e�.�C��wp	�����ss��m���&��R:O>���6�s�$@O(�-o�oެ�����G�}������°�-�9B�������w�;�@���Gۢ��.�I�7������Ad?���8��4��g����2���-�]��\7��<��^��ݛ�L5������� �8���=U�`�;J��$���m��*e�ҟ3q������b�/��fc����7L���~N���TpT�"f�J�gA+Qg� {_�Cm�v�ŒJ������=.[�H� &&t��s��om� 2c�%�k] `��@�>2�ϝ(�������$}�NK�_t�!��<3ۈz?��;H��봼.}�|̢\�Y���8�T���x�(N �:��fI;,d����d]�O1J��9Y�8��먔���\��-d�~Y|�?E��Y�~�qޅ5��U� �c�7�yk7�zL#�ry*`RmB��Yf��ײ�ZCַc�:��7۰$lK�-I˥�5��y�w�vR��G���!�����TN�w{q�?��][���h�{���y��)C�laGn8S�S��8�kt�G&֛�^"YW��/$mh�8/ ��׋S���#��-��}���!t�:	�-���7O�h�����m��F���(�Q�dخJ7�w<�V>!��6N�6�����G|?� HC�p�����7�2 �M{��Pd���h��<�	���yF�H�%B�j��S�03X�܆f�����ĩ.?N��V�%^�=�������v9Xb��%�E7�A���G,��K3�L��Ї�]O��:-�K��~(�+�=C*_}������5!�Վ��q�LOY�`�R�K%C��'�Zk$% ��i�H5O�M���?@֚�7X����y��"����S.�]�o��:}�=���Z�����hg�D>�3���{���FsY�䢥rML��Q��w�d��K�D�[�wvЍ-�"�V<���~����1���ʽ�.C�5z54�Α�ؤX�3�ƢaS���>�'���#���~���Cl8jɄ&Qn��勝n�i7�00�_k|1I}rr���vq뎈�S�uFVC��q�� �y1^���.<����rB�dړ��d̄�4�o_� M�<���(�Ey.�E���L���P��])VŬ-{0���Fe�_�
����Ϋ|@�=�Ħ���a����E�*�qp8���}B������G�u����]B���+�;Tv&�P0�9�`��[�#���X�,�]�?�s��ȍJ��;~n@�Շٯ��}���H�ڪ� �>&|=��*|�V�ex���w| �s`z#J`�.m(�	�8A�|$.js�RW�xy`-9>�cq�g�O?ǧ|Qۥ�tk�i�2�F�1;��^,�r���A"�EH佌86�.&�!V��֙>�I[�\�����6�����8�bl�N��y�cw,�" H��y$���e�5�P�S��UJ���yy+Nx�ԛ�3��l�&E��I}�C�M,/���#vG��͡�{3��z�B7�6Df��ڑ�3H�:����Z�rz��[	�G� -��"W���]�e�cF���3)j��+Z�v¥��LawZ9�b<���&PB_�U����p�x�22[�̟β�2��?d��a����{2�b7>ڃ�=�L�Lu�dʓ�
��4��4��Gؾ�`�s��{�𢲖�~���X�'߁�%B���2�����H��]Biء�����a����@b�GSb����j�dX49���8��	4Yɚ�r�F���`��|n�
���V9�o�<۳A|ĸX{:D�m1����}V��a�z���8T_�G����Z��8  dyz �7)u	n�C=������J^j������Ez�.�)��x������ri]Φliw<kxX�4b��1�]�s�y�j�2����`ɥK���ji�u�3��Q�-��[�κ�q��,����0i�G�UQj�� E��}��:�����xf��*-�ʶ��=�,�b���j���)��d� �d+�Ų}�+K*Т[����Wpҵ�#<(���m�L���&ʧdm=�e`�8"����gM��x��J���F��,���KQ�	�{$������iV��~
�2>I�)�����td�Z�\H��I�ٔ�ݨa( �*J���7��1�S kBCGgET&�POI��I�Ί�=c����*#�%�<\���|�
���On+���%�`_R���T �z$&��E5�������7�5��0�C��CE�v����=�=���l#�&|3��K��'��(��H��ǳ▮p�i �zx�h��i����մ�%h����g�b��)Πwߑ�PGysw��Y��|��
S����5�{�<�y���wu�3�'�C���ݘy�-xq��W��4'{�2��x0��l�NU&L�g������G�2�b�_��V��}ژÅ���qi�U�A�
�YRjl]�~8���G4�6�������$���s��i(
���f@�D���� �^�lo�J�NAg�h�����-w�Rp��U�6롢Ef���4I���۩C���t3%�M*��]�r}`N3��cH��'�eL$xsu��C^�G]��UؓfkVU��(ө�Vՙ�9�׼��HM���qY���p��2r aTbJU�r{���7~�O6���I�.���	"_R�B��Jއ.��{�A@�/mT# �nFB���B5[=�� k� �f\��Wes
�w�e�B�~�G�M$^�L^������㓴�� =2_|��0����Tm{cU�5�v�F�1�(c�;)U�f���`���8�5������*�f��t�EE-J��p�x�B��}�c�s��7^�Z����;B/��H�4�1ݖY��ﭶN!
y�U�b&��a�����aU^�q���\�mg�%h
���1n��� ��퉋������*�M^��Q��y�)`T�Y������T���Zgv��[��r��W?�Ǻ.�|�P�Tj�;q=�&�5��d.�:<��mߛ;4"y0J�9��b�Br/z���J["!ÖEOZ�䶧A����Yc�x�{+@�P}Z�k���
����N(���$�)����Z{Z�>��FL�E��c��n��2.���Y�(����Ŗa�Sa:�`ɻUc���w��T�U�"q�
��Z+`���A�&��c�s�z�QF|M۱�}͏쿜�r\AJa��8�T���u�I�ڀ�5?�$��OS��� ����e�c�<AМ��y�|��p�V��4����Ad��K�=��	�2��8�z��*�U�J��	PH^LEL�N�Ҭ�R���ڳ���X�����xd�,J���A��P0B��-���a�E��?W�h�tW�]����!(�2�oU��Q�ǈ�}t��(� �E<���7�O�		4���s�j�Yxx+Hu5S$�)�
K��'M��֬AB���*����^�(Nu};��.?��7�5�������)5_{3v��K��RxI�ȴ�sw̑`�����<�e�J��L�����	X�����x�L��35^5&n�11�zw�>�n��ZP.�@�̋K�� �IN��շ��H�͍��~���F3���
>�`,E���Q���F���$k�צ������4� ���Hn��:�f���,�`���[9�>�Ⱦ�*1��N#y��VO��y��k3O�=�=ï|�)��9�6pRƫ���%��u�=��8�����V������'�T)Ϛ��'-�0DH��ZS���#���D����RU��;��jç�?�r�0DZȒ�j��%���F��}Ƚ7ٕgGj$M�m�pجu	��M.(��%�ׯi^ֆR�+�' y�+�9���\E�À�&�z�E8�N�nV����֛;��� >�U����M�!��HS+���w�������;����F@~���+���W�YQ�r-�,�w0k�5�uL��<��ۃUoȾ�����~�����x�[!�
1���:�zCRa�
�NhpkR�ôs��W���G�ي���x�� 5�d�ي�1��8Qc�5۸-��s��l�B��8-oS���Z��Ǯݕ�~�E�l�Q��}�R9*e�H�?��N"E�����w�t�aG��!Ix~���p{�p�`�l:Rz0�_v���
�����:�eպ:_��ٓ�����8�z}��S����P������h��s�x�'��}��(�U(��;f���r`���ғ��B�F�ɺ�]�p��&�V��&����{(����Ё��k�y;�+܇؅�L�r8v����� %�G��9&��#�dK����n�o].j�8�}>$OM2uJ�(�D!��f�4����9����{�/�x�5t��/N��rJ�w�j�e���ՂIyQg�5㻊Q�ri8Fu��/�*�2�S����
]׎uluA��_��
L�����F������x�h|h��"j��u�@Ω
�ľ%^�34�?���̠Ud�G����Vʞ���u�j�t"a��ߡLb�C����{��D���W��M
�$�e5v}��Th������w7�+���?|����NڌQ�luM����6;$�S�rR�Xg��g��7�R���@��
�� 	�!ȕz�h�f�@���S�:D
����Z�O�U��%�C��0'D"@�G�+k�����񈾣�`������!+nj�A�A���F`��+\6��8'�I%i�L���ȡ�$��U���$4b�?�A6�i��n]ckϩ������{�\��ތf��O[��%�a~$�e������E��5B�� �E�Z�#�B�����]��r��e8+A�Z}b� �D�@��{S#��~ VDQ :�,��6��D��0D�$g,x�Z�[/��G�Ni%Hh8�:�e,Q����y#"��Q��!>��[ 8�|sQ��Qy�C7TRj0(C0:"Wgўb��Q�q$�Wb)��F5����Ų� 9,��}Q�n"�m�a/��5l��+Ø�0�Ǯ���lV�		�'��=��s@洳݅�ц�R|;Eal0�I�QԱ�J�}���UژD�$��΄V�6�	(;��P6B��&h,�-�R?�J*;>cAQb#�V��㟌��2�������~��J?[����CQV0�
�~���S3
�¾�Пlv!��O���Y!�ۨH@����:-RMO�zE�`:`1୨�'IH����1��;s%-.	 nM��ە���O���7�`���yV�Wk�[�hx�� �l��n����=+�^��⺃���y�1�qV�u��vr�ȧ��<~o�%itche�'��'�x�Ӑ�+4 ���O�����E�����ի��
2�~XeP�_��n��0���8�޵�lY��v-G�MF�q��h	K�8a�10�]�l`�K�ot�O��W���F�k�7V�k�O�;�t�zb�|�X~�0�1"f�b)�K���X)����%ʁ �uB|B�ӡ�c���R�HW��~kGt93�� T��^kre�L�~����n��x7�Y����0O4���}xr�����ta�|%��w3]_�'Ns��H��b.N��L��f��n3���n{8�Aib�*�4�*�z��&n���2�"m7.�3H��םɊj�dY6	n�V��n \��n��w#9_�D��J[ajIp��q�ْ�|ڢaGjͼe5t����@)�u��{unL�d8���ԃ�6J�0����q1ک�֧�8�6u<ӠW�,�-_�дU��E�ۂ����K!�.��� ��
�d����ѩ��f4IC�2�t���0&�Y\s�,�c�*<��u խ	� �h�^w���,��9E��$�+�
YNM��2�H�LS��փ�ס=JNɖmfI1<�j
>)��ց���o�Y8\g��|�gm���='�WJ�DIsĘռЄ=p��%߽�w��ρ{/�w���6 ��T�i����D�6q*�E�S�����'$?�n����$��R���Zf���1�(Y��=L�cq�C@f5f!zt�<�G���J�Ţ˓���Cgc	�|�R�7ߢ��Y(l;�;���W�S�rg�h X7��[����zE"Ӑ��_S�q�h��0�!T&�0�2�&xR�ɸd*�q���B�����iSh!Lv)��|)��6��1!
��
��t��*�Z�ja����ؤ�<{��X~����������ț8��w1מ��L��?R���ʪ]��q�{���w����"�a���Ƕ��4��?�:2|���@||��Ҝ%���08�V���o�XBd���� ў~���ت���a5��#�O{�Ԉ�H�� ��5ρ�2�-�UAZ��39�HS���Rb��RJ�	XZ�=j?��/�H/�]�q/���M��Ug_���X�����X,��f����3�L��`��Rq6� �v��lzY ߽o��ۣ?�G��܄����E��!�l?%�I�y�d=�i!�oQ�&����q&=u�e�j�F���� C�ѥCN�>Ѓ��B��7&�T�/�i���zw)6p��R�T)4�w�/��3�z��C4�b��5 U��-��yG��6��Th}�)�b������kBw��kB\A 7ʣ��D�PUT�OLe�s7[�'��\��f)X���E�:yu�-lX��ak���/hT�v�&�х-��Eα�ʋ�M�r��&E�k�qf#�4��.��jx�M����W��M���Q}�=B��R+��������y�x�����A.n��GI���cŹ�M��:d�m��zB�n�~)���{F>�(�Z���;���h����-�W���T��5_���yn.Dk,�܈��	C��PqOuH$�Ds?�O��Ϣ�Y��?V+�8�+��L�,���FEF�s8�y3��\�'<�q��|Q}v�Z���CQ<<��.�i�J2���?��Mf]n[{�j�+��D/W�;E_�aq��(�v�Ӛ:�LG��0���]�aG�L�j[�m�%-#��ש��xܦvD�0��V|Ǣ�%vy�r�����wu}���N�njA��k��B�f?fk(���N2vk���y
�r	�)t,|Fm{U M'����?I�DI,��ʴ���mG�ڠ�� ����O�v��o%�KP��pD}�[Ა��kx����3���j�|�$���?J�v�}��)N-Nu�$�C��� <z��[q�n;C�����u�\qD��R����S�xw-���޺��y�ڜ�W�Sc_xH�}������ksd!��s4����c�Aʓh�s�Pf1����ySzA% �������~��X݄���c�x4G��`(�1���@�_�������ɝV�-m5��"����_K����K��3��k������l	5���}�K�uc`�6� e�u�x�v���$X8\�u����[)w�5�t�����~��`���. �e�&޻�������n�����2?���ARѣ�A���ч��)Ƭ_���.b��D7�"{�)t��ȻM~��g�G��B�Ѱ���1%nR{�28��U�2�ވ�f[��%��m��)��U�J�b�2 <q.<���'_NM�=�#f���1� �e�.!,�^�����4����� ͥ����/��^���t���<��˘`ᬬ3[m�jh�K.7/��t�w����b�U�="fo ��H�L8W�y�>��Z�3r���� a��gbTe�59Ҫ��'��<�̢�'�+�N'wA� ���o ����x���z",˜�C��3$ip*4��2�؟`\C���ϥSj�D�P�sJ�uʣ�lI���w6����j%]@
/�#	[i��j�Ѵc�i-�N�j*�)�G�1��m;�%�R,T��X�E�d�8��z���C��L��W�x�LF=����������!�&B�y��"������Y�Q+Gఋ<��o�(�>���� 珓r�o(�sG6j�3H9O%g ��(0�y��Y����FKd	��Z��ߵL�
t�D��!��f�W�i�:c�;On]$�)a�������e�S���悅ڝ�WW�-�sR�H<Q+E.���HpGmH��1xdDWf��q~��;�����Ő���J^�� �f�I?��4���O~��M[����O�_��x'��|+	��o@Bs�i�ݗHiUF���Mx��N~`���^�L"c����7b9C��~���C{��\�o�Ȕ}
� ���j-��g}N+*I֝����Ě����Ѻ� C�j��|+�kꈻ%͇1��ǵ\�ƱHb�n�̋w�:y���n*���W~�0U�9����q|���ʜ���Z>�f�5\ªPǶ��Jqc�a�D�܊����t�M�} �V�v ���"��AP*�y��-BW����^�h[��N6���VpN��k��Q`�6Π�z���
�%W��_c$��T�>Ǿ�s��::�\���������-�\/�ȭDN�ԏ��%�>0?gJz:��o��ed��է�q�0��2�LL�����w�U��Nx����\iK{�*zv��t*���7b�ˬR��)E�k��S�m�N�m��6��Z�+Y�1�Ah��yw}��_��#X�ɐO٩/���ϝ�);儲��Z�T��k�#�&��+'�6�W���[�ij�l�Yee�*5�֩��c�+���hI5�\=ݑ%��Q��x�w��!�P���ݩ�'y��5r�I��7�c��O�P���i��J[�����!�9��9c*��$	��ۘz�������~�>:&,�G�V�K�^_���-}f9��|j;�L�����*5��4�zJ��L��}�>��J@�b�x#D�׀e�2�F��`��@vw>f����^�:D�
t�TZ���Cʵ�������w�'����WJo�f�N�j�����d��z��N����l����mjC8�;����H6E�02HQ�S�B�3���Q�!�Gy�����H%W\\�W���s^�,bLiC�
������m�4�[wv�;�2/1�r�5�b���[�woTʔ �*~@�sy�̭򥝞b+F��
��?Ǡ������y�o��ᦶ�������l�$x9���6	Qa�By��Mς�u��x�G�+���<Od؜��>U�2�g�rf�bm���a	)�/��Z,fT��*s�������`�_��C��^���ݫ'V�X��߰&ʘ�+J;餃!�Q�O{�&�,�	z��V��6`�y��s!�T¸'���0݌fh��m4*�5���?��C5X��1�Ƙ' M���BX���}�?]l73�N?���.zL�U?�u#�.~~dHَ��=��ə�l%ܱD���g�<!�w)�*@R V%� ��Od��I�[��;�͛L7�z�L�vu�j�t�5,���������6$�j��w��[L��=�-(�g�	���րW�+��a�MW��f-�@�k ���9��I4D��
Dդ�UY״�e�u%�%\��O`������P[���2*����ޗ(�G��َ����G��Ȱ�D�}m@�a�Y١��S��%2D��R�?mʞ��Wb>�vW6J�����}���C�k�]���d�p���cwo��_�^x�PFy�o%H��P�ru��>/Q�B������t����V�� �R��wt;�������IfK�*)���0���p��,��Y��T��j��yB�J�R�E��>��{:S�������F�Hs��/�w�Pˉ���U��S|刿��?b:F�d���%�b����C��PvL�2^��/�&��])�AV�>�_K�S򚗨�G���v`Q�3��q�K��j��tQ���w�����ڊP|�z������-�!��v����L8K/[�;��tR�	jV}S㯳��dp{�v�ѡS�����ٯ�����	�bml��<���+T���l3�[?`��������[��4��/y�/=Hp�D'a޴4m� ֊4`u���TK@��U퀄[���$��ب�x~����͍�  ��\{7N�4��VU'X��p�KYy=X������Y�F��e�K'"RE��Gz !�����:�_N�K���Xͼ?������Bv�N�+
�Ui�q���	�U�p�=x`�9X,� ��p&2���Ҏ���n���jc�wi��j��@^�4��&�%J����E ���%�+>�M@�.Vt~���X�v��bd�Aж�Y.4j<.� 7�*�\u8Z����*�e͝�I��[��O,@1k,��m�^h�v�ȋ_׬�E����Z���M	������鰝��.�\�2fe�`a5�u���U6���,ˉ������'���M8��Q���o�zJ�lѕ��E�D`��z�g��Ё��qZYߏ!=ڪO�X3�L� ��\x�q,�U�3�'I�'�E��7��e}�#�(3�#SmNj`���k5��I0��0Z?��V�N�T!�q65|�_�l~���7|�6H1{��x��?������j�T�!�>���+�	��q�U�Rk���q��������U? ��z���yJ��_cmY(ѩ��e�j����Ǵ�sD�AI^��s�/�=V�	@���o�z�<
�'�;$����*��4Hf����ڨ_1A�V�#��O�$\�?����w_��ݳ�1E���|���/��gT�OՈX�<��66P
[ �"cUYc���nhg���B�]p#�/�U*�P4
�`&G�@\�� I�s��=ڹ�n�gS�~��K-���p���P"�o�la��D�N�������p�Q�6~Ϡ��J�k��z�@�yv!'��)��{�5'� .��X���5fU�`P��ZMMӈPå�rK�[��
�������j�b�����0�R��*!Y8�����!4��=�?�?Ψ���Px��������iA��X[e*V9Wo��yO�+)�S�z���)	�w�ۼ�F!�;�6Ǹ ȟ�W����Z�ש�*Y�%�w�ɑ�<'�t��/6��Z���m;�@!��'�]>�]��-�\��5��8n�":D���n?��`I_��Ѵ� TћN3��*��QÂR%o�4�b>�>�LBN�ц��P\N�c��J7ɾ������ެkO㖋�﵌���s��\��sݡ���Or���0-i�&�P�����Acc\my�VM����E�v�<��>T���ZَE���BcqO�e��(A�d����ɹ�Ji��04\�i	WꎩV���u��c[��V�9����?q�c!�Q�	�z�E�w����Vt���;�d��Df++�Gz����"ﴡ��_��T�j�:Hޖ��O�@+�	��`ݳfP��$�����b �v�H�E�~odeOմ���g�?k�t��́P�a�������eƉ$�A��0�DX���c��p>)ǵi�a�hx����cxI���$��2�BN�t��~	m�	�s�y����"��F�ɜ�9����?"�����>HG[��&��i�ʤLQ�E�����;�]lub��z*�S��A!��ud�a1�U6i1ߦ��ۅ�s���IGH.��������� ����Gb>'�a\G��>̾���p��Z[ȽP����X����я�t�B�ϵ��[�T���`u���� 
��"����p�\W{�����92	O5���� �m ����TAo�!�>���
��v2/���Κt@�"��ސ�9�f���9!k5����=U�G4HeE����C����4���l�l0�)T�=*C���V��� ��5ס�(�y�x�^ҏ��!S|9b�*t4�ӫ0�	��WƝ�L��,m�}�}��=͒\L�₂Q��e4�ګ鵓,gQ��M�O'ӣK�Rus�>������8<�.>��a�<��� Of}�5[�ku�FB�9E-���@Tv�u��#�:��,Thu���܂�}���Y2��S��s�$��\4��ɝ��8T�dKIҰW<�C���剹�$�*<U���p��7]m�.'dn�k����~z���[�.H�*�>0�*�A�t��9��#E�p�S�tԑ\!���L��%���0w��+����5c�2�j^I�|��`����y?���_�E-@��OՆ��� �GO��#�pi��;/���rZQN��鐢i�M�7[�=�*�5`���ZM3-�`���G�B�".J砎6tF_�t�j�z�_��!�	����0�珙����Rc�V�@v��.�T4�ii��&��>�3_��>G�硐X��>��:7w��J}��E��A�_N�ԳtFe�m���G�"��S�?�Ru����A���x0�mu��^ C�׫jP�y��/����V*�]�|�35�����߯0��G��f	�J� ��i���iYda�j0�s������Ĭ}~���
�&P\&��Y��X�����/8���������ZY��'x��i��T]Z�]���z�x)P��2� �@�-/��>6&ؕ �.��}j�lMvɄ2�4�F���I�QK�C�<btM�Ya���-�Q{�������ro����Q^>
�u�BC�AU��9I�-+��M��ݬ��A�8r�w�BZ^v��\�:]��Cڒ���]�B *o��}3h��W�+�������~�1%��l{�ǅ\��Iy��B#�ӄ`�����Z�6=��m�r�W�Ӓ���������@|y�.#4����jz��[����M{ �î5�0���0��	U|��r#���D�}f��]��(�H�Kwt�f��U����f�	#��Ө�e��f�<պ�6��������!��h�Q���=XK�L^��<�����,oE���_f�4��Nf��M��I?�1f�S�8�גN�g���iB_k`1	�Ɔ���"sK|	bG�*#Kp���f�۹* ���˕)�g�%&P!@Ɋ�?�I<�C�x+��H��i�a�67�Cp�$@A��z(4�;��jTr�4��T����ks�3�*���q�p�X�,&+˞Z�i��_(�u��p�iC���.pz&T�u��~9%�<�Ć �	>��+U��j� ���=j�H5[
�x�|��b&�)D�2��I��G�.�́6�()&?}k{�@�PC��v�t=��?� �P]�#�B�B���0La�a�k_*�,V��:�F=v�<-MF�R��R3嶿��P�qLP�4|�����{�LpR�'#^0	2�s~\s�a�#�ѫN�z�֎P��(������,p�à`�Y9�Xt��/�L��e#�@���mp�%�8S'h�4-V�����d^R��y/�I�D;H/"'"cM���l$P}��=�͛{�f�Y>��R|v�
��*�'�p�mP3=�m��^�=�N���Aw��T�E;���$z�~N�F5�'3͜�B$����"�!��*�_��9��fJog
%-ׂ�������?q�I{�L(�9g��߄}�y����U�eĖ�R�[]�r�	_&������[&�&�Jh�Г�I8M�cÁ�YcGm��(m�u�xe�����gp�?F��j��I�)�I9�h}���������6	�}��Ѩ�j��u�^�a�oӻ��ջ�ά8co��)SGht����VюԤ?��yh��TH��.|L��%�'�O(ͪ�g�[nb���<�-qyKQ%Lj]��q��l�LL2�Gn8p��ޡ_A_�p �=�"�z�QY0��l������E�x �=)����,F�㚘����#��R�+��E ��st�=���?���f_qb�g��RrV��qBp��{q<0_\f�R�4Z�XK6}�[�X�0;�}{1�ō0B}���2�QIArD8�x� ac;o:��,o�(�i�	��\:
��Ĉ���s���V���>Ar'*pM1 "�b��nH�_�_r�h% �oHR454\ivZ�ԫH	��^EpE=E
�2z�6��j�~��Ӓ�_a�M)��ӢD$o}�g}�����!/�eb�!^!퓜ǤƑ3D�2���;n����]���[�>���	V&뫲cIK|���Sj+����5Nz9[3 I%%t�l�@�1�.�,]�W`����|z*�H�F6�tZ��a�LM��ed���]չ׺Hj�Z�9��ˬ��͌um�V��d��A`r�s������R˷��7�
�R�=����+�d�Ym��v#��������'k����!���[x���i��<�uq=-��eՖk�9,�{�*���^���)��0m7l��i�$��y®�M� �,��]�=���I�;�4[Y�MJ��{��A�?���e�J��J�/�����qVU�*
�#Grƾ���x4>yl�3'�{O����y!��
K�.����t�����(N���W;�#i<mH�K��<�u��zOЮ�˨�����֥cq÷�'r��m�H�MJ��e�\OrnvǺk�k�>�GҞ5K�+,qB�qz��Qf����1��`�-�<�q,��4�Te9-��&6q�sa%���,��f�VT4�KB4�!��">%�%�#��Ʈ�\�#O25#�/7*	�V�����1i�+��kZ�*���y!Hi�{��0�|�*�U#�JMa߫R&�p�Ei�<�\�PU̿��紥��3W7S������S�`�c��"����e������sn̲�4�� �/ �t�ǫ�}#lMs�g%��V�ؐ�(��Ό֏���X��Y�9��X��K'w�yd�)Ɔz+����JN'�p��Na�3D�+k#�V�:��SI�������c-Ė�CB��؀�v���ZJ�2Y>7� � ���ͷ���cA����&����e���d��N���D(j�'I��F*ԟj�ķCS�S�n$ov���dn�h_�?/b\c�Ak�"I�Hq*Z6���L��= �]�0�ӦG�/M��u�U낵��"��l��wlA~����M�`<W9	%�CjSl����(&Dҧ��e��V#@�эv�-1����&��dM�=^ob�C�*�4϶;#'�4t�җ�����0{���Z��E����?y�[��0,�X���k�;��C��[��a,P� JE������s�����H�_�B%U.B�4'N :�Q��h�"��pM�K�p?�m�K�q9<s�̖��n�Xgj��W]��V]�fKW�<a�`��a3\\�T4١p�A���(2�_iˏ�u
)�Ny�q�4~��{��O3��s������b�������O��m�
nH�ʗ���/k/���1J���.�"�u�}{} 2�/V)�T�����ߏ�^�I�&בD&.�[1�O��0w!�f��$��N違�D�T�} `��wiSG��.]~@�(��¶�/Lit�U�#x�1��4���u3�;�:;"�h�fI��*�I��qX��#�4�e�v�T�]�����@a�m��Z��Ci6��u���o�\ⲓ�bmDr5:y�F�4��3IxV��) 3ڸ��������'I&8�o�N��H�؛�7v�T�����iߚ|B���+{A�X ��bjU�!�?�퓓�p�MT%�����z �aj7�-��ЙQ�B/�j#߾���<�)��â	,��0�.�ގ߆�x�G��h��dt	؅� A_C�\*�%�E�%4�VM`�	� tU��?�Lϻ��zL�e���L�EMn�1���5�Ӭ�z�l|\�j��Ux��H� �ْ�L����.댢�h���N�si�F��ʬ�"T4���^��'��2r{�#db�x�f�&|WM��p��O��J���AM���!�����c���܍�78IL+�(������������Ph�ޒ�6���/���`�2��,- ��;���xw�V�/BF��mR3J����#x�/�����<?K3��ɃT�WK�/��H5j�`�Ê��B���e<g3���)��|�Ddc1e1��
R{R#����^��t�i/]�>U�lS���]�ܸ�V����E�kW�ִ���)5K,,������n��h@Zh��uY%v���i��	�J}_vߟ�&PFt\�����;%��t�>��A�Q	Л���G⏁R���{�0�h�#�0bf��0H	 ���%X�,�X�\��L�D�B�oS�5�.DM(��j�U͇6�Gj���q:�]�J̧�� �{�"�����[�g�`��9�MBo-v�H�z���4��}'&V� )��	ܹLI�T��3�ɗ'�$���Ľ�1��CI#b�θ��
V��I�O���Ȣs}��mDv�2�3G�AHr�1��c(�۞7��v��������'MK��0椹�G�Zc� ��򮱚�eA䘥4���)0r�xk���vKs+����m�Tº���LkE>���U�;g�o�����]o��-��M�v�o���o��պ��4������W�t�B�M���E�wTN�V�ڣfV7�j��cqL! ���D{y__	�/c�鉙"�����nXB���݆�i��V���8�č]�}͚��q�k�,V˷n��w5��
� ������f�^	�(�(�c1�c��i@�We�]V����H�[������7?�A�ψ�o�Up�ml	3j����I�xv����J��I|0�ϋ�<n�W�Ht΋��^�A��ڠ�U7�~A�<D��$xU�C���!�7m��s����x���C�ի�m˙e�b �ڦ����I֋�*U$�S�f?���LLˉ˟6���l׿��N� �Z-'s�7H�F���f�#�a�b�X��8���2X���w��ɜ�"����u��?��+�5���V#l��s;{�6��Q��e��r:����!Z���z�b�֩}���n�o4�'�t	�	Ö����6&�}��'���atl\M|9�yb����&sp�,!���1[ԣ7&�"h�e2�[Mo����\��ǿ ��so�@�Z�̉����l�l����
kk���������������!W�G���p��_F���������$��OS�4ї�e	�@WHv���1�]��.�l.�+����k�`2�[Fq#E��K��\-�1C�X�����ay�<ED�eU��n¡�p? ,�@:��Y�uQ{��f�:���iޚ����j�?o
�3�Pz����.<���a����bzMw�!/i�:�~� H��(f��X%@�Z/�/Ѣ��L��7��H���:�*P:�;�
� 4p��#A�w�>C�f�/f����߃Ï2�f�6}�c�$���jce^G����=y�&�_dt��b�����)� �;暌g姨c��Ő�2��q���c�Vh�$K��-�+s�	���>�f�U�ǀk�=^��3f"J��Ǝ�d�#���ّ����i21{��e*���=ٲ�n�!�Qq�Wnb�m�	�y�� �s��7�;\�GjnR^#�[! �(�r�2��]��bQ�k6U�j�=M���,1#w�kK�YV+�Ly�iNO���'���@��Lب�`��J�8�Ybm�'� A�J}�2��AP�?��o�W@��,��z{���4���еhmd��i�d�NA��� �%0�ꙕ��Zy4�!�^lj�M?w�WEbZ�hiG^��-�{"��g�-�:"���z���`�<G?������鎲���(�	&���?�rTR�B��S�CJ[-��+���%�a,�c4�� �D��[Ey �j���{I;t{ۇ�N���~N����Q������π��cR��[�.]<�$��|��{^���h$���8�!.�8��-	X57ٓ��\J��h��'ϒ~ƅ���F�82KAF8Aq�&t7ӡ����U�!�f���I�C9"m��KU���"2hU�	�C���*�K��q��m��1?-��X�8����~�@��14���W����ke>[��܅�4)����Xvi���O��h)yE�p�<��ĩ��x�+����y/�ՁUc����g�tcLW�r�2��#i\���'�o�v�),�ufma	<�f$4/��I�������n���;���iyBpB�J_I\�J�v�QX�_��P�x�o��x��ػ&��
 -�o�w�	����G��xg�y����),�!��� �l��0�5@�`FTq�|�9�9	c �Йj�!qq�=��~G�j�Oo��O`�8����쒕�q2���qC ����a7�1C[	%��r{p3v��#A1��g��1�:3��&��{ݦ3���kVP�f71"���O����k��z����f���3�&}�&��AeO��^(mc�?�J�;Zx���G���uػ$j�	��z&U�K��=�:��4N]��\OnE(�+�d�pP��������x9�vӟ����=+�*u�����8����5A�����u@�'.���js�&u��SY��Y_*��]i��0�jj�j�Z~��H���#P[��]$�`�!,�%�L9b�D�L���љ�7~s�`�g�@?���M�|;���ϧ�`_(+��ˆsm(����"f9�5�)�ӪX0�$�2�ni��)Y�=Y�F���j!v&�o6�n�`�t`�
q9�D���n�5�\�d Ș�2�C�����7��w$��L�L�3���dι�̑�E8o��\�������2�uco� e@&?i���?PH��b�qP���9qo){6�0զ�H���ý\D;�E������bÎ�U�2m�st�!�z��%���F�QB��S� �YT�'��[�c��9�\}�z�A��!�����������pN�{C�qൊ6�Ȣ��.�i�n���J�_��\�	qs���`ϝ�HAԡB,63�)�~G�+��o�M�9�6e6�a��#oH]O�*U�@U �����v��}J�I��ӵP�l98 �]��/�L&
��\��U��P�L4�+�s�9R%9�6���Imd�
��л�(�F�8E�ΕK�{VG	��䥻��@?��
�+QUV��| ���?-eg��yW$����^i��UC~#���"��w؍�� �3�K�R&$�O���g��\9t11�R�d��"͘���&m�W�7Pi�ݖ���R�<���6�T.<��L���6���3�rR�%��|J��(Rvl�Ep�B��Z�(� �r�BK���D���d��;��q/�K�LO�a�Co:�.��P�U�=��ԛ�#��$'� �A �}���t˵��9ˠ�8n/.�K�#c?�6`���*��r�7$�4��@�9	y�U�+H���ڇ9�@�t�sCW�(#g[�X����j쓀N���^�A���X	U0�OS�2�����Yn�����Q���_����(�Z�Y-�-�'f��������@1S��V���u�[H������+ի�Lx��:H�`&��`�ܠE�G���c5_�U���ßi��"��Ԥ�},
����q�v��K`X�R���{����J���gIɬ	}�i|��P�+��_2Fָdeot��n�0Q:`	����^�g�h|��\R2��l\ݧ���2�KT��Є��x$���U+���i\s��vi�r�R���V�-��y���h����~�ן�x��t��g!�ꑞ����Zdv�C1�|	�
���ød#�.���1h=vhW�Њ��X��v�$]d�qA۳
1�w�[l��#W-8\m����>�=��~���|�o2%�O����m���ݬ�,�4�稒��sN,|�5ϑ١Π��i͵���ꮲ:��8�mr��Ğ�g��PY�#�l���_���7��c�2/�p+��X϶�s�V>b��ȳ�Uw�"�7p�����D@<�� �?�O$Z��6���r�����'F"r�$�]�k1���e�@9�7{Ū�?�^�{^as��`2�&c2�. ��nԽ�\�Ȋ~���Jg�Bȍ����d�x��X��tr�2�|�rP#5ɕ��q1�?�Т��g��&��.�}/F�)��b�s�zRx�-r�`���O�y@^���Jh�^U �%�� �!дX4��(�`��cj��ҳ<Ed��B�ҫ�^�i�1A��#�i+^�W�����L��`)��7���"�̊���G������3�k8UR,��*<d���шt�
]�L���1�ڵ��&����q"�0��ͻ�0�@p�ߘ~���%|���k�͘EX��2��>ZRs��q��Rd�t�������i2�E� E���T�XJO�?>�[�����A�S��AK2�e�@�js�I��>)a��]�����R���i	�%�A��H���É�ʦ�F�xo�O�)��m]c��q"�#������E�᫘����P�((0n@w�Cd�Ae!<��Emg���bo�X��ό�e}��DF0<6��oT(��)2l9k_����v*�e'��-�Z߆��(�u���>���vme��W�N;ωע���1�e\+�D8��S��:���XG}��Kr�*jX�.���G���0�����Ȍ/b;Ե#�<��R1��*�:j��B��ą峦4�����܆�>.� �uf�%g�٢�~�,�4v���#oU�L�r����}�4���%#�RY�vj�!�+�-
6f���p�M�3�a���D���A�L�1�؜җ�	U�\km��6�����W:���pP�I���U3���.7d�ok_�L�ɤl��[,$�6'�H���5:;v��r�T�n���,�+��~"�����ux�e�)�lQ�ZuZ�8�y��������(<O-��t�\=2�����}�1x���QM�D	s���C�^&�Hz�2ߗ0�g:�dЂ޹衋-C{�7LNy��VΤz��������F�a�Ƶl���<���d��ӾBoO'�������(�sP�	~����Sp��l��"c ��)�ј"��
]�+���%�鸜>�D�E
�{aY~�1ξ˖���Z�, #	_�;AA���cdY��Y�q{�ֺ�eJ�y��|���	�.]�m�K�펖1�9����T0�����ٕL��@�[ȟ�q� �6��"I��wD����N�D6�zBs�BX�4˯�][��Jz����e�D�s�k�F�?M$������)&H�1�m����R�3i�Y��b����y��]��N���]��E����:�O͔G��������}�IB��&F��D�Q�w���<�*��u�Խ�G�-��K4�DA8�^G�c[(v����;�-/�6��$�2w�(��c~�h�f�V%���;d�FF�٢˛��8װ/Q�%��D��)p��\m>��r_��޵_E|E.6��J-#m��W�D�0zc����}.S������`]"�;)��vٻB���D���8�|��
�������G=#ss�q
Ag�Kr2������C[��VuP �j�.s��<E������E�m�:���B"��%������ȃO�.u�Nx�%L�kU��-���	���?�ؔ�2�H�K�������r�] ]��S]X�Od�P��ȼ���b��x}�K��-��� ��4�)|��܋������ޣ��}pa��;����:~ �����.�inD���.Ĵ���g1@��1jg��8'�鲩K�Nh�BP�v"%)����{�pG���U:�p^Z��]�fUvD}M�6R�x�_w֧qA?���j���3�F�ܸ)8�14�̟��ܐ��ˁrM&G�ûz������ &�Z�$Ue�b6�	�-�c�R�ҭ�C<�<�������5PdjPL�w����`> � &j��"�N�LTVl�}�����{��)����p�Js�����$��J���v�����mm���?��=-��p��o�U|H�j^��WX��mY]4�W|:G��wd廒Y���eD�M���f�;��!����d�՝��~����U��� ��
E
]#�B��������%#A���A,���;a?�H$Z;�ڔ�u�h�[]D�|��2r �Z���E3���SSd%�)��s�1�x5��u�#�S�ժ�ץ�O��0��$E��z?���jy(s.�0�W�����d*V$U���E�6���� ��|�R*|�Qe�`���^x�|��30�ȅZ��3� e� cZФd���at��i��{�z�i��bI�[ceI!�99�0��r7���ZB��lCu��
:�8��bB�e['0 �)ߎ������G�	�ER�zRl���0�Z}M�T��i��_@;R�x������x"1���?�)F��+�W�[�q�*K^a��7�w?mi�=1Ħ8_��h�F���3Z���v@,�pk�I< �lj�}���_�[����O�z}n�9ԯ��@O�W���� �a����El�?�j4��lz]�d:��x�Y�ɣ�������]r/�P��{�����f���\X���`Ew#�w7��B� �%V!��"�M���q<u��5Q!t�&�`�06+�	S�u�!�t*0���{��P�5+��:�4����5/��;<g(�]m�$�|0����D"�� hYL�}g�:�ZתC����j
|�M[����BE��|��Y�1�I����1W(��V+��0�Q7�����6 ���v��E�g��j���AZQ�'�m��7&&�zf�uտ��7E��=�j�~e�d
�b����&���V�os��%�@܋
�y�٩>�i^��n���m��e{4-#Y�� O��5(N���-˚w��i��`ɉ�3�l��F�������g;�N-����g�_ń�p�"u�+�6o�C��.؇�4|�;OP�4.��n��g!��Q�mɁ�5��̳���%zL;��@��]����s�|� }�z�^��]ސd&}�`Ш�ܳn��a������آ��B
��V5������ ����ք�_gI2ж�� ��ם_S� ���lMQ�"��I�Yp�|!h��ƌ��"�{5��y>t��6B�Xh�ְ��r<�Չ�L�Q7]�ݛk6�H}�LO��K� d��.$��6:���d4Xjk77�*����O�w�G��ez���V���(�-���OaZ�z���sի���
x�]u���U�
gT��^�ӽ�A���qIpJ����;��*7/���1f5'>���C��#K�C����k�����/�CY�ǂO���,����T�Z�I��������«������vU|��(�A̮6Z������,'�1,���c(�7�!>*�ܳ-H��^ur�*�I�f��������vE͖9�M��J���>�*3%YHц"�É6+�5�=�Sv$
�:�8&�W��_��
ܜڧ�F�E^���<q�T�e�O���
@ߑeu��9�Ŏ�%����נ1LSx�C��\,C�2�{N��8��'Ȓ���'�J6���1 �;i�#:�5��uMI�}Z;&���zt�\?F��}멁|��̎�%��y�2O�_^�l zUs?q���A�h+�=�ZV6�e-���%��#��Q԰����?
&����)rE�ɡ|��$G���$z�]�Ǒ� UȔ�}��I�&
3�<[�";*9%�yl`��hM�2���d�ߘtO TB[���~]:D��(j�肁�8ZԂU��{�0,��877�!���Dx��>[���!��Kˌ�A��kw=�h ��ר���������/��Ap�r���Mus�۴v,�@M��Tq�3[��,g�<���� �`���6�hN��aj	v�i��ݾ���E��ET�$ס�o�����������Ϗ�W{)0ܖ����`���G� ��[\���!�4m.v�Em�7���^Y��ʎ �E�Ȫu��2��x�Q���6n�(��������R/k�sP�v�[����OT���'V<��Љ���B�`��3�ۢ���iῂD�b�y��wVI��\�/a0%F&,wT2Pa�.�S1=��&&�������V�r�æˀ�-�۹�N�j���9���1-f�tW:��}-���V B2�F_���[XlX U?�m�n-�x0��*O��.�c}M���ob�!�� c�d��RݎOlI�if�<QSM��֧�F���� ߞ���׈o*����g�z��p����1A�������f��M�5ƴs�4GŢH�E�24�cc�\Ͳ<��a�,0��r�Z��lr|}���` /~�X�KAM�£j	��c�#��uCQ;I�y�%�z�ё�K��W�S��?�n��W�4!m��ղT���t��*����n_��@�z��^±�9��H7��ÚP�7���!�J�0�?�D�Җ��z.*e���C���Orr������J��琺�'�#6q�����bV��<�y�Hԫ"���}�ɤD��p1���1�z�����+f/L�U�Q����1뉠���N�ו����B\'jF�=w��9�겷�-v�!V+k�5j�`�����l��'�@�	<�6y�T��X�3v|΢SW�y3+G�����^Q��ͣkvRς��%��j�>��8h������]qO�U)��j6��ʤ#��V�7Vk�ދE������H���Q��>�ҍ �w+@�ȯv�O'E�b�35�r��P�"�2�Xٵ�d̫�Qq.|V'�NL�Χ�<z��Q�<��q��a�:��|I~�[�5U��S\������䩫��_�/iq�n�tg�&!�\|�/��ZN�'s��M$	�g��Ȋ���M�+��eKL�O�]�<�;l�}HAМ�F�=�����)v�_P�h��F8��Ѽ���]ka/���>�4v�@��t�>lUH��_��o9XX�
���� Vl������e,A�w�\UFqX��#�!`��H�v�stlv������g�2 �jү5B_[��S�]�0F~4m�� J�O[M$�]ݧ����$����þ[��G�P��ǐ��5���!�H��R���8��ЧJ�ҵ?��<�1Z}��*�N�<f���T�q�,��|���tjQ�ekR���t�p9Kg�z�>}'�L��酼孉s�G:�4���llz����@%�.���ȷȦ��=w��>v5�z}�L��69>�U)_�fR��rZ4q�1���N��6�-��ą���7�[{B-6M{�����o�����B�X�k�9s�B`�@䰛9R�rc��(����@^��UΆ$���ٹ��}�Kʣ����7x/[<�'��%��	�ŵ�"���V���a�()
���M�D�w~gD!�x�E�Wt�c��L}��D��'��ȔL�n�;n�v���̈́��z�s5"���������b�v�s�yi��L�dO�Na�����H[���Ǽ<�����[��N�ϰ�6 ,�����R<O�+�;eʰ�	>^����|������}X
n}�����[�]l�!T"���C�n�ާ������4'a����k��j8���fB��%H;�l֭���ڰ6�a���Z�(4��Q�4b;�\k9�2���!�#T��0C�����%%U���swr�� 5gY�)y%=��<��H��z�|4�=��i ��Ю��6�?��"r}�Y��7,,%6���tS���M���90fP�愴I�8'�E���'}�&��$R�҂ �!�|�5�1�6��h����G*B�J� ƟYYN��=�U� �V�"Nv�ٺ�_�v^@��~��=<p�y��Ӡ�Ɉz���ϰ��6ˬ5%��NBW��n�r:r�/���s�k�����v�Ch;�	i� �����#J<X�Y��Fk	|�S�3L��/�t��Գ�Ւ��a��0x{>}$��k��xG���+|aR!AH��.9&��(\�.g�^p.bFN�Ë)VQS��b~�P8��촿Ro��e�N�sx�e���w�O���P+�p�A����������=9���;��8G�<����5�%R�|'�,C�?��d��h�w�j�iHG����}p;u@���g��*����2�t�i�׵g����埻���J~�q�6�O�ϥ~Nj�u��xe5��%,_���o
U�_��ۥ(���brH����A���,��܅���r �m
�+*bcD����Sa��)���ZlB�����+����9bE_�4�n+�.��Mȗ�IЄ-�]��n��5�qo�G� =�|�׎�bR���+ �	���m�w)\�qD��%���X���T;��	N�>퇄G�ލ�u�c������w��������<Y��1S4<���2��ݏ��2�g@�-~K�{����>������ç��m��:Ϣ*�����ڽ]��ٖ����b0���h[+ %��t�8"]#͗dZ$�L*R�`sUZ+�=�Ҟ��� %�W#�	�X�)��4i�.�:��s��ܦ��K�"E�﹦�M~����_4����	\�/o�~Z��Ne�.��l�^N�����`8Fb�m���u�l�*���nem�Ү��iU1�-�2�6/����ح��RJ�䎥�C{?�(�?fs��`�*i��j�Qg5���E<^Qqi݋�>o;�q-�g��vA�m5x瓴���w���uֶ��_��~�Be��^ �H��@����a(������{�����h�@���~8�-%�F�`�S,������>v���e,N�3�&'K���i] (|��A����	y�"����VEK��7o偷�xh֞���N9�9W��� ���S�`��5��iH��F���4�c�㕰$�>�Sm�:����k�j9~�4���q1=��&̾�� Wv�Q���`�g7��H��x�;�m�g-j��k�'�~B�!l����_�x����~.��A��a��9P"4�.��wgD���}�z�N짒��� �2��Hu%d�~^8���͝�߄��ȬAY���������q*�j,#-���c�oƨ�D�^Fr���G��������<����BL=V����?2����@8\��v�a9m���,����9��Ex�4$6RT�@� ��K�l4��Gj�=��Y�.��̭O����s�gQ�7���O�Kp)���I��3ߣ��\���2p�_��Y5�t%쩵�GK�j�I\3�s?ov��<���*���#Mꊳ,�S�ѭ�~�PǨt�䦮��������f��A�ڈ�Ձo��9�+�3�Mx�J�*�'Y��3�7��Z�q�X9Lv3�Y�_�)�\���~"uj^���X�'�S�r}��W8Ve��Åq�k���@XvH�wF��h.@g^}��q��������T�q���|X��y�܂�U�ٺ2l���u�&� 
�Z��'I�x�xX8���i)��s�(�UD�ZVL�+�S����G¼��G����3�<���å�.A�\����C`?++���ҧ/��t�v&����mfnp�:8��P�}H�[�W(f�q"
Y��?��Y=`;n��N(Slʞ��0]9�Mif�y�Z��R��;�"\�wC�I� {ߕ�D[������W�����[8j\�i��:r]�cs7�\�	��F��Nne��OЧ6ץ w��-qR]%LZi>ZR�T�&�ؚ�C��Y��w'��ܬ){�{��#[�i)!��,i.����vQ�P��T�����d�G������0V\-tȃ���A�����
�gŀ���]�mHV�v��X�+�����Q��AS9�p�	�f)�y*&z��1
{31՟�:��~'�Q���wO�4[�f)�<��oBT^A����h����L.N;	�� N�^L�R�5Q �^j /[��5��yZ��@RL�d!��i|�����s�<��u�q��G���!]�u�!xvš�{|��2�n�i����R�d�i�� ����lt�0��u��<Eۖ�`�@<<�3%â�'�'͐{)�RSd���YG�u9������.#s�+8ח���G�W|�9*�1�k���β�jI���ӵ<S5� 7ć���w��B?���)B����4@Y��$�؉!�U�Z·]N�w�DB&#�p����[�CZ�ɻ��`��=!�������sm^��M���#@�'���
TH�9����e^D_1t�J((���CR,�N��j?+�ѵU<b��E$�k�VyaRgRj����m��2����'_А(ܪ}"���Knb)C9q�[Ʀ6��Ġ�