��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn<����d�{�Tn�l�ed�Bn��zX�C�*�g�P���;ҡ�dq5�t"�&-�6=K��ƾ[7���%��0B���$��X�L&~�w`�"b��i\&VC���J�vj�:���]����VVS j��qՓI�A��W�S�l����C�Z�W�.�養c��X�6��%���?|��4c���{���A�'L�����) �5�L��-Ӎ���u�x��|�\;�����[H��\gb�Aq|�md�.m)�0��ѭS"��2;´�8��rε����\q��#SB�M���w��\�7Q���& �]u���O���L���ly3��ͽP�ɀVs��(�n�����B�R2����=� ���V���o1�W~���^8�S^���u {JD��b� P[eG\�!'�Sgqe��5�^�~է�Z��88�wu{�?�.� W���k�z���Õ�;T�}�g�c��9zV�����U�u�%|ť���H�3��l���,+6�b%pyX`\��M�\��ߡ"�k�Ӝ�7W�İvs�/� �p���m��Z��Nl���c�*��y�]�r���3���\2��e%u��Պ��:���`���mꅻ����m�������%��q��.A�j�5��0W���9>Q�M�MH�OX�@�#�j�"��6�1�䁉�be��[��#�B_�f�b�}*����C��P�Hs�Rh ��L�۬F�L�"��U�5�?-4�R��'SQ�5P��)  <��ȫ
ڝ��%����zA�Qt5
[���)�1%�iw��n�!�[���Z�ض�W̎�ґ 0-�Ҟ	���o�\ε�B$[�r܉��q����8�iYDH��A_�<�R�~r��o\�I���C\�π]Z���D��n.�,���$�Y���8�g��� ���Rn랼��=?ng]iUN|�w��$x�
��~$��ip p3���h���eH���3�c��&
���ݭd����ʴ��
;CU��-��`���9�?"�.%F�PT�V�2�&ur��{RP�~�_�M1�:)��л�C5l���o~���]�&+�����|��P��	��*����p��/����z���`:13�ɄJ:���Z�HI_�WۍљQ�	O�Z�\7��xи�tԝ��י)l' �5��/�U�I�0�fڗ<���MmHo���ì���Š7�zU���d'u��>�3`T���%��VM��>b�P���yH܉���%���dŪ@E��|� n*�lC�[��AE�ap���.���q�h���y?�o��E��4a(ٶG$�����>�4�Ԙ�K�7���ti��D���D(� z����n�ڳ�.�l�{~O���^�u��%����"�(#�\�(�]���-n�a����Z�~ܪ���|���WcT8�ʜ��ll�:�J+�c�����BQ��r�C������|I+�݇Y�t�b�ώ�v��eGW ��*`H�E���3Q#/����H�Y_ã6����?�m�fٹ!}��ܻ]��)%��s`�SEo=��6��䕴Z������e���%����1��dm-T~1,ZF]��vz���l=���V�S���e^6D7���.'"W�mS�/*)�u0uSׄ�Q�'H~�v�L"�F­QT��0W��7�m{�M�e`@�L2���@�S+*�'�}ؿ+^���D�����rD�%�ٛ����Nv�S�P�����!���%b�1�x�ݼU�M�������u�}�4���R6Dx���@�x��^�i�\�mG6�$�ڔ"�b��8D��e��;۲Uy�]B��b�������"�� W4D�{��8��Ȅw����&��L�ꖻ�pCf�M�Őa<������܇.�Y�X���3�,�H��l^����J��8��'Tz��K�~-!	�ȱ]�"2��J}9�@lp.$���*�쾟&h�|{�=7�S�G�<2L�ujj#ViX�#T�O�[ؾ�"R�PcTr�R��R>���(�m���7�'�l@`"}WcA��m���yo��JZ�xY�G�p%�2�(�
S�x8=i*��1������3�<�6�����c�����٢:�c��X��<t�� )���7S|��"�nE�κR��'tB~���	�#֘? �7֩�잼M�ܻ&&A�����l~�����8��i�������芃,Vbݗzi�A~����)��ܬ�rr�z��urg:QX����4�.�L�Xw �ާ�b��ױB�������/�����8�8�Id��~�MR�\�%�ihOS�g��E�3�&��pR�g�)���i������ES��L�v�r��q-"�q�|d�]n��?yw)t"2& ����������,~zHǲ��7���G�ٙ�_G��fN�����J7��Y�A���|�$|�,�:b��ӄd+q3�~)�(��{zc�~T����ʡ"z/ѷ=��w���+�c �<��ǔ�<]$�?��Yd��t�Ve
��2�~�Yr�4���G!Y4d�k�I��Z�fr�N�U�#��H��1�q;+q���fD�]o;�w�79;Y"=W��G����μ67���䕸��\R҅n��sR��XV������
�-7�nP�� �hd�$�56�\���S���E�JgU]<�s0 I�ű�נk��f;jb��!�b��&�&e�L�}|	�,6���hI]D2�YS8~�Cz��8Oo9'!��d�b\/䯕�"����D+�u6`nm�kQJg��`r�����xYOŋ�KXy�C����~�K�j�kL{v�B�c٫�*��G�����A0��'�3]�)���B�'��F,���48�Z��-��Š�9tib?����h�;���+)Nt�#�ц� �Iy67.��6B���8ؖ�E!�K"ؚfD�D3`��Y�����OX��!�8��fzb�s��l!8�.��C��t!���tp�����gX��.00�"��Oa���=��'�#�#Lcoo������"�+ T{a�����N�o���Kp��p�%�DP�:��!��F�4�I|�ρӬ������	�������!l��У�W,lY2�1��@Y�����
����?i#�.�J�]*�Fz֝�ٰ���#�*��vM�J_gCە�#x��"�%�ˠ��r�:|A83���C@I0��*����_x�)�%�Ϯo"ܲ
�P�����$>�Ek�߰��Y2P��jea���aL�w]�C�X�a������P@��[F�f���Zi��ܺ6� k�a���]�s3%���|�����zR�չՁ�w�8�6�������� vp�(���TũEm�b��ιc7Eu���^���Ѐ��9�BH��{���������E�>h����.��fT ��guN$9����:��/����p�cd7�Ar9�0�g{)�B��
�L�1�i���IN�n�t��<]rVR=�a�z}Љ�Q�!�}i��F�E���q�Á��P���I�9AB.H�hAR�<H�1�/k=�e�ڋ����LZA�M��Il�������#�;�9�,���7���a�����&���p���YY�P����/�H��D��[8ꇼ��G�\Pt>��ּ�(��P^&�t|I�2(�uO^w���`X<�QCroɾ��� Z>�����k5CӬ��4���N�J�^�(��h��XdOM�ay;i(�F�'"t������
.�@LߴEc��D�Z�^��oA�+��,C��L׃�ɱk6UO@β����@������8K%������|B\�^��o�!�Xܓ�0��iC�1I\�&�H,��x~�L�_���ٰkO:���k�B诐�����8���Ԉ_�����V�y��t��i���w~If(x���8C�|���:�{�M"��w�S��2q9�/I��9�s=��v�>�ql0��w���6��;hR ;nC��6I��Zh.���I4\ʴ����`��������Hf(v[�s��3���nj�>���W[oښ��M�s<��RB�SD2��PC�T��Om���VFG�Ѳh�2�цKi�@����Ե3�C��Z����]�Ji7��]ڪ9����1�nu��oݤ�`y!��~�7�x����-��1F]��*!+��f��$j�c�����t�OX5\��J%���+Q�x�7��A���k���\���;�l���J;���c�oჴ� 뵅��c�����3f&�������t��2����D����{�b�����	��a�5+¢����]��|Օ�=�^ƣuf�3Y�O8�J.���d�38Te�j3�ky�T��Uz��)]6�����-&p�}^�վ~X}nu� -�]�2QA@j �Q�Ɉ��Hk˕&�0�-��Y�y�`U��ǲ�������j�s6;d4�8�/� f�ɕg���)4Q�W!mP��vh[�V9SF|�U�p�N�h���Jݬn���/���-������gN�a��A���S`�+�)O,�OV��/oQM<R祹\F	#���[��쏘�mB����4��e���.��/y�~´���k��W�+��"{������6� [T���K�~���WS�c�ݍ�d�|HRb�ي<Ie���+Q]�щ�;z�&��y����>H���I��~[ba-(�w X�q-�/"�~�'���1����%Z�| (�DL;�;w�֝���q'��e�q<�k�`��~��X*��#g�-��(��E�%��u��Z;�R�l#ۨ����.�U D��Ӿ������}��}FN� ׺~���s�B�q�L�0\��vnl�bx��fW5��?����T6��`�$&�y�E浟^Grd o��u��i�َ5����Es�U�9?}Q��
��P��m��������M���0��<F[EN �ԇ=+�z��C�Lk[�|FooxWav���Z��C��(I\��6��A� ��>���y�pA\@�s�����m��J�gN�����)�6�T��Z�(/�^�]�xd��y�O��"��\->J���G�L��}�+9��A|��fyU�7��Z�Pa9��	m�Q��c(�T�͈�`�Z�ɠ>��g�xÐˇC��`���Ԯk �;$�p�7_r�d"X�,�9/-6���)͍�3�b�ad�SC�1`c��"���ó��߿�Fm.�m����)炮��ub�2���T�V�k��c5P/�\��ٶ�$e�����!�@Q,��o����cv����H��#�D���he#����x��&�p��D}*\�>3O�����%#Œ
������aD)�n�����_���JV�PXR�r!�pbg%�?E����T��|(�D@Y�lf��j�����lMi�1�����c���u��k��J<Zf�x����R�0���z��^T���o`U��*oQ�=8���ؼ����Z������P�1F8�K�_��2�Y^Pe�ݢ���T�GX0����C�}w�����=�h;�D8��㶉��
�^am��u������d`ΐ39�߅���i�"��m/��_�K���H��� P�)M�% ��/�	����H�N_��0�x��fpw�*Z9ھm��!�s��O���0.���R��	�#Zs���U�Q�,c2������J���?�-�D��)�sV�S����N01rߕŨw�_9�c)���Ct= ��>SAݰ�^�Ƌ��*�������j��{�����ⓄҶp��C��k����[�:����(�Cz��	�!A�̘��0�,�ٹ�"�A@��6����	4
��=�e�}R�I%μ@��ː�N�;��g���޽���]27`��h������P��)��7�������鯐�?zٿ=;�mt'�V�Ůͫ�W�ы|{1fFes�3�o1���b]'}�up�!!b�����-*���$��I�"-^;������B��'�+wc�vPzu><c��s�)��w=ˑƥ���v����m&�f�dD�o�۹fʢ�0λ˨��M<O�����әB6�J�]/w�Iy`@��:3��ؕ��v��( 7\�>Q�>�f���J��с���.R��;��"/)J;qېk�=GXoڳ�=�0�Ǐ�_R�\a�j�r�o,�DP)�`�7��-Ă����j��X�d�@����i6�ɟ��#JL=�$�9��O��-��R��ޮ�>�)��������tu}��"�7.ی}��@,L6ʦe���fT�XEU��'#@^�W�	�+xj��z��r������c��-�?�u���N5���L(��x�}�e�XZ�l�� n�x��	��_��kw�J��}�G��K�ՙ�3������
�j���#\W�Oʐ�I����6�i+�#�Jbk�u��U($��H�9�]�T����|&"��>z8�Z����%m���ɜ%}���xq�FjҾ���ብ]����h�8�ǆiɩ �Gt=����o@����Â�;�2��~�}-��N��&��r4�̤X�=${W��ף�&�"�A��J�سſ���BX�q�1�w����]�t�m�<+�������(������2�I�� 92�ě��رOh����Y�m��$P��`oaV�\u<�L���b��6V����/�I�L���S��Y)�&��{ڌ?8��sP��4��D�F��S��܀�<^���mk�0��W�����c��	V�-%L>bj�� $r[�e���������)Li���Y�Yca�b5��@*c\8u=vl�O���T���V{�F@��{�Naj;��ZV��1L.FQ �-���Q]�.l!beFjjmE��E#8���x��UV�;_̄�|�.Ӟ��2��@����eK��+�4�F=��ז�x��T��H�
ӒaF�F$%Nn+��)�I��O��`mL+`��4#�@U�pQ�|�I�M�Ȝ�Eɤ�쌆m
y� Ȑ7eh��bP 
n�P�����b�=�1G�D~����݀d�F�9#�����@��}���_g��w_A2�H`��Z��ٱ�|;E�n;�����1���m�N���kE�#&�Im����"�h@���}{r�W��(�.Tr�4$� ��&7�՛�	����Ю���5��b���5��Wji�����~�y5�>!�f��a�1�i�uo |O0����7z$�Kyi�W_;s~��$G��%��l�j�d6�����$��B�Q��[����$�QE�F��l2��F&+�E
L��=��!����;�2B|Y��Kc/��Þv��w�tQ�2�c��t�����k�+��~���}��!�q3j����ji@�<ʽ�	����Y�	o��Ns��d��ల���=��E!���-t�J��F`M6uqEB�C�bM�F6Eզ��g/i��b�q��#�{�-Z����zL�e!�t�jl�� BE�i&i
����g�uT���L$]j>�u`�����$�d=�C��$X�H2����a�IkG9�g�J�[;��u9�� �'�T&M�Yx%�I?��B/Z^f�E&/����0XQ{mmڸNv�8��0�}�=ߠ٩�=W+�]�
�1K���2�Ǔ�y�I���hJ�L��۫#���[}�P��`����"�6�m�bxO�2�yo�,�N�p�֞�`���	z���j�$=�\PԈ�'kYY�_m)�?x�$�M�nӶoc��bF�1�`!o�*#�&�~�Mm�<c��@�VUj�ᎎ�O(9rP`<��Ck
D#&n��~�dT�~ۯœ���+�[`����/1�m;�'9�9/$�ڹ���X��S��i�GVK	�Ɩ��q�oܪ�������ӝ�A��z%2�����U㋝�cǃ�>.r�(ȭ��
�{��]Ų:l~!F�_? �jC{3c��^�A�����M�(�<Ӥ��Fh�n��q��xF�_X<�nr@ע��l�O���^�ߙ0A����D�h��*��\dC�"q;�xZˌ��b"U�tp�uF|��[�[o�sJ�l�J���qё$�늈��c���/��s}�`Ϥ�V�pZT`�ǃ̙��*CE0��$c;��#���U� ��~����6�"��vVz�ڶl�vȦt�g�x�/��us�v�����j�;ը�9�NRl�}�R������!0�/�I���޿�ꔏ�����A@b�J>d�0�p��x���S�挣���ƥ�L�z���ށs;×�o
�,Z�hC:6I��G��!��i"Ĭ�<,:�g"�A�ic�X��,iJx���>�s0/\�[�ӑ�t�A�}|�Q%M�,jn\�Xj���k{�4���;�lO�XY~p�. Ec�apqo=nj��'�S�K�����bNk-ê=/��7ig���8^�z��oz1�,���K0�ǩqs6_ї|Y��~��(�]b_�J��I%H�U	Vד����Ex��4Z[�̓�����7��,C\�hG)�(�YӐ*IF5;�kyo���Ã�z��%UAʟs�&��Ӂ�	�H2�$s)���ۯ��s7A8�W��3�*r�n��ؼx���>��"��#Z�m��PJ5b�Mw��� ����rUC�IX����+IUi��!�Q����q�SR�!�����QH�kA�n(B��8h�hDLr�'���E�w,�ح9|�c�ć����P�\����\�4���?�pe,0n�|�{�a�n1$����Z�e�<��K� � ��Y~�]�XCU��Ys�Q6��Ew�TeI2,9AXl�����S�K�v'�q�V�-U�\�f�q����;�t߾R5�>�{g� ���P"�aF8.�ҥ���_�0�3��'Q�[E0(��ft����:(҃F����he�L���䍂Ŏ�ţP?��"L0����&����ʎ�� L���䊷mu=8xL���#8�u�G��[~[K璬�1�o.�Ǵ�y�ܸ]� �0��d��� ��ncԸi��.�ߵ��0��<r��w�'�����HA�A�s5Y(%���	�g��V�PJ��	F		��e�@�KHN�{�&� 1�CPU����-�0���+��gE�٤��$�J��2��/��{��dЃ�s�y�L(ට��c�����[&�I�9�#�l[����"��$�e��D_���sSj��d���K(+x���cʾ�?��&�D	b��{ˇ�a)�ͦ�k�O��^'� ?+��ڮԙ5��2�5n8���*-�~�y��J�v��R+�rw�"$��K�?�p�l��� �F%��AQ}����>����'bK�&6s��[�E�QP5Ǡ2�Y�����y�0cyu��- R쁭e��n���e���c��O�7��=M�,�6cg�a���}s�.�������2��%̣5i�{�ر ��kx���d{�V��?�p���]����t6�n�݆�6�j�������tC��r�\�'�S�(Q� ��_�^�8a���uKLԂ�S>��'�jCJ��r��Ǆ���<���v����	�^��#�#Wbl���Y%1��vk��<��9�Gq�(
��vu��a� CWASs~��������NiݾR���i̜�س�|�VƜ���6�Z��
~/.� vV�}���b�T��
�Z�a�Y��h��4�2�`zcEH���\3@�gw=I��o_>/Lx�a���l��\�4� e�i;긻c��\-BQHa�ٞ{�����%��ŀ���0���}�c��Jz�禋jI�oDK}���섺����<��f�97&lϱ���g֢�
׹���d��l��#����+K��~�"� ��S\Pm0�rc�p�'(l�Za�2�ݥ�F���$��@�~��1#u�RBy�@;�a�Y@�o�{�,���(���X��=�Tڡy���7��Aw$pU"�V:Ĕ�W�[�܃U�!z�bJ��!oUB����������	�.�SA��d��F���,�T�p�s�f��3�%�a����C\MD�0k/)��ܧb�ϩg��<l�V
�H���� CKg/�D�?�5n�V}���C9���;��2;A�����s�Y@�/(��Q��{D'Z�UO�2�G�s�N�4��Yإl�Z�؜G\��gmKZ��K]Kn����P�Z%�e�	^��G���%���-c�n��ATɪ�K��(?d��MIw/ ~��D�+����{��y8t��U�=P���h����z��R���X!U>�o�_�Qb���M�sP��$���\��љ��Sʈek�Z�<�}��h��퓖 �k��nS�@�����a�}�����6[f�/7	�� ����a�S4� �4e��1�*m;��!'=������A٣u�^���2j2��5?$��dx���Eħ]����K���L��
qS��
�[,O�)(c��F"EM$���خݸ!�b[�݋^���՗Q�Fv�E`��&�X���~\���@J��qe��2��ˌ�� V��XG�:&�_�M|(�!���<��G��LV �US%IY_iI��XѴ�O���)9��<./v�>�&P�ҝ<��^���pI�SQ;4X{�D
4�'8�7pT���&��>�]��TkSq�`/�[1C+����@�-�����R������Q�&�:�&]����Z��ֲ�C_�ݬL24@�JV�&N�L=�˵��Vr�3�+���D�1IZ�_&�i�w��"ag.��]v�����%
w�d����7;�J4I�F�J��,��ʫ�l�H�0 ����I!څB-�"���ŵ�z(k.���XI�W��a 6n��뙡�>���0�-�W�@b���,1 pS&퇂��Է�7�N��Bb�L��Bbg)��j�I ���6�]�I-����}bhN&[�/����R�Hm��dg���h��S�!M9�A��᥵˯�7��D�l��� Zr��\ۙ^�y7mD���XL�*өx������#G�y�f����<3��&=��g"�dP־�)�V���㳼�YlO>e0]�lRj�雦�۰��w0���&�(�s�k�������wM���ٸ�Q��� Z0��nZwA��ud����	ӝS��X �I@�/V�%��L��Q~����4��ړ.&\�ո����&&ch;�W���m�
�/4ئ�N4���$.�ҤV+3{��g���z�d��ᑖ������fw�!p�	�'|�h6X�ˑծ%���f��1�&d;8����q�Ui��͙�f����է�%M��<�Ne�j�1(J��{�=N ;1�C��oCi˩N�IBi�c��~��z��a�;�T>Q�����Slǒޟ�,�w�\N�!�o�#��| ��lh��)��3<�	#;�@�ai��]y'8�/=A#q�b�K�)�U5X�u�yw����Lhm37gMZƊÔ�U���+� X���ȋ����d �K׈=>��ZeHs��������]������-�캍Q6��ȁ��P4~����`�u �\���G�=_�m_��}��#b ���1v4I���k&��Nx5�^ټ2�,��|�=��R�(+��a� ��ʼh�7�e�M�{.gM�r�9��jV�[�+=��	D�B�$�^Vt����X�4{�	�2u� 	v_�jN�hƭ�9������Z�$���^��+i����_�^�K��0������o���<�lf|;�ٿ���G-L�����1�y����9�����O��["l�Dpw�	Q��j!�z7��܂�� t
L<jՐ�&Χ{�	R�\M�
�P�s_U�������2�ڹq���x�qh#�6��1��M�����3ˑs
�xv�N�>�
r�3�/�>}��ӧ�S5��<���r��@{�p����|$A���V��@��B�w_�� h �D�y�jU4�A@ G�Q6��Ɯb���AK(rWҁ��5m2�f_�C��"�"���=�4�$M�J�W�����d�e�s�G:�%k��U�V7-�J�6���=��S�B�� ]�\����q�/����;7�,�s?�4����7g��(XB�vf|y����%�ac���jW���\q9����QHvtv�{��':M�KN�&�6�]dm�h_|�>s~��e�ݕ2(�s���7$���A1��$��4����g!3��)�˃�<��t�(�5f�<a�4�(��4�p]�*<��/6�z�t�����]l����m���%�􏫉n�$쯦���&C���q�dy���ޟ�n��(���p2�|8���dI�B��׊�G� ��`�r�e��_\}��@�?��R|�����Ɔ���p�m��A�@���C!��h����RC��;j�6z�F@Xe��Y�ѲS�v��]p�5~�c�.7����$'��I��B^ h:B_��k���O������j�����F1@j��R#P��%��Y���MW�	�&��il�Д3��(�����408@W�?�0�t�MQ&���(sw%������	3kT�Á'�Q�E�r��o.�� �xL��*:U!�5��l��)д;wK`�r0�*9��+Z��d��̂�&/����rH�v�v3��|��M���EsйB����%Ղ��݋�80��8�~�4�:��<{�~��k�x���A�{Co>� g��vv*Ff�j:y~,����ɳ���0trXCxE�7<�j��b��x�E�vxdu`�A�(���ϼ��J�*,D�p3Ԍ	UI���k��/rN"CC�e")�
"C�F��a�~��#|�T��`���	����q�ۻ�7���co�u��U�ԙ�_��ڳ=�����io�V�.�����k�$I�^\�Ӈ�&
�~x���g����G̸�Dl��������ڐI��Ҵ�ɰ�t}^�@�7�
B�W�����1�z��n���G���q��8VZ I9�]7��Ų)��b.�-(�j_��xM1����R�},�>&��1Xl��݆��y� ;����"��|�{-x�������Izo{,�8��Ԡ����6��iJ�i���DA�"��}��Yu�[u+a��h��cY�t�aJ23�4�4�4����n����;��
�qgΡ�ab������XO���W�����I�ZA�>�(Z��v��<��{3��8�X�����^n;x�3��n��>HÆ���#��G�nX_��Qv$��	�s3l���>5��#q�+ď�-�QJߧ��Ț�?�P����@6���h���=���c����׷��ov�@ID);�u�@L��Q8H��1�I�o���ِ�\y'�`� ��a�B���<��n�׎F�l횆�Xщ�n�n�q��T���g3s�=�ì��iX{뛬�"���@����ٸ��D�<�u�e�Z+�1��ۊY-J�G���q��bj�8cN̑`g�cdblh�Re^�d�'ux�5$?Ꚙ^P�u(�W�s�ks�o�o���L��D�硫'5���Н�k�`�"�G��<ɟ�A���
u��.�cQȮw=�֕)!�r��+l�ަx�d���3j3���{)���e��9����ؓ87�lWo���vY�7����[���_̖>�#ٷv�1��0Ҡ0��yr��.��d;FLMx��D��<�oy�]��ؔ|�L9{����	8�����&��8*�)i�}^��w!<i�v�CGQ�9���
]�Ri,��K�S�&����T�0;8�~(4N�m�s��I$�0�vA���T�� ��B�N�18631�q��Ft�뇓w���������"VB�c�.F�5��(v2����G�zp 9#�`�������V�v0�ە'e.>`�d(qHaэ����@i��a�d�moZv8��$otn3zD+�9��O�@|��`�X��x�k	���Gl�{W9P�u7b��)xIp�XT�XzN��׺���
k��i�8���a�4M.��u��#��o��J5���  G��	h�W��E*b�v�`g�Կ�mp��~�z��S����m{�QalR��,�a-������^�1���*C��"�˨���%�����4�k�_�h+�wN�:��ͤ3J�ƀ �Ⱦ���m=ם��L�"�`���B7E��HC�%�Q@��]<&�/���-Q(��ft��>�եq��v
��N�g�u�����kϡ6�&��-�ֶ�J�P�^r�t]E#���*�Q�C-䓅�������d�x�;�c�!>�gvիF��c�j����x3�*�,�r��RCk^0�#��'�KC��V�y�\Ud��.��J%��$��3Z�E&j�HYtع4uu��o���7�J�i�3Q�{B�6�wL���l�\^�A�?��r�n�&��$%6��˱w-~�f������l j"���I����uIJ�~H����{RZV�<[�t�洧`8ԴQ��[��6�!;�K����{ !���Z�08N�!��%[�e:�c�*<I�H<(�|D��D�!�@w �J�s�ך��Kz�OOT �����P�bn�6����z�T
"����Љ�4b����R�c5��I@ahMӅ�,:��(v��[[��V�m0��f�Ղ�.�����lG2[>���+O^�bg���hg�-d��]mV]\�3�����Q�DL��ư`�6��CyJ��M�NPI�&�&���DE�Ý�ϔ�����f�vj/J#6��IP#�_�U��|ѹ?�������4��:#{�&�{0N/6��ߋ!Wr G�h���Z��j�fa�9)�{<<�@�K��K�'q����3�e0�w9���@軉��ыRz����k8:8�<�^��ϟ���`m�~��J�]l2���Z���@��2�o|@���b3Rn�C��k$5=�ˤc����O#��|o���[�@�j��0{\����-N�M�z!��B�|乳�:�m���?5\θ4� ���d�[�����A�� �l�z�2�9G��u.���rb�����h������v�����P���ACr��X���I�463&� �0��������u�%����G;�&@�[)��|���\kYZ���K\'W�N���x2e�CD��e�f��_?�%�Dt��Q�gM@� ���A�e5Pj����R����ul��ԓ��yO����ǧ�'j1Щ��?�N���1V�}�1N~=%(k�9��͏�������IB�'�^�W/n%�{(U:[Y�O~�k&��;�+��=�g-�����b�'�p��?�!�Ih�d�7��_ ���w�gv�K�{�6��{���J�z���g�TJ�*�B�$�G
���Y,A���~%�Q�>iy'w^m�׺�OUp9n]'������N�� !M7���K��+�J+�x���4��(3�Y��u��$�Z1�F}�e�^�5aO�Ƽ�_nD�T敂t;�Y��{����t�v�@�<��j�S������O%�������S�;�kTJ)�VNݼV�[`u�6�V���K��*�k�ށcв�(�O�!E1d�f���h���ya��Y_��ư��݌�Gђ��s��.6��m
|/����jd	�d�B���R] ���X7md�"-À(�lyK�/�N"q���6�E���|�}���J^|����8�x�ϭ`�c.f���W��p���v"<Ò�ϣd06ĵ�i$4 KSd�uD*qє��V��m����?��D���3����<�C�t�<�Ӄ����x�n˙k��=6���J�*`�r�:�^Ǐ��!�ю<�J9x�����/|*��ұ����;��l��L�_u;iE`�܃���&�5D�¼ɵ	����0�
?{�M |�a���_kz	�uƣH~���Dϻ0�<�$�ŒF�-�|(<����<nHꈜ_�ҩ���B��0��D��֦�X���7 �\Q�tg�>�TO�w�wʙ�/��GYg;�7���!;7��>���0�����dXa��fxk �N�A�?�?Sc�ӊ|%��)m���V�������Ƽ�B?�����"��SeԼ�'�����O���o劸=�����9��=�3�ԇ_Bo�x#8>�q(�8|<io���ܖ&#zẌ́!*�s�D���	@WRs��C�,� �[�ۙO�0i��\�ܰ�l阗N.�:p� y(�HD����;T�9az��loF0`��{�ʳ5��W1��`��`�g��I)���.��V	`l��S�� ��z�s���挀!2�b1�%D���c�U<9����������1:Iu�R�:<8HTs�k�05P֚)/�xMRc�d���-.W1���҄����N-�+����x?�ɦ616I�J̵Eb�!y�����(�^���[w��45F����C3`�"�Ӗ_O\X�q�Zw%)�hb$P�GƁ�21�ɯW��-��z��<7�'���}/�;{��H_���F�S�n���w[7[3V&��pϐF|���f����-�c�PE�e�-攝5^k�]��V���z)6kC=�8#��	-�;Vq7��dh1D����ڸ��"ٻg�'��L�M�h4P�p���[xo~Dm��>���7.%`��
��3m�23}?�LӇ-$Ǣc���\���E�s�v�7���<00�|�GNX��R��)w��H�$ خ%([<U��?g9����جg��n7iL����x���� Gz�4lq9�]������� ;G���p�Uliz�� �� �2�����WZ�m������(�Ӥk?��e�P;�5����d`p�,���&�7�Xw>1�Ǩ�M�5w�Cp:�͋��LN����}�^���z���I+�Q}\#Jc��5�E�"O�R����o�@d���� Iϴ�yn/<�V7�E�n��K�i�16A�)��`W��a�'�0E��wD���4�{������-tv�qYK|��|��}n�����<@蠩f%�G+r_i���et�`�7&Щ�=Sb��A�~C^�mҕXJ@�k@�m7Ƒ��J7��K�6Sb���A���An��r�Cn� x0��6}i�193IZ�����8����ޮq/�K�<��; J�zN�c�'��/��a�*׾���d��V8��Z���)��ל�0�ǘ$h��ć�?�:�GD &~O�]s=��e�����=CG�N���)Dٮ����ƃ�WR��Lp��1S4��IT<*��.L���������劄�/.�`c�ק��`-󬭗��V����p	oů=._��^_�
P��=�]�.6C����V2<[}�g74,Kx�TwYOf�,Z.a�3��9}�]|���؆���l�M 2�9����M���k�c%����&��I`դ*�����D. �R>��*�.1SǧЛ����D�˙V��Ba���M��,EL���8��b����n��E1Ȏ�a���$$���m�)A��}�!h�U���b@v?�r�l��r����*��l��Ľ��u�H.04���RU��0�+.�#�"B��gc���AWpdI��dTY�p������?I�61O��mz�N���gE� ��P�vi^��dc�(i��]�<��Y�p�ı�'��f?�#�\k]:�A�v���
_��di�ߤk\IN��mN��,���5�{���+F$��~��(`E��"�����xb$�O�Z�0_�],����|k���մ���!G������qX�BG<�S"�J�&x5���]mh�9�n����>0�y/y@�X�c���g���h{Tx1w�T�:���M��,
�Ŀ���s�yg0�v�����5�D���Ģ���z�f��4��t�]/�g=��K�C�$N-�L��]Mxap_���+b�^�y�!6��p#��͠��<���[̣��3�Bi�\9��(`�-�1�II�K���G�fD��L�^M4���}����=˨�L�y�Ө�s�ַ-N
U瘃���pw�mKHP���<V\�2�	��L6��7�=�A�H3z_�3�Z�R��C���Uc��� t�V�Xq� x}&Q�-X�Z�^nخA[��nr2�d���/2sC1a*�/^k`�)6M������W�5Y|8I����Yeq�#�Pds�Ӣ~z�ȓ*�
S	5JF��2�ڦ�,�� sC��b�Z
�ދ����(�����v��29FX��y��T0��b=��X}5� ��_[B?|%�v�h�c.�U���f������N��+��Sm^�#��upܐa^���2��ahN�I���"4�s��U@���Z�L�0��V�;6���������7��{�����ߕ�v~,�=��.0��zbu�iF t�D�یEz>-��g�^�����/H��p]D�b�FY��ܾ����i�'��i�^�4�a���vOs'h��E�N���I����Ah�Z��:�0�e3�g=��w`�*)����&�X͎�ء�[K�|{���q���_/{� ��nì���9���aY ��0հ�e����M9.���y�݀�+��m�5��]��h��K
r'bJ����/���@P��$�������@�ƞ�&�\ ǋ�H�^��7c�]�2&ܩ��e���(�Y�Ohõ�Ǖlh�?�\Qg��n+^w��ȫ�h�=�5�|g�kE[����~$�x�@jnɊ��m������2Ĩ�_�,�[��E��tL8���?��SPR��`�f\�Gc�A5h���r��������y�q�L�2 �^�1I��NB{(���5��ę:E1���k��;�%a���vאKm�N��xz���ϊ"�?������@u{�v�ٷ�@)/I��)�;�d����'b��Z��Ϭ�n����[�@� ��Z]V/�ʫ�6�Vo[S@n��*��#Dd���H���4�$�*0��A����:��*1�F%Y�m�5�I�#D5�P�1�����d���e�)��/��-(���۲��?��8�&i`F����ͪ���\�4���`��o�:��X��J�x�o��::)3���	mGYq�r�e}���T�$��[c�X��s6�_�#��