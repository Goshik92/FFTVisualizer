��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@���$U[H_#�/8�y��,��F��`G�m6f�f�aiI`������tC����dl���=eZ��^�٭����B�FYĸX�G�����݁�]}~�s�cC�_�V?o6���p!��#��9~̢z�x	����M�8�DӅ>q 6��n��  �	���Oi����P�ª�ج�9���Q3��eS�&�ʟ۹����:�V�ۂZ/'m}�Dv�Cf��)B
�n�ݘ�I`���e,����i�����r���+=���%{��V�ݴ����{��L�����3,{���<�@�3��N�0X )b�t��~����=����y��(�l\�m\���?��B�*"Rߎ�R�ʃ��t�6
dw=y`j�2�e��J������^��ò��-ƀ˘��yqXy��1Ȓ��h*�׈��.�T	森�y% \PU�*AH��i����Q��w�YH�#�k:����db�s叢]����8�Q�
���d]�5�h�Vr�(��C�c���¸޽`f���Y���#�:D?��.Ĥ_��5c����D�Q�{\l�M3�r�������
n��b�������6AZ3���r���%���Ly����7?i4p@�tƛW "�o`α����n0��dv�qnh9!��П4��[� k:{��ERS4�ۇ1"5�E:ԄxDL��AFqDu ��b��e���6ϛn�?;$�=_�t�s�RL8��""#�Z=vv|�g�t�嗻CYY���m�n���
����|�E}������aS0"d��*�q��h��a�9��Xy��1uY-6��Af�����F_���Ԩ��|�Ч���_�y��\ g��H(����|�&�D��F���Vv��&Y�kP;T�7چ>�tH�w[���W|��5u�S�p��[
�>���B ��{�t� и~h�j,^@0��Ƙ���(6�ɉw�ި�Q�D�je������g�����M��i |�pȈnЏ4<�Ը/�%�{��ٯ[���>�;[�R.����&�+z4q}�l��M��F�U��&������g6MN��ȕ8��Jm��s0:q��`d�]̽Bi��Kj�[5>0��VU���Ii|M.T ��V��(���sl����V4�$L{֥��%U�����ynl��!� ����<T	���&��.��{�9�����\��?$��xf��h)�~��[�7A����}$`��(Ņ���m�$r6K!�S���YD�e^��v�J8S-}�q0M|�|���E2K
� �QPȓ����*�І��.cʙ��s
�rp���6dj���x��'�m�x�����������=30�3[ W� ��q���-ĳ�����g;�e�i2�I�a�ļ��`[��GpPhY����yM9{��7��־=-���m<�Ձ�u6�S2g�wF��#�5;\�8*g﻽�d[����-�Fn
M�<�gRЁ����q����1��m���T�ǂ�|CL��W��-�Qá�Q�s"k:ה��:��°�Xq#Iޞ �����w��f؆?��~�b�h���"�jȡl�߿�~�����Ts��s�&��?���P�y�6渚4�׸����6�l+�U�".�f}�V�c�@�C�!������4,��^sv���p��~�I��z*�1�T?�WS�&B��/�$��FRG���JBH����呐T	�
�Z�>1�b�$Omba��]���>�QR�:����S�� �@�V��q����jڇ�f������v��x�C+^2ږ���9 q<���
)pvT�=b��=�$dB�,���3c�|�"N�\\�}��M(��y���V  ����Ŵ����٧���sy�q���ӷ�r(Iy�F��=����R{��|����iv��͇�pdJ�X2�L=����2B���&"�kh�7�(I㫁�zƚD{�R�SA��X$؋eF���*jw�%�UR*�L�Wf��jOE��9#DI3{���%g�Pa9�dU+D�qHͭ�E�� �'�쎫�������� ��yЧr��/����_Gߦ����1�	_���մ�{ʿ �/?��#�?-s��#�Ŏ�9�Uq�_P��mJ^A��di���)�e�XF��h)s��rx�I�f�#8��k[3����,[�u�3�:#���n.G��g}��⟺��!˱O�66�XF��-rÀ�F�e���i��r"E�b:��y���Ƹg~����5e��>�]��2	Z@�_~Z��q��7�cc��(��AeEɱ��{Ð+��.����H����fO���狊k�f`6Dp�<<�i'�\�iY��XkxO�L�������"JEX,�0M��ό��7`�.R�u�̯�I��b�<�1���{�0�=��f{%�z�}��R�w�X�����	X�VJu����e��O�#�(c�=rW�Q�|{	�ګ5��j�Sl���2���i3�a4K8�<��4wh6��wa��7�ԡ�6�ͨo�O: ��e��V�<�Ae��*ҟ�si�����|eCD2�m�k���>@1�<���A@'�LuMCf��$i�������#�]��K�4Mm�w^Pmwmi'�U�%O�H�����d��#QH��8z��!�]/Vx݁x.r��nc�B$T�kWhXxC�Lr�����s�_��T.<!ݓjX,��1`����� K�4��9Y~�+�S,���̜��;]�bEG�ѱ Z�8�$�m8K�k'z�w<l��y�����(�k�+�p�͐�+l}�2[�]����A��P
��c�F�E�1~��2[N��ꄴ�Q�^ ]>&x�[
Z���;�e���>9߰B!�TzX��םl�$��J?�v%QK2.F5�x͊�%(�}b3��X�r���_R��*_�a����-2SXr�?0�n_3{�:��r0I�B$���Z�}�`W���T�Զ���Ղ�e.���y˧�:����M�)�V"�E�K�g�u���J�/J�v�j�+#g|ԓ0���%Xh\�V�wܟ��&�=�k��L��7~���!���u^�r"��ַ��n������0wj�A�t� �]�Ũ�u4����Д(�Pf�<�v��:�c�&H�c_]�1�Y<�+����C��T[���w��]hr-�Q�9_(��1�Wk�G��\A��zx�9�F�fȶ� �o)��=��c�\g�\]�A"mi��D��\�w��PAn�%ъ��cwJ����Q�30hR:����܄��ϗ�^�U����#����q�V�͝e�z���e�j�u�[3���S<���qĒ��KT����#ՠѐw��l��"�I��d	���>`��FU;����H��z�A��o1W{�.ZI��u���o>���u�u�R�U���0���ém2�'5r�E1��8�t���F��>��Q@���
�~�$ u�v�F[��Ҋ�5=�L����pk�?M�@}����x�O����{�NaA��2�]����)�dw��$eqj�N%�$F����z����x����v+�Q~�ޡ�}�3e�ŝ�}�j��Y:m��ɏ��?h�ʮ(#m��aAĄ��vKLʾ��!���>�s� �}�>��W�GjD�W3~�q9-�%j&�v�вO�0m� ��W��o���*�n��%�jr���B�@zY3��Ϥ*c7s�Cm��b��br���|�SV�����_��&���c��[H�h�챸�^�g­h��c�� ڦ\��P�9o$
Cpٯ-�w�}dD�N�*d����@I�"��VG:���~�G�U��;��wуk�Hz�A�-�_�uW5\^L3�"j��mi��}��^����Cm~UqN��͆��P����֕7k��R^�!!�
s���ut?+��C�gv�	��$YA�J6�,�;'��<�:(E�l/����JȜ��\�>?k�=�dhJČ