��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����)n �n�NP/x,�Fu��D,�C�)��j�vR�������|�]K�U;���A@A�qY@@բ���e�̍�gF<E�0�z� n��Yaex�1��p�+ [�B��;$ţ!
�_�c�>�Ή4�k-�e�M�}Y.tצ"[^`㻬Kg(5�f��#��D-s�q:�0eP�%����+���ݐ��j\�8��n�p������xo��|�v ��o���o�4,٫'.Kq��$�q��\�6R
4�q0����R�R� :P~�آ@�����Sx,[��0�$���E7ٷP�g����w��Ϗ?\x��%�2Ç�n�Z������eʔ�/�w(¦.o��z�2y�m��#��S�F:�..!U1��#U"�SF��A~S#��?;�
�~&�Ҝ*��N*D��bg�K�JsL�ql���dD���p�1�79F�ryσ��zp�+���W(`$� ���Mk�S�<6����%ү!LxGp�̓\�J7M��d��$ �)�.$JxK��\)�ZU�<!�R������#_�r-q�HJrEѢ�*�C:�&�D~�/���F�������^����S�C[;�Z�5����RŤ�Q�a��ߺ�b����+t��h�]�*Ԑ�;��C#��]�r����2���?]�g��Ϛh�D�;�<��l��W��4hJ>NeH.ř�!?=x,����p��dAdp��}�X�=���y �w�S����0C3U����&;5E�� �����>�ݢo��Vr�����m�4��q�=��Ҧ+$�HIgKp�PB�F}6��GXz���x��b��)~#�_�U#�=4����q�ȣ�&P@ ^\����(L��V�:�������e��`�R�Q*���=W1&�ݳ��C��b�k�,F3��2	]�]^�-��ʯ;fg��GG�7f�.��~i��������Fچ����I$�Y�@�Ӈs�d7h�)~.���0���t�h�:�����8m�Z�"��Oޏ_8��n�B"kk�|�TƢWv�S3y?��ߨ㳦D���2e|
���Z��"ĭt҄�X�����Z�W�Z^~wx]b�[�+i-ja�T/�"(���Ѕ�K<e㹌��N9���Q���G���e<�ˉbbN�ۀp@��1���F�ec���@�֨p���\r����_n��� �-�[���4�6`�%�cU�ܥ��E��HR�E$��B4�!4���@�%T�Xh����E��<RT?��x�nsg���`#hn]{��'�ж�b!�jW��ż̎���=͉�<i=g;�6��Cb��_�C�H�7�{>a����Կ������W�f��V����Ò�P'���K�A���Kb����7�>�
=���4�#�X�8NCs[��(XE�0˲u�C�U?1=d��D�5��*^A�Lt�;��D�.6{����h�!D�ٝZ�����S:��lj .&d��/�8��S��f�j��Թ���!��h�P��wL��c_3��j�c��2�a���o����8�J�����y�U�b��k�cxt+�11b�+hj64��1A����K\�2�N_�}c�5����=\-����ԾD�<�/�k���>�=�o� �*wnY"f<�UYFGO���"�%�f�ȥ�������z���uO��C�h]z21��隚4�5�<�G��"�ڇȭ����Tr������٥b��͠�T6kY%�Q��D�0C�F�01CFQZsbO7���C[4���s��f8����`��������'Ă�®�5�2.*&]��ot��#ݴ`Ǳ��\����1_i��n1�k�A���-HG�0Q���>b��"�wz�]�h�mڒ�G�C���,��ʠ�m	��T��W�o�	�1�(���a�nJ�� L ��>*_�j����_@xX5�e��������&�00���Ԝ���<x�pE^)j��K�t���^Ӿ���*�g +vR�>��~k\"f����/���}�Ƣ��L�[Ӡ�5,�;�:��g�=N*��+��Ei#�5���e����U�ru��wO<D���j��*������^v�2q�9/���d�?vR1��ӢVW��r_��;��M�hR�O��c�W-f��"�~/2�rQ�v&�Q�?g�V�T[�:�(te�.^7}aFň����9߄wP^krk��@�d��L�1޳M������\�p}�.�)��7� ��w~������I�5�L��7�05��'���Z%z��D�y��Ԏ{V<���tX�۠�O�� BeP��Rq��U���Ҷ1��xW�	+�z*q8�a�#%ߒ�8n������	)n��[��W�@� Uov5�<=
 �!�$2��.�Xv7ר�g�s��M��x�H��\�'"T������+.���K�����#�pVX��?]�u��[��m�aQJ�m��ĭ��hj��i�c�k&ڼ4�m�u���ztD���.5mF`m|M�o�`�^&���,�c�=�Mi}�"2����ʋ���4a%�bO�JԂ{�Wۮay�Q��+VXx��ަtFg�+fg=��F(��ȹW�56�i~c�zZiXc�ޤ$�D�YUla�Q�<n�ѝb� ��e�����1�,"����]a��`t)I������@Uڮ�㓴�>ZAwӟ5ja�L�ۧ[�^)�ѡ�	��Ht�ݸ�vB3�����;�T�Du�A��V��*�������-���N:�x궭��0��e14(�3(���jdvM���X��G�s�U��5�(b�KN��ȵ	n&+��u��i��C��ʫ��2έ�`��5%���7e�(�Rz��~��d�� `�S��QXּe��u��ɦ]����*�/�ˆn����#�>vg���"x�$=�u-�<Hlԕ��4/�M!��_o�;&�|n9��˱M�\}E(�b|�vW�	=�_���>�3��v�̌�},i,�浵L�r�c]2���Ͽr_B��%�	��v�P0�κ�$��u5:�H���=V���#�Kt�Ƙ�|>��6h}cE�f.�G�6����|�<ڷyE��/YI�Z�1�r���0]���A3��J��_71Zt1�S4=+C�����1�$X����x�y0_4Ϗ^\i�ˈ���"�(:���O�\��e�3�����"N[<	U;�	b�5��t~	��ҍ*]� �~	Ƌ8�\=�\]\��lڸ�O��lU0,�#��`��Ji��u���a`���	��"���k�q��=|<�ɋ=���;�y@�#� ݳZP��)�	���w}��T3$ҕ�ft��O�#+:�ɞB��f#��8�O�1<t'*��.�Mڅ}����zK���ߏ(�-k䬸�r�0Bg�B�,�ۨ�}V�ۏ��e�g��|�jf����<�D�5�v���aFZl隵���O
�E(4�ޠ�с�������].��ꍨ~��e0&�����փ��)�Ǖ��KG���s��4�v�s�����mT�.�n"Nh���w!jf
�w����Xz����ZԹ�4�.�x[3�o�~��u����љX?c�ā�8�v'���]ݭ���":�P �"�	ݞ'�X�����{#����j�h�)���?8Z&0�yaet����O�x���m���1�.��y��6g8�E�����~&����1��K�T��J[
]8�7����.Syq{띭D�	ӳW��)if�ɩ~;�*��vhy=<6Bo��m��m��6���ث݀����M��2��b�lף�}��m�X��I�8�]�g���2h�Pp�D6��������a��{�װ�:�H�m��ç�n��T��$s`��W�:�V4���0hMpF�eڝU��K� ��!V�:@�+��>1�r�c%��K��f	�wu6�@�<<)T�:��r K�^#�suߊ��e��ٌ�#M���úrQ�h� k^~D~��ԩ���<�M�7>]�V��������+�G��Nl�NxL��b0��z�U�8=�b(T�}�}�*ﲫ�i����'P9!��_��Z@:\%$cWj�˥�4!���I��&\'c�"�QJ�AQ��=��ecg褙gb�Y�+ҷ���Ҵ��Tx�ʐg��V;}GJ����R���B���p�$��'I��F��OÙ�@��o��wv����EGL����t��ϟoȮ/| ��DjV���uE���z�!F���� aB�"���4��\		�w�ts�͒��ș�)��m�fr�J ������X`z�:t��4���bN�5ed�*�&Lx̉G�1�������Y���E�EYC��r�h���Wr�8��N