��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ����"WYj����i� �N�7A!�@<e�]ң�;��5D�監p�.� ^+��Rk0;Õ\z�7PF���p�e��	��j�kdD/���1M���(���T�e+qr)zD���FWkV��������\���mk�*
`�R���	j�' �� m�cD���9:�DhT]�����۶�����i����ޙ%��d7ܷ��	�:���U��(�����#���wv�pFc�o�m?���<�δ�7P����( ��(�����1���o.O����BE�l�pSX�m����
'j�ߑ?�a\����3!���Dꁖ�0��N��I�SV�����q�u͟'.+�}������t��l�1|��}��%��ؑ�)�0PS�"�`���I�5)�"�;d��i�='R�X��Mp��4�zf�~o�덖vUlr��"Dt��צ�Mt�o�3�=Y.G �B`A'��2c|�o�V�憺Z�=!�������*�������3ni@$��c\��zq�H3��Yj������P��� eSH ��Ǡ,!�D��]���A}F&����vQzqR
_�ؼ�M�{�k�v�|�nl��Fi�J8KĨ	a^m����JRjt0��)�#6}w4��s�_E(RI�:�r����s`m���
Y�,�B���}0�]Hz�,^�y�e�މ����;S�fg�ozmyQ��K]JX�H�\�:4aTxI;r��m7I��G���O��o����������C����bDC���@w:�<�;��vA�!C.�uTj���^��~aŁ?>�C���v.��5N^������OBͅ����X��! m���݉���P���� ko	�b�f}�����@y\�	9҉���E��g?�GR:������N��o��"��؏�?7��X&�po�U��X�7�f4 ��qE�/�m�U�\$�ѷ�7��Eг���c*ʧv�̻�|d�7�A!YҼ�¿�b�VH$�~K_���勮��;�<Q���sxP�0��hϑ/W;�,�d�q�]���-%�>�ᕯ-���t3^ ��{i��>�E_O�����[EV�E�`�o��@wި5��?�U�� z���Ϝli��'.���O36Du���hb�q���C$(��VdNkU�`�mi�
_���9r %�'�(��b�Q����ە���bȞ�9��:|��ܲK�$Z(��Өr��Wٞ����ŵ)��NU�����3��-y��˔�+1!Ñ��i��'��[e��m����0hjv���E�	ymRGK ^U:AeΏ�I
��|x�
�)�8��-���]_���n�M���,!q�Aa��0dm8L��,�F��FI��]�9����&�=��1����xgYJ\�k,N�}�ŭ�|�7syӳV%H7z�?Xi�5I}�30Cž�z�ɢ5o6��WSR�`�Z��r�~B�ˁ���ܲ,��^������Mȡ��k&��|���~f6�N�E���\n���I��j�I�����JKNM�Hðl�Y���bz��K���|{v|����gL�R�N{rCk��z2/�v�����+�:Y���Ӹ:��'�OS�z�8�k�XfSOHmNC��1�0M?a}�.(� �� N��a��m�aE��C��e��)�(��fVi�7���@��h���
v'���x�A�C��EW�ߝ7�A!����l���[wZ�`Xhȭ��/؏d�٠�n�f�#�g�R]�٭uRd`:A�Y;�W�d����"�|�Z���(}"��C
wz��2p��|\�.�hS�7��ߐOw������m ��x�;N���p~Z�o�P�1bma���V3	[�p�ű��Z��,�tF�2 �ړ��/i�%$�be��(L�R���P��VK6S�BϗٙwY��I��� Nw���Pm�m���h��f�ySX�v��h�A��[�F[�qB������Y�n�����~�Z��"~b���I�D�H���Z��� e��<�����'��������Xҙ��u- -`H/O�^	��O�;S��?oK�(B�N������*F^�9�V0d��S�/ߌs��v�}��T:��x�bL��l�.�z�4�%&;��j�(�v^��b�ڌAF��,N^��)%&������5rvX�B��V[$�]A��
��O<
v�=MM�G�s�=RW��9n�R5�(�դb��hƺ�'Z\Q�8����ZEO���-�`��ꂪ��#VҔ`d[��[�5�h5n6ϧU���b�V��[(/�LퟋJr�Vh5�R�](s�ٶ���Ny4��m%I�Yx���>� E����z��.Pb"���$�<�@ѣ陙�O�^I9R-#V��T�؈�"�����n��uA�R-�8�-ú�>c�L/��VM�	��L�ۥSc�J���9O+�(�ne��)�?R)1e0=:6(GئF�]�ߋקcG-<��f��Y�L��vi�����h�X%�d@��V�@�d��@��
-�%8�$�8	�jg�9���8��p7td���;t���Խ��:�sAӄ�(lf�z�2!�M�s�|
oez���lEe �ȸ:�At{���kv� Q�XWA�9H�G,8�PV��ٕ��~��y�m([�e��1�i�NYPJ����1�+&�č[VIe�1��G:&2:�P2�nǀ���Mv�m��r� ��؇�*��>7!�!D��+ŻuV �'0�oa<��v=���`����SXBs��E+R��� XM�n6���Z�e�64{�*4+Ϫ6��9Ϡߍy��i�Lq� d�罒)�'���V�lU�)�t���,���S����:��(fԧ���v��c��_�d����G���a�A������RTx5�����׼,��8}�������A�O��/=�qu��f�X�g���bը��O��LY���sB��+�R/A�h��C��u�v"�:�"�b(���56��g+�&��ԃ��:;�!�il�,��Y3�جm~��h#�#YήO1�r��{w���yg~��i��W����X��*��c�8$�	�L� �k���vpC���f��(�Z��0�29�v�FN&�^A�3|�ڋ%~):�~�Wf*����*�=��؟1�O�9}�{��V�e$X���^T���+�ɜъF#�+;��@�16l@BDJP��z��1ߚ�5_ꔜ���w�GMb:O��kf��UԔ�| En"2��u7���B89�%2�e�%`r<x�W{%��]�!���e֊be*R6U�fY�-�;���=�8cF�^�3�<�CQ��;�*��i�㘡�R8�0A�!zG,Y�;�rS;=�P�r���_P�]�D�_��[^���xo��[ߨC�&�R�&m�n�}'�W:dB��q�� �����G'ު�{<�CL�߫�F��)TS���j��(J7��k.�Ej7���_H���_.-很��2�yki~㼃i�]>��l�Lp�Ph��s��f�V;4N����9o _/`Ȝ��3�ٍ�}�g��C�)$kP���xq���u��(ڌR�7|�p��d���;����3���`���!�W�?B��יz��&_ڿ4������Jg8�����z����2F�C�y`?��Yt��eM�d��4�&j�#�{␍��5o|HN��	 ����n�؃m�B�䛔?��rGn��F�/a,n�����ޭ��9�Ń2� c�؃�ɾ��[>�-tk�$�Ͻ����V�-}{�Q�"u�;�'�i�Ǿ��q������L��*���&CE�7}��&�#�Ր���q�/����پ9(��;��)�{����3Q���Y&���ZXΓ Q��<�3	j�i��捔�J�UX�P��@�:R��0���@��ҁ�ᜈزЯ!0�j�.zt�.
-�#�m������ d��	�7� ��?S�Va9��8��ƍ���0���3�V�m��p�w�N�&��/?�h���7��8H����;Ugݚ_�(�4g�;8�_ʵ�f���a�Y���.P�o�*�����®�ԣ���=�����ު<s�s��ChT}��°Rk�k�`����`��SO�bǬ�o�U�3�F4�dK�N�t��;E(O=��A+��Oel��x|��J��1W7��/�e I'��P�)��1��+��{�.'P�p�9}R�9y� �O}6�k^�GA)B�E$����p&�`���d5����`?���:U�jE�@ �O�~/��'	�`~vZ{*�����fy�I"ص���C'S�9F�8�ߨ(w�
,���5G0�X�)�
�n��^�+%�1BZ�f����_��R&qi���b�x5/��n�d(�d�ǆ�-t���*�4����o],Gg��� ,i����$(&�������B:��BɉD��1�+��@���T��|v��$W�B��Z�B�\�V)w�(¸};��F�60��y4^��21'�|�N�v{�±�r�4�ce�Q���F��:)�5��0���O?ww�剔CA�	0�>� �6�4WI�~��C�ݫT��%n-�Y`���Q���G�)�M����b�M��L����t���ϯ�Uq�v!�ܛ� ne��7����԰[�3���Z���Z.�>�B�;1츅�]b��$I1n3��hT� #��%ؒ���T�)�A�c�J�wۅo�^W��W�7<�8��R�ۖ �b��△��$^��S='�5*�q���)w�~h��(*^z���@ ��g,~��4�;�bD�e4�Y��o"�O��-�m�P����h�GR<�r��i��4�w�I�C�v�є���q�z<f��e_�FO+�/����)š���S���M��9�(�Q�Μ��B ?*�o���{�d�H��4^0Ǭ&�>�F5-!e�J�$�c�P�NH階P'�'�s[�!/wftD��?Uj����x����Z�=x� m˚�M����`^�.T��"��fl�������yh%�
t���_Uc	��Z�\�;Y2�#ݷ��j><�Uc�%�o�yF���no���0�<��M���(�b�e�.������a9�	u](�����c��xt��U>\�Mv{g@�1{b/�ay�D�CXi-�ȹ���|������	��/:�uF�y�ȥ�1D*&�p�����P��K�¬׮�q������pi!B/&5��22#R|��X}$S�DU��Y�f�twۭ����Ѡn{���\��AU⧣�HS�(O���,C�Ah��`酽�HN���-�E��1����8[X�,��<�W��$˓�,n�2���i[Q�@-w)E�}�:��֛ۤk�k��]�Kk�_�ݒ�2�w#!�f/u���[5р�Tc��옒s���r�Fsl���r�F�q�N�yx�BR/��/�Jm��#�U��;|���i0���+�&��=K�.C%��u��� �$4^�1�a�D�'[(�MFf�ᝉ%�ʱ�]���4�'�N�:�3��LY{Z��(a���`�	�A#��&7P릵���B������Fc����>!� t�~	���B?u��cp��'���I0���4�Ar���)�P�{�zyM���M�ɪe�ty"����[�*G�׳9�*�5��#d�ML�Q��0O�1ѥ��&ca��Kk�Z�F��W��.�4��*p���l��~$P!Ni�޲S�a#vV�8����<�`c�4��,
�<�%lT��=m۷@�ݖ=c䰝�)r%���V��B�h�˦����P8o��[��.�B��W+^���"6�V:t�X�?�V���p@9P^{���(U�4^��I��S1L3�Y�W�i��?�i��!�]]*�՟";|+v�����Kg��c+�hW7I�f�*�&�����_ ��e|���ʎĽO��OBN�U�;�m�>��/���`�*���e������@�~8a0`e��.�3l���z!Ҡ,i���櫾���*�ưydKs�ԡv����*S���塠ڿ��3�X�g��)T9��zz~�p#�j����:��$�<�ĤV���%�4��b#㫡�>�(߅d�e�.5�g+��eM8җz���s�_dϲEm�9�L���4�rO�C�ދ�է�Q�8�����6|3�~���.RAy���D�F�5���@ר�5e8�æsD&��v<��U)�l�z۬O㖕Y�����Ș��ÑZ������j�K�m��|�y�(%���QG�r��[Ł:� �մD�/?虒w�%�[ⲱ�5�䷬���A�y����J�����(EA�r�\�S���8I��
,�'�Tk�y��k�Z��ZE��JA2U��Q�7sa�$˕u��������쑣��\�Ǌ�Fnh�0�dq/?�Y���o�u�Xj��.��#��g]� D	̅)��Y��E�Je�5ب�[�|������4S	E\#���
."�r:��{	���Y� �;�Q߆+�I����J��J&���X�����qa�% qɑ�
���j�sاS�#\�������r$jB�%bWTƛ����F6�J/(�s^�*Z��B�qq��6C��g�%5��)'g#$�qCבOl:^D~N���4!�$�&�r��wT�e�̃qO9+ϝE_�s����̵�>c����l}���?�}٠,��
�~�^�}x<Bg����pY�`�H_�6�䔲?��t��(��{��w8�T�����v<�߱�_&[�?��O["/Az�9�ۈ�c�r�=��q
�RX�˳��TH��L�<�ٴ��ӝ�#8�`��)�lO�ާ^�N�$�3t\�s�ڦ��d����*^��f͢Wn�^&L�+�n�YC~Yf�/���*�
�{T�>OD)�4�|��?a�ڙ7e�(����^&�d�Q���%���0Yo9�֧|�F�f� /x��w,%�u�U�(�U�RE^ԴD���0�h��Ŭ�}mB��W��Y'bN�D ]�Ĺ|Ḍ�|��&f�������0؄��
[�ԅ/�#�M����_;�={�6�lȠc#�g�q	=�^<��Oz�-�K����==b	�5�q�1�&c�V�=^]?JW�$A���ġB2�!M�����Wт6�Q*fu��6�u�ǻq;��s��H��,.Nj�XE�凷5 j5H1}��$�q�4��2��x�lNi`p�cI�I�lo�U��>d:3A�(���-T6�B�D5�(лfy/G�@ ڭ������FM��,?��8��)*��W���-P����8-���4`,G��ĳ���z�i�}ѷ���Kg9� %��a�vw�%'��W�Ak<��*�P�������8U��T�WfW�c1Pj]��a܏����P='�~���0F���T|��\�]��S۱ˁ'3�����{��V���fc}ɉ8Y���az�:�2A���t�<Xڠ�2@HL8��8$h9���������u��� �y@b;?X:;B ' I�ҝV�ᰓ�C-dB�OL�iԒ4�
i��ىH�`1����b��	�Ǐ4�v�B������`!!SZ��ٸ�c�PU!��H9���e9���;�HPy���y)@ob�	5-C-�	-�T
��]/��:QI؁�nO�'A��O�#�5��P�a

�Lh^�ʵ�e��k�)���S�E�-�xb��-�i�VVl�")�~$�?"�?�'12
2T�ޕS��N�T���7��@�����'-鑯:@~#կ�Z��K���	��%-�AP0�X�E��̙��{}�1�6jT��s=#p�wQ��O2	H�72��'���.�W� �h;��.Lpr��;`ct���WʅC\�����M�J�{Q6ˣK)�5�Ou�D?�B�e�#�?�0p����F>�Q~�'S��@@;p�>AK��0ӷ�P���1;��P8�d���~���K_�ޑ�'�މ[i��s�_>��"�\.)��b�����њب��d��A�+���c>��m1GWۅ�l�&���&�Z+7a��c<8�QE�0��Y6�>����}|�K�}e��EH���rޡ���Q��"�e�����bS>/��}*�'�_�`8��Eh;b��"�NL���|.5��4�u���*�II-Լ��O�p�=�A>�U�8��f��.�D�P����n�;��Mk���3�;�Npv�N�4�=W�#R{ޖ�y%	���Y�Pe�pg�۔����E�D�u�Q07�=+�(�տ˻p�.a3�B̸%�q¬]�B�'nf�>�w��- gX:Ƽ�0�?dw3q��s��o�p�gB�M>���@�.[
��"����aB*$=�<��O�V�`̈�}��Y���6EB�X���.`��"j߫�~�YqDmCRt��m����3#A)��{hUz��eJ�@���q�h�����m�!�`�GP�B�r �<-m�^��J�G̽x̓p1�����y�o�<�Yjz�
����4���-�*��E4��C+D��ni`�_��r�Ɗ[��F�|Pt][��	n���_c��	�F-LnW��؂,r|�%�}N;����?O}�E���Q�10
\r�EnD��a��F��M\�'�`�
G����Қ�@!�9�e�&��&0�r�y�x�_�6�|��k��v<Y�	5�ޖ0d������S�vP�U#�Ⱦ�E
�1�>�+1�v��L���RS�hU�G�CI;ɡRȃ˾�SOX�^zv�Ɵ�e�=pS� �}���K�y=y�r����Щ�M�o�����0�n֯����?��=����!]�f�w����1��������>z�
ƨ^@�)�F�
# JUp�{��
��%���3�X,����`r�		�n=y�VQ�J:f�
5����=���,,
�K�-���)0���W�m��V�nV����;���"#|�	�����d�Zf܄t�A젬��s�P��B D�Z�j���)ؚ������=^�iΨ��w�9C���^ot��~��\{��U��=ϽI��Ǳ��eb��+�.�2Fe��ҙ��$�����B���eg��\7�Db�w�R�Oր�kZxz�Y����Ӥ���^%��6�������q��8�j�nt��RmH�����Gu��
1U����	�Ǵm!Ǜ�d* ��ˑ/��aL�&�vB1� �7�n�ϧ�-�$/�-��L㱚�
7���e�^�(�<@��8�A�>������`;�`��B��Fc�(����a6m�g}��R��;۸�'��z�WHDu#�Nc}���^RUg���i-vLJ�-��f����JP�|j��c'j �p��H�x8)�شˢ��0l��ݴ�� >���>rz��d�;S�9�DӲx�ơV!���KWQ�1�RP�+%�_�]񤂎aB���x%�޶�7h��җ���N	����M�*q��\A��ԣh֏-�����f�|6������ӭ�P�[H�p��Y�_ya\�;�⸳��#���7qC{L!G�!Y��4���K�!P5D�ꍳ��]������J�8��ضV@���C���b��!l�Os�Ix���:��87ﻠ��]gp��"٦��āj��.�����=���=�pbWrM�����O�{��T���lY�����l_ZZ�;�ADNR��kP��b�i��m��b�E��K�<�	t������C�SɈ�,���l����QO�0��&��OY�^��xS:癅�k7�Ve�#���VN�:�*UH��=�5�(�������%��6�o���.�;}��_m3�^^$FU�q���]�o߾�:�!]����L�i�ڀyy�R��I�����Ò�gF���4���a
���/}�����wf�nn)p|J�T,?X.u��J����k�!��E�h�E�*0��rmL����@i��L÷�~E	���� ^ $��u��D�������lv��а3YTiN�B䴫 ſ���;8�7M��An��z��a�O7���@lr4� L]�ƴ�oOM��t
9�&�}�w�xh h�S/~z���'�j�q�Q})x/���1�99�N:N�kq�6�e��h���z��uJ�d;��c�u�n�_�25�]���-�.��0f�E��R���<�ƭ�k��.W
�qY��g�>���4�{"m�*��{N�($�D�nd��1�1eܼ�~z�h� ����C���I]l�̂8B��XjXQ�ё�$=�s�󬺲����w9o�����1��+^��YqP:��+�I
:�c��.bH��;i:�v���1"�2Ѻ$�VS@ A[�dK�I�CF�����\��0H��Y*,�;5 �jT͓ 1(@���`���`y�j����,��@��Q��hs f�ٖl�t�z�����_4@�2��wФB���jFW�xb{��'K~�W�e�
Û�l&�w)1��A,UU@��N]�8�4�b�WU)ؼ٘{̸�V��9��B����b��ŋUS��Y�7DD]��"[��ދL�
ׇ긦QxF7�X�3�|&�_)@��%˕@�� $mKh�SpM�U�����`���c3ʇ=�V�3eV�y���#�m��Ǧ}�Ǹ�	I�2ܖ̹�h���IVQ�Ĭɢl�ֹ�q��D4��gҵ��w�[��&	�S៶�`��ɳ����؟�����c��I����weM`�QB�����V�p�e*c�z�w:D��F,�Diq�W��j	�� FGo8>�Z{��<J5vr'�2��9�)?����1����Ǚ��D�f-Ta��O�5�; �S��櫍�[�u���*�U8*��)���\�P�=�FQ^���4�EM�q�@t�u�c������Sy�4���	Z���t:�N�+�T���1��9 r]������L���� �ck��G��]�8�� ���`�gԔH�l	z����` �>��F���jT���g�u \��.t?�d�P��N5���5�`GH{�5Y�=gc蠊XY�jpX��Գ�Wo�:>	2Yv)�jjeHq>�z�s��P��}�~�ȓ�=�o�Vl"Pax/����R&�d�HA$k9�D}j)X�zhН8ۇgZ��!g项�$+��U�qh��9]��,�SB��]
��Ȏ��2RM��>ǧCō�%a!��`�$�����"����!��`�����9X����!����F�`D#G���. �3\9�&k�>CH�:��o���ǯWo�+�F��P�����D�8��H�oN�p����G4���(0�uBҁN4����䍠#��B�wD_�W���Nsz�)����͚g.�डY΃���zN3�^eesӡ�pT)��[��}a	�y�{�,v!Ky����F�K{^��i��k�t��Qt
���7��5(�w�P[57]+-L63-U�ҎҹR]�^�2j�+�/,EQz�b��	`v�{���N`����5q����5���GM����� �_vжB����sQk�\�5ECַ����s�6�{=m�9�$q�G�"�H����i(��^ ��!}i����j+��p����Q[��Hp���,JX#�@9m��tl�z�kr|�2�d��'E)�>_U�ە��b�BT�U���/Q��n��P3�$J2��.v�o��U3��:��)ܨQb����t-��={h6�2;5h��o�ȸMC0H�)�?N1��*��9��Q���yN��u���LZ��8�fl҃^�N�x����[���)D��ڍ�S�����Ն��K�}����	�=�طd���C\�C^j�GT��=��z��<��=m&r@�\�x�D{��� �2m�I�l~C��.�bc�`	d����N������w ^��DC� AvXlGnV�}�Fφ��\k8�ygwX�ݨ� &�z�H<t��ӟ^�)ݳ�҅�eу����B� ���4�*g硱G������8/�d�Nz8 �U�����g��Ek�Bo��\%�fh�4���ê�8� ������l��s6�~�g|.����}��X�`�D׏�2
�)���o�~��tQ��o4�$��+k�j޸�';��[��v0
^�5S�� )S��[�G!��Y.�U;��&�����"z��:&'=x~�ʊ��$����kEA(�ҕM1������� �3!Ǻ%d�|
��P����4�w����Q�{۳B�D>*���6�_=�t�� G��`�#ځ��oSEۓ�O0a9�{'��G L��2߼��k֢t�=j	���S����C�- B�I��хF�Lڂ6��*�X��.B�?<&��˿���I�:^��[&x���{_�^��us��Ag�� -���!�rN�F˹]��E����c�5��j�4&�ı���H��E��0�������]!D���&/2C` ��6���u��@�ͣ^�9��I���*����%�8#9�VX�R�8$3Mc����N4�J����,�~ۨrq�w�Q��[̋X*}����xWl�f�P��DFJ�UYP�'�7T������ڳi�B�2P�]6�������`{|�Bj�1Z�b��*0���������8����8�\�(����z���4�����e��ƙ�S:?>��:Wmk�H�����0`�8Z'%�Qn� R��P���q�O�ipt�*��**_�� �1���ߺn��9���c��y@!�9��"��/������p�!2�#���d~��钛�:�%��Z�.��ͬb���qU�8�������Լ���J��V+�Z����Wڥ��Y,8�����������#
�"�}��`vg�ђ�]ǧ�:p���
�S���Wn���6�����C
O��Ru ��O#���-M6�$�����P;�
;(���8��~�9�U�3&kxX+f�ĈQt��L�����g=��y�*��d�m�Яޤ���8�B�)zp
�{m�J'G��%�\�Nݓ>jF3gy���P��@�9�3�׸���u/���W2��G����~��Z��w�������T&*����A�����;c3�ɘ|;��R���:�A��UJ�s~-C�.M�/	�����Oqo�d�)��Nl4�Q�~�'��:�ޝt�w�j?\yC�gQ�Tq�(�mzY&#�^��ȡ |-��g�:���I�UHB
WX�����
�Y���r�>���$Q�q 0H)'+bh/�y�1oY����N)�..����R3u����:S�5�<>ݢ���
�}�c�n��c6�̮S��d��Cs�UP�_��>A/���Tڗ����&���7��k�X�j�Ciw=��<�s����c��(� ��R���B���ZJ��x=��T����"�����L�PD��@$V�<6��5@&�# Q��X�Z����~iU�R���`�07��� e���9Nü�Nj�yغ�6�k��f�	RO���C�K?~I8 /T ��/���v�Y�si�*Ki:LC�_�(e���2*��4-~��E,�Ԋ�Gl[�4��W�v~=
V�����Gqa����][5�<�Y9{G�7$v����m�Z�q�� A���d���ǚ�%CClɈ�(��Y�(u��W�uO���o!��e;)'e�Z�:�"e����B��_��:=��h��)hhi[�S�����m$1#�������~�V���e
Pv8|2]L�~�JR�;��(���8�.�We�yUp�R����Gj �J���ȎaB�o..z[�Jui�f�)4,X���#91̮�}����g,d��΁m�
5������\;�{��Q�:�����D�+�ٹ�v	�_�l?�:��A�s�\}y��ڜW^�����;2xU�(/�����w�rQ�E0_�U����+}� B�3�2�z�ު�5<�m��MT�(���e��/}�UN��Ls��9�me��J��o�cM~��SB5.�W������v+���m�r��x��$���J%���]>K����!�^7�%<�%Mf�/�'RH�lkW� 3&�׼������M��żʿ/����䳞���Ɩ��L-��Rz�h �ۑ�C�EІ���,UT�8xu3&�Ⱥ��nƖI��O��8s����VXx�!c1k�@y,��{k�";��z�>�X���y�U�\.�d�5��7�����>�
Nr�j�S<C3|���?��S)�,5�i*$B�_��Ǩد<���Ʊ��i&�I�RTʱ�^6+��n�(��jnD7d W��+��f�T+e��/���J+|������\}�F3-h�ؓ��֒�\l�J�����1��#�"�믇L
��N�<��� �@~�P]&�Z5{K*&[��w��L�dʻ�
�*��LԦ���w���VW�V ����Ӿ�I[����֋4�֚�e������O�Բ�-�����C�cR���8&���=p&;]��4�ؼ��0�l�W]C0#r0��ܞ!K)���(�l��f�am�m5�=QE�c�QpQ�6U$�r냇��Q�	�>p������f/ f��`�$qb�y.OG[vv�Ύgw����=��̮���}��$��m�3��+Ch���xΦ^�ɹ2kq��=@���h�OoZa�v�P�ڸ�컊�I�g�kM��I��d��� .�Q#��a	л������"���ɧ���� ',�tU5�?.='}�=˝ǭ<��(WctU8dYQ0Z���v3�w��� �����rh����X��@0pЩ1�_
㣒�-�cI�H�q �9��:@�����uZ�A	����He"��c�����:��1
�u�;쿨��j�m����Hʵ�6eZ�v}�*fל�%ɜ'��x�Th��,�S�!\D}p]�s��*&���u�k��g�B)z�&+h�.�A����1��sRw�'�_�I	�n��ds���n�B�_������������wdV��
��Lt)��^�+C�BZ@0�j�S�=��%Ә^Q�۟+�vd��[�R����ր������pݢԵ ����F�|�ž5f�gyu�G@����r��i��+��]ƙ�H]�s{�'�Z|:U�O�./%Y��"���0��F=�т����l.�a��yo� �5�c�:���d�Rܸa|E�8�M��UIG�^u�.>k�^u�jW&@�A������W�u	�����
85���]�2�1�j�nD�e^s*G&��'�̙��o�8��@�p;�������P	��	iZ���
���J`0�"��N:1X���%/� ,L���*E�W�vs
��[���&.���Y ���2��{?4C����!�p���xs��GJ%�*&�x��CZvZ� ��fGQ6t�X�?�~mC*kUgXDn`TT�9��w���c���Ùk��(�n�G�{�> �3	Z������ěQGIKy-Mf�s>�Ԁ��7^�}��\���M��㙳��Z饎��dud�V�>2�#N@�oҴZ�]�.=���\�>D��=ɜF��D�Шň-<�[*'�.�,*u_X|r5!��c5���'k��]��(ᥳ܌�b�G��&��Q�{�\���1�)�2H���3C�li�Ml�S�2݅�ؒ۠�V��h��s$���铍d0�,)]q�+���!E�w�Nq�3�PuVJ-V�n2)�tȥ Qi��Y��	�0}�+��Q̟E˅�%.� 1(��D��څ�6=Ù
p��	CϠt�	�4�m�K�y=��[�t�.�$��g��,W��|����֭��ug����~㳦͝|u�L�3�ӟk���/]�
=$O��	�s����v���˳P�0�^�@�uD24�Nm���g'��|��^��>�pOf�r�M����>�,r���bO��B���b��+�d)�^�t����W�mH.Ϲ�dS�����Vγj*��M:S�Ŭ:�&ظTZ�x|r)�Z?y�6��=:��/8`Uj������N���m�=��Ђ�[ߟQ.��vP�~�w��j�<�b�$���G�o��5�H�.Տ�>x�P����@����`�nk�^ui	����K�,��릧��A�쀧�K�e��4C�dj���>�3�OŖ	`_����-��Yǌ#�/��nO �.6[܇ G�A����m*0��#�0/4fƙ��Em��l��
�#�Î�Yx�Q�[@�g@�QN���xu(�O��=|R7,� �2$��+d�~�}�����Õ0j�AǢv,�,��j,
�vXo�i�*ʩ?��΍(c2|V M��.K��4g����J#��:<�s�Q�����2k=$�b��'�r����r�g�HG����3X}��ȣ"�<�;�)m��2X���S��q�<���_XD�ɦ��E�n%�zW̺��&F/(m��^�=�Uj}�4	�׋�no�����V5��X�� ��=@>�����!�w�u̲I7qL��ґ���w�3��m�<�S���N���C�s]0�+-��g��yQ�lD3o���� �\�P�u��y��M�!��ǎwܻ�~��s�W����R��ZS}�^Dʺ6ar.w
�j���Q�I*i���t%�i�x��1���8�՗�}��Ε〽>P7���g8tV߿�t0No�|&�%昹9#��Rټ�y�ӳ�k��X<0�;�Y�w�!�M{j��V6����1g6�?��&��"׊9��;*؁u��޸�CI0���E='N�fe�/��y�Di"�{/��;�E���+cS���v�mx�b����*HJ����Yz̡����XM)�]9��@�&r86���.ZBT��o`���-;&E)�mL����Z�t{mm���
�03�, F"����0:����A	��M������d������)a ^����g	�ge�=
���D1�c�_��!W.a43�˚an������z�uE@����a�+B���ǾЖ���!MP~��c�N̮�wBB��{j���*J�ײ�]�p�d��3��V@Q�<e�ځ��{ކ�Pa�?��h�G�� �F�C�M~�{�<s�S�������8%T7�E����g�Q)��T�ӗ�����z��S�L��!�7�v��{L���?`���
(�5z�J�g�~N�Tw� �2�,��2�U���$ɏZ�$l�i�yGi��Z\�jJ~��>�?��Q&���Ԃ�哧+\I��G]�ވI�Y@�s{��i)nn�H%����������_a��*W���gb���n����h�b�1�WO�dYs�[t?՛ʅIv�}��f�f1L57�<���+`��y��|�>�"����:�7�Uէp]�r�C��l��<~ŵ�����V����?��%,A��Jw�6�L�xA�e�?����n��Gg�e�6�n�t�p;����S⅛��-/Ff�kPP
w;'�N�ң�G:�R?{�E�?P�|V�/��h��_�����h�� �$��-y�Ö�Ba�4�ҸM4���D�Ƒs[,	 q�J�����L1a�*J$���d���]�F�#"dS�^��e3[��3��� �R�K��9|k�(�v^��b���_#i��L��:Tc���Nr�1��B�G��k���tQ��L�\�_��G՛k���H/��.7&�?Rb*G��	\X�*�!/�����{M�\�٩ۂ���"emc�d45Q1��wQ���B1�<N��=���G#�[�0h[��`Mj�Y�7/��ﴗ��{���3�[L:��
C�뙴j�
��=����{@d0�ڱ]�e�}�`92��X@N�]%���9t]���V��Z����~���px�T�J�	.z�e�����ykJ��GG4�(N\:4ֻD�Ð�.�ed!�ҋS��>?����vH��b���c@d-4,nd��}��))8��bKs��lĂ����f��nh5�W�"����&L�ϩ�-,�S��r�i0/��-���b>3��[���q+f�餫�IB��	�\����@��wj�~��Z�m�DSt�El,��{�2�;���dPx�Тm�%��]\����QW��ylOA��,�6�.F�U��:\�lm��on�������Kr���3�
+�+$X��}ikL#�[�k���oŇ(
oR�[ti���S%Z	(�W�l(r9�q3���*v?>�fv��A�p�@?�9��p
~��"�/���>1�3g�kHip�vgE�_�J����0a�\�F�Q�}���w����|�-�
�d��2xkÚ^�ɠ�s�Q�}�pZΓ!�ׂ��WգlMY;<#���x�
>�q��kM�+??=N��ͱ����jڝ����4WK�oa�LWԔ
�3&9:�� �g�EׄA�x�E9ǉ[7�DD/�T3C����Z�I),��~�
h�}?*�$�5�ִ�^b�<�T�"�g:?`:��]b�*'����Юf�9�6ppR{oR?w%44��?���,Q\�O��$�����(�n#>M�e~�`�����B=;�̃��b4�Htn!��w��h�
��Ԡv���J�\�5���$�_o�D��]`- ��ӧ�H��:�:����`��ٲ���ѹ1��&E�EPȗ�+���CW9��R]���or��
�+Q��� ���P�,��L/�,�y�0Ij�"
k8�m[��n��'��1��'��B/2�q��>y�0$������u�k��v>m�A_����z��y��L�r�4$��ٌp����5ʉ�*���ؒ�����㇅r������"�{w����t�������2L=�z�Ѡ��C���A&�;��I�ƹz�C{�H���(�[�B%h���o�n���Z�W[e'U#��xS�H���#���	�,6<t.��M|�a�%��39�x�S���so�Ҥ����Ko�ae��R���wAn�M?����J3<G�R�Vwa}��CӲ�; e	�@�ܺfY�+�H ��#8!�}��h�m$P>��!���y&]1�s�,�Ⅲ���2xm��)fI�1�wd�E�@6.~�ipT�Cg�R�Hr�e��K�~��~��u�zIK�Tj6?���7�?����
��?5]_P�v�L�	/M�ER|j��J�}�7Ң� ���Y�ݲycg<�z2��F�Ci?( � ��d��{3C�}�Fҵ5�U#�xt X�Uy`:C���9�{e�g�睖�}j���}R٩�J����Qڶ��"���8�jbjf��g"m����U�n�)�Lu�$"�Dx*,"��6�ժ����\�q%�����h�+i8lu[��.�V�ej�47�w��7T7��.��3^�_��u:83�5h@#�Ԩ���������8s"�@�`�h�tBʮP(�U����~�[��lC�BlDl��M�J:o$	�]��o<�	�;9-�t��K���	S����
��m��gPe	� O��t��>�36�p����'�A���L�N���c�=JȄ��z_v�W7Q�O�ow�[l�����I��_D�\�W E�<���������g�%�8l�R�=N��Vن� <�䏫�y]�-&�� �׷��5S$�7�>�|��g���N����N����u�G��G8o���Svz���~��/I�|�`}�������{�$-���ZI<7|�������iƑ[�a2�"*����#m���
��)���K��Ϫ�-�^�6* ��g��:��:*OR��y��"u�~�U����k�U%hM�0�p��Z����5L`�=��[�ӤB߅��4����$*l�����Q �h�Ďg�W�A�ǩ\�ϛ�S�Z��t�A7�d��B
���7l�b�!���I��`��^_Ai���/ޙ�x򰝩�Ok�+��EbܐŚV�u �����������3����jj,��t0�,����눿� ��5�9��3( �.�쀲�ݦ�c��`�Je�[���3�e����6,?����#���+Z�fc����&��yژ��k�����S��5E�a©(��6[8��ϲs�}5L��
�M:���#������ �H��(�]m�?����=M2TY��|�I�*��&�&��+���������?2�l�s��	��y��C6�ϯ��;�2X~6B}����d~���{�*Ҥ́xU8���&(����� �zX�'m�ʲ�j�D��u�[���0�Bp�ɦ���5�{�?���"��>�p�(.��V�(u�Ϫ�A����gD��%mՉ-���;���Ty��'���9�ܑR"�����S��n�{m�xμ
1�xM��$V�i�{�m�~^�ԯr|�w�&���<��ܤZ4���*�FAW��H�p�8��<��_�s�acb�c�0+Ɓ'�VX�X�b=p��.\�"��R(��L��f2I8%����n�|��E���4�r>��K)n9�j�����v�5__��6�K+�NO�q�p��]�o��t�)�i�9[�Xެ-�_�4:�<̋ި�ii:{Q�1��� B�Ԡ��q�)P큭n���ۖ���Q��;A`B�Q|ɲ,ЌQi�˩\e�wV�����O�Ӕ����2���g`��5��,��8��\b�$�o ����Ahv(���"nRZY�rNa&�4k�������DL�0tyͷ-xH*Я(�L(t��q>!���c�֝xH��$k5��*�� ]aϰ�]|E׋"*���9�g8a�bwJ|�'�
']�e��.��~�f�o�h����eGRE���� P,R�ݨ&��&0�uj+Nk�|��I��ʝ��|-3w�y�3�"�x,w�z�9����T��k��~�t7�
A��<���h�(@��PHt�E�;gMT5Z�c�f<��<�}nև��.FX:#�t\�?k�GC��
�(uPZ4�$D��4�qߩ��Am=����v�z��A��A���q���{
�g��^o���x^�Ώ��gf��)8�hj51�ｮX-ە-�&ĝ�g�Nd��~�ΖL=R�Q$�ϰŏ�2I�FY��M?Hc�O�vC93�$8�H�{�?�����.#�7aI�T�M��(�Kj�(/�H��l��LA�	�*��#������9�d ��@\��~�WM��n!������`Ŝ��|9a����ʴ=��p�)���I���Y�.�4�u������jU� �4Z��G�B�89xp�	ٮ=\�'9�8��?c☫|����W��MmM��	ǗQ��`ի!jA��sԹp��=*bH������e�[��9&�hB.�#�}hxG��'��UR��ϐс���e�֗Rڜ�?u2u�r��l�:q���m
p3��w���A�Vȭ��l��3�S�}R�Z~TP�8_S���bm��F�����ќQ2Տf��ڈ�:��6��>N����!C
��(T���ޣ��ߋ� a8�,�<���������r��6`n{4�Fa?�!pmRtk�#$Hv%w��xx��M��r��c�-$��G*'�̀�:�T�,�U�w,c[��w@��)&h[Hg����\2O�~�zXŤ�� �!�'�#�#)MU�Á���I���  00��]ϯ<���5�-�;�8 燼���:o=g�.ؽ����@	�O���C2��M��e0n_Moʣ���0wT���`Nb���)(�Eg��)�J7�eM�����M<������ڭ�����O����;QR������Y�S��-��U׋��of-�P&��	�P���������B����R�	ڎ�Y�c"@$�/7>u�e�s\�;.}���~v�+KG���8Q����s�E}���\�θ�V�]�6:Ld��w��Ǜ
l/��a*�f�=��Ck�O��G\$���2�w�󲮚��*+�ݲg�}RK&������y�����K�i�ה^��N�-�ҵԭXL�7��o`Q)->!��z��e���	O�|QS���*��p��� �H)����RS_'U���]Y��iB>�q�&Of`10����Z��7�vY<h�m�Y[fӑ�T`!7�t]����;�p��J���$��k��.��5-����Ѳ�[{{i�K�B��X���Ol���r/��J��d�t��B=s���t`z��W����[��g�Q+��� U��sW�<>4{i�	�0[Ͳ	���O=DgyO����ߩٔyĺ�DWz��`��e������ܽ��8c��{���B�o�l=r� �q����r��O�(B�,yܾ��B��S�;�U�ғL�7��_ϛ��5���Z�CCf��ftQW�l�����I[��6�o�t��_
����@��jX��x��~���E�����!����;���k�E��Q���$�Q/�*�P&8�-t*�M����7���˫��i��I^ֽ<�M1�JG�A�\�Ө��oh�g����f�I1��(S