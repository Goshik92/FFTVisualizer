��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn�}�SP穟g�b/mk�p�u|� VNY��֞x�u�ׂ�B>����ˑn�+�ϒ�%:➄a��G:L�~� M���SM��
���lJ��$o�d ۪�7%Uf�&��C�6n�z�
`�i7���.X�q����e����> _��N֍�j��p�.kK��Gc���(j?�B1�Q�d,3�*����k�khy���Q�p��z�cU�͘r�?�R�z����2}�Hz��U Ɲ`�<S(�.��_�b��/{����|y3[&�7�*�xg�NC�
�=h�?Z�?!?��fp�,zK�k���i��-%@��iY� u�Vvb��e���d�\��֧������w#��F#��*Zj<��n��h�����kd5TL�y�XWB�6�p�ܘ����-��ޝБ�08k3f��X��+��=���]}x�+��c��;����ox����L9'F %�(G�l!@U���ڳ��>�p{���gM�����?>׌�G,�������L�כ��� ��M6�Qe���y}ۓ�G9y=0:��%FȆ�	β�F޸��w�6�t�.L�lT*�E)A~�<��iS�b�,d_��������WI�����7:�}��=�1Y�������qN�IdƖ����[���P"��A��Z= �w@�K`��#N�$��8��������㟞� ���$>��=gi���]�����#�K�//�b#/���s<��?�zְ��W2�7�'�O�b��`Z���v�	\V�B��������r^\�r�5-je�g��4��h4+�m�������@s_�o0Ń�9�.H��6i�� ���*�}��S�쪞����M׹j\61� 8j(���sm�opw�~��@�ƾ��������6iW�\���
�F�n�V��|�2ŎLU>�}�v��L�3���	UL�%�,,a������e ̅�a�35P$w�hq��B8�CyP�,��os���U�;]�G��ѭd��00�c�ڜ��bA�$` kl��}I�pL�� �>�@8�J����씴R�_Z�e��kF�&@�a%�9�>��\�J��ـ.�Q�х�O�=���J�<��ެ=s�"�r�	�@s��G�n�wL���k�v�S�I�$�>��;0��	ɬ~/�����Je�l3��#�(��5W�Vk2�1.C���T��}�>��.|)��q�C�o.�7�\��S����o&�D)�,�����FFx��,�B,���b@meB"�!90!�V��K���x��� S�,l7��&8��P�_��錢	�̤��[nz���K�3>:�C�@أ�62��|�'vND	�qc�eZ�y�,A��} /I�(>��������>j�Z��۳��Fe�$;��]���0!Nz�R���3m{�I�� 6���!�ҀD]��H�v�r�(��@g��ɕ@�)�6C�pn��`�2��~WW�u�m�͘�H&wۓb��(Ƀ��xc��m��>�����:�5o��Vma����	w�e�^w�l����l�Cz���;�Ι&ƩOj����i�P��F����Ɠ#4L~^o��E3ڜ����#z�}��J�A�ߡʊ��2sk�0k��l�`��u�ݞ.������^��a��I�q1r��}c��\] Ý��"��X�z�ʒStf�_`�$���u�	�jٷ�R��A����m@�N@:��dJ�>%�R-B��rj�ls$�4�3/��B��A�f�_CƧ&�e��YP�Mp���P!�N.�}��~*�ӽMR�}��yu��J�:�
���5%3s�q�
jK%l���)b���S{�ʋ�ekD��L��Y�)��6FG�66=�}�'���sD�;-tU�/|�>��A.q�sp�a�uB�&���������_����G�.#�t��!='�ը�;��A�]��~_��)S�f�����a���v�49�x)� 9�զ��$��>�L�B�:�p�����u�cd�e�$���g9G<��Z����:o\���B�WzXX�o�����M��@��$�o��$��\_$P��n�z��e�"Y|`*��Yn8*a\�t�N�$�j�8�^y�ġZ� ��#b(�II�;�R��s��O�Sl<ȥ
W��ac(���w�>�'#ȳ�d�������+��BE)��Q`b���D����G���
J��v�"���}�>�nN{i�Y���Z�Y&��"(����P#)�ޝ��^
���Pa#U�e�	G9�3�I���걹�V�֞�8C�W�iV���3B�+�����HM���D:���lAǑ��lY}w���s)�������6�s�u;� �8ã:��:��(�^ͩ/���_=��8�(�r�#�I��A�Ru�����N����^%]��\���bn��Ybj�����;�L�d���&r �i�B||��I�Y�Vc]�(���x\��Λs�a4�*ˎ�vO�+�q��
�NWI+��˫�>3o��V�t砍��u����(O.���x1��R7�27C�=/zk;�c߻���+�5�'�B����F$?��.�5Lr� e�-��D��9�M�<WK-|FX�.�?�9Z��F^GZ�jÛ��[�pf7�5$� �ؾ�K�f����ɱ�\��rmƮ��?�놚��3��~�$W3r�2�7���x�5�ń�0=ͤy'V��=&�>�e��L%�v�h��t���qh-B��I&�ω2>��ʚ�����}�L}�9R�;�Q�ο�5���? �=�ף܀g�W�R���q��s�Yʯ��W"��iΡ7�eP����:~:�8�~�癇��B��4��}�Z���~� �8�k4�s���e"VM�<�j�7bd{Ax{�<�2�!���x�w>5�h�\���V�h�{VX��9�����g���~7��Un�鲕�V�}ZK��,)eiw3Mk�U*�
�F���:��&��:�M;f�EʤP�;qk
���q�]����5S�����y]�TRc�1��B�ￋ�Y�|�
M���>lZ �,�n��I�Dԙ��nh��{֚f�a^��F���)�z��AFHW�9��:��z��$=��i���g�ؠT
��j.�L҆-���+��-#�s�W�]���0|l���T�'�'gMp�&��`��i��	��o�D|RG`�2�S���4G�����r����l㯭x6����f@�z��	 ���ыe�xk&�ꊩ�_��Ӥ�k�Pæ'�ыQCU#qky������>mC���`�����t�!�mIP�(�]��¡��&�DObeh�ud�
���H��v�v��,�Y�E)��?%1\�f�EC���
�#6��eDS^�p��A4����+��rtiBT�WOh� �ڻq蕾�;�y�)�}8?m1FM�D�F_ޟ�|���)ԭd��_��p�۰���w���7���8b�c��NЎ'KJ�ǵ��ؚ!8{��Ar���_yd�f���IY֓|�,�2c�M����%-	Aؼp�x����P< UZ�1�6z�B����{Rrұ���j���}J��SID`s{�a��"�U�L�~������㵌���q���FF�t�_�K�@q��Lρ��>�S��`�53,W8*�o9��!�Fz��*�������C��vfHq�,���qKq��H����#�aˊ0�(t��r�!����_�ؑ��)Q�]{��kyXԾc�(/��JX��$�.S��eYI����g1��\������	6L��b��ٞ/0|�RKC�+���窢&��n��!�x��0����-i�L��W��ֱl�����u�0���t�yR�6ͣb�kHy2N����� 8	�Q������2����2�W,���&-�p����dL�JK�����4�'�Y�ܖ�!�e5͡�{��͉�-a���6���i~6���H�m4B9�Ӳ����u���9}�,<���W��J���OK9�el.�1���H�����{��^��`��[�d)5b�K� Ӥ�TD���$�����]i�P^]�	%�@��:�.P����S6��N�1_�4�}�z~Sѻ<;ZF�����ر�h�2E")��E�-��G���c�Zr�]N�r.��w�J�Z(�I��ɦi���'#w�&�nlzml%�'v�I]�q�g=�j����� ')P��K$O[�k����R�]Kq^V�Z�<ڄL�
��go6��_x[:�}�����(_���H=��嵅���:��s�؄�=�-�d+
~�zXY{<�n�YÐm����{O~C+Ah��F8m-G'�t���i��z̐�d)��'l���〿��U�4���ްֳ�զ�3���Hʭ����2Ϙg ���4��Re.��h릶�Ȅ�+k�_��/_=��~1w��(�7s�=�z_�1���}�H��w�~)���ڸ9-X���Wk��&���f~��C�gs�'��Z��C0`�؅O���[ҳ�1����$nh�������h�*���ch�:�E�����e-]7-U��*0}�Ar됃f�}X�]�ք�Q��@<aÉ3���ۭr��5�T��#2�O>I�'yA�7ژ�Ƹ��ҫum�܋����Y�Y�W���q�s�+�(���W���1I���w-�e�(��$N���x� �b�׮�M�!�<u�"5��/��g�S
]I�ȇ��L� UBޡ6�]x���Lxut�u����ƥ��@�uh<�Jo���2�̘����p݀ue�,k�:hG����9��1�G."}�T�*F��;��Vy�#�].�[�0��&F���f*�-U�8��Q��P� �'��v@�/Z�����W+�{F4���4?�R���6(��C;�LW�sY�SB�u�r�����ϗ�M"�J:�L ğ�64؎�%�Dm  ���u��{x ���B��}� W�^2@���Ll�I�EE��T薁q�n'�e���47�0j��0=�ۿ��>l���W�z�������쒚��e�ޑT��BDz��`���k�C2,O��C\��q.�Xi��x��#ur�=ܾݷ�8�V��fHI�..$��?;m�c����Jf�����m����k�|�����7:ڽ��۠i�ӖK!���Aq�/?.��ld]_/���S� ��}�}�A�g�Ҿt%�R��t�	��ss���~gi��#�91���L�p2��o�	���7��"�'��{n��;.V��݆�Xٸ�a��\X�90?2b���kF�t���$�9�/2 �\�a�"��X�M��^6⑺��[��d���\4����1[���l��wD�/�Ei&�6��s������B3>�*-��w��|O�)qE{�<,$h�;�Qi��}�;��}`�PP�̓�����=��Ś]'�� �9X�$�1��5�?c�d���Op7���p�WGg �sydr����Z��E�a�d#�[�c���Q��=o��UB',���+9p��f1�s��3 B���yE'F�!�����)ep������@�J���;��c�^�i�~����m�(gE�R�0B�r���'�f�~x���	�v��km�c&��
�� LN��{���M϶C�-$�`�_�Y�=U���#
L��\�OƢ�&+����<����!əJ��z��k�t������3F�vk�� ��
&���p8��z�f��J�wy��	��G5�T�$�ɝo��M�
�Abu6 ��C�7U���i����Q�R��ۺ��2�*��*=&IPi<s���y:��j��P��u'/�L�|>��$�GN}�+6��#5�"!Kj%��_ b�m��]���օv8\E���-r��J4&W��zIm+TA±�
�w��znetu~O��o��2���$�G^�#<���	6me�Tz��w�!Ş (�-�W���ĎU"�nE/0��
"oeϫ���h�e.x�b�[*P׻цd�fdyሚ3Zx�R����_{��aen]$"�� �	#^����� aF7B1x��C_��)-:tu�\0$�������7xے:?�3�W;7\Q'M���\�V
[4�+Z}� �/͌��*�ƳǠW|Ї��T����#fB3>��z����<����;�Y,"v������"��D���ʏP��/���=*#�0�Эד��GX��:�Ffq�g�����/hɹM���,�աj� >ּ�7�{��!�C TX��<�,����B2�+�i�V!DI~5 L�2нQ0�DW[O�Ɇ�w�Fbq`����(P^V�o������m�"�D��~e6�Un�ߑO�	}��F�W�ܠk0�� <A��!,��c�v `r�M*���F�H4Ss�qf��$�~i� �S���<�&��Nֈ����?m'����iY�|֋ �
^c	<T1
��[f�����7����z�ɔ�ز��*��Bȳ��������j����މO���@�$~�@K}ᮕ&E5
��ad���Ύ�u3�;n.�h�n	� �����
�,����t^e��0���5tN>��x�!r0�|;�pLSC��]�a�Φ�,�1��</G!��h�	ʞzMQ��1g)a�f
҅��}�
+Hj�7�oN���gDN�"�q^�;�U�?�wu���b��h1��Q�T���v8�Q��mQu/�;������D�xj�����v�h���8� �op��5GtR������p�q~4.��@~P��Ԗ�W�Mڷ2�����is�w� ӗ����o���N��(���6��·�+��Q:��m��}��P[�������i��������[�^�?s���������Q�P�j([����s3�A3��;�
�)T���v��)hRh���d�EK����������2J�OI�7%�aw�]te|��UF]�LM:���Z�W�����dH���tJ*�g�qPG�Џ� >[y��^��׶��齦!C���X��y�㟤ߔݔ?���{�G��͓;��F2r�2��U���Y���\�_�<�m�X�v�N	�߯��j��)�ix8�ϰ��i�����k�!�W8/AO u܊���N����#{�ɥ��4�6ax�̼:�4Ѯ�ފ
,	��RcP4��f�T���,�4����oR)?3�0�b����95��[- �_e�)���p��R7DDW�%�I4SS&��^�"��P�_G�����<Z}#rg�m�2UĐ�q""���p��z}�A%k����6���zF�R_���eF�ϔ�)�=�n^)AsR�ܰ�3�v��^9G��N��W;����?�7�Dߑ]~R���������5R��#�9		�j�#�����\i<�"�බ�=�ء��/p$�i8���Ԡgۯh5*l���,�]_���!;�T�fǦ��M-������P{��ewsW	;���hu�i�&Z3
�X��"�����)]�2j> V�M��o"�D�_�J"?����G��̋Ć����TX�G<M�qe�}3z;�A���̷$n,�S�JᳪF��cG�����H�U��{Vտt�StS�l����眊}�H��d����K���-���%'?R�/fx�Y�G����,+������ ����(��b=|UN�50@���~�};\+Ӂ������1�`o���Ԙ*�C�Y>O��ZZ��'�;�[�|^��I��r��� F$�hk��so�����Nk��- ���x(6|���X�#��\q���bH�t�;�3��H#�U�u6r(>�9Ml�79��)W;�s�B�?� �6<{��WcmX��M��1�Pw{�F4�#b�!I�r��N+R���H�튗��7!���W�,ؚ}Y����*L��:��X���Yz�U5�ƚ2N;&��X�����G$���p�fY�\u���3�,Īlg%Fqb�LP�J�Y��d���0\?I����5��a�P�Lu����G|Y{v
�T 
������<hEՇ�r�����gl^H\��4̈́���
��:c�Z3,���~�6�+�����G�;%{ N[Z-��K�OVcX�����	n*�H
�)Ǫ3��=���~�Vh��{�j��D��ϤaQ��یp��=N�0��Oȹ���E������@K����N>l��ˏ��C�Ӊ��!�p���tz-��(��"$�e�V&�`Р�������[d+���B�n�}�������.w?+��\�V�Ҁ�X��f�"B�P]�)x�����2S;���0�)�~��=^rB���O`s�ls��ͫ���nI�W��<��Re	 8�(�8>R�.��(Р~�j/a���A�L$�~��j�=B�'�1�C<��͋-�}�+!4����w���yA
����?�S�����f�9�%�b�U���|�.�2�B9���t�q�AdM��N��{U]]B@I`|��<s�@�.
��4�&��4[���b���	6M��b	�M_A�s
�س2"���q�����7�|�g��ٲ��� � �ha�{w�⚽*P�E�S:吭��/�F��|/����1vkm6~Й�Hܞ8j�#j#��'9�-*��)���5&A���`��0K��� ��K`�:��'�/T���r�r>��r�c~��=e�.���	ٓ��9�T[̀���^Y������,되@�t����x����'�~��8�{1���u7�C�U<��O�C�h!����]Ų���bUѮ���@A�"�x��ڛq�
�z|+�r�~������F��~���W�ox ꢺ
��N�>�L��oLm�gOw�-�N�:~:;'*{����Ӌ,\{�x�Rl�AM����'�|��8/��܈�kɆ�6�f�O�o����y0�>)@ƅ7s� KR�z"�J��@�غ4���Kt�D�@K�ԉ�e�;���)Ek�*��V3�N�����-1�3c�`������4��R$=,�^.R�рPkA>X�P��֫sPA��k=F�:���S��pX�
P��ʟe�0ƻSKu;XR�P(������38NEL0r�Y� 'R�����L��^�'��G��������6G��8�`|=�;��oOEX[E9��e򠁯��\�;<�dL���$�ʋ���7Lw͇�����z�<C�h1b�1�!�x�RB��M�	�.�C�	�;������tuL*�����'��M��:����;&�����6�E:�˂��s����mQ���wC���ӭ��(��d7dZ32�������D�S]��m��yU�:�<˧�`=��c-�w�H�8���0���-���ɑ�Z��п� �&s���c&^}�V�-�s�r��-�_5���;-��x�GL�M�6$�D6���zI��E?M��M� y_՗5�a,�j.��2�x8bbX/�@jt�����x4�c����^ދ��A�(��%�g�8})�Ov� ���>�K��:"�>���z��Q�Q��XgbtAN<�uX��'
������ԤP��Z��g^��U�A����WN��R�x����%x�3��6&��a y�����TӒ��'R��U�:W��*��B|�ӎ��"B �.?��z������=�$�|�~��
5��Z����" sک����|����OӃ��w�X�Be��mzp����hN ��g�O�u� ab�ƣX�ml��z�#���D�%��iS�Q3��fP�DW��.MW�B��ArFd��L���u���0�b�v�ւAa���g�[��&K�Dl����Y�^��<be�ưg����3ֶ�!!�Ւ�tMD�L��<{�ٮ2�c]8��	���;�zȅu�R����D}���-���%$�z�i8���x��I*%�Z�l��]t�N��	W�/���]s��W�䉪������!��ޙܢ����H �m]o�10�w+�H%PM�M���f��s��1e�"�Oi�}N�X*�Ix�j�~��ڕ6 �M$���ݓn��C�]�$G�yr�Q}���B��� ��e�w*����X��P��1���F1ﻊ�N���!�P<��N����j�Xₜ�09j�dZ�۬Yb�����t�ɋ�P9���R��f���dH±�P�-��lx��|�������EU����Q�\�`�UD5�a⯷Տ3} R�L ��D�� *���G�-:��:L��E�VW�}����VgLsb�m|��)�\�Eg���Ǯ�w�i}`,���Y��PKI���Bŧ�p�8��)�r�B�`���X�6E��}�o=8+�>a�0X�L�l���v��E��@9ǕK ,��_�\ނ�Ji�Tr�!A�3T��e��`�3,\μ��2[�p��Kf���Xrk��E������I~W�$�3�l"$P&��
�3R�����Z�	�$Mc>gɡ�	n@2�wj�1=����0�1-��q�A�M�+(8���,�W�4w����I��	ҦQL�_�s�2�?=%�LP {?�xr�Z�Z���׊^�7I���U�.5)Do�2����HЅ8p|�K�e����q �r�K�Jޛ1aN�e�-� F�|<w���J+�yd�#�~���*���fE�}�#����\
h��S A ���[M���7q|8��S-�	z��2���Ҭ�����U��{1���ǳ[�\Q��PyȚw)*s���"� �G#P3*!�I*cG��E>�#���5I���`�`m0@��y�P�*��{#���/{NV��Q�q�����M.�4kg�YN��&�V�d�Y\s�������1��� �	�+N|�T71|���!�`z��&EY<��\~N!l����+��Ν
�Ƒ���4?��x1���\dy޻�K��H6]��)ea~��DB�S`��~���hJ2BFǹX�ΐT�����G��3�z�1W�c�'���G�Ir*�V޾�z;�A��^)Y�9m��X�̞�=��|�=�3�<��ʝ��9$�����
�AR�ݫLB��o�J�p�� PT�łXKd6��3x���X�^�g�Hs���~%Z�1�&J��w���U
��,X|����(R��*�g3�I&$���M��t*ga�@�s)!�A�u�&��>wL�t�����bX0Uq췯yy�V�G�Q��'6bq$�_�W߶@�S��5�<���3����G����:�7���Q{�[;ɀ4c�E�a'����	Ş�I�Ƣ���Gy�>�[;��I>�3�7y*=�*<��s����څ6tm���+���NW�H>s'0=�\�B�o�"ɭ��?�? ������b��XT�@��� } ��oV���9Z_�څ(>�F��i��Em�h��w���y-�ǋsq�u��m`����9(���3;�\NQF4�5�B1���ęR rY&���4\��s��N�������j�H`�����H:�|�޸�>��X�9Q�$����;����Rs�:s�ŭA�R�mfp
���\��hO�Y�ajME�&E ?�7�OHrO�y@��+QKL|�ڟa.d,u�R^�3;���7V_W+�q\��O��N9��y �zx��,�����A\����sJA1�C1ܐ�)��K;<e����C�$ݛ4]X$��c��J%��f�mf���(��5��<��d�k�K���&S��e�O�G���`��N���p�q:�8W�Pxth�Z�!C� ީz�s��g�M��#��HI���Z�m�g>�ZD��	���>wD�C��־bs��L�Ѵ��H��g������7*�"-f�m3	�	q���D�,�5�4e���.3]�t�'E%ܕ	Q���̯��;6�O+�E�A>��Ԛh{���=�)/�� �SY*1o4�[�[!j
:�O��@.3���!t�4
��;�h�ZF��(,3���,���JQ�~_���C��ݺ�n/+��C��sO�p)ٕ�?� ��Ju��p����J��?��aْۣP�=��CGg��A�Oŏw�ۤTn�만5_W�h��o	 �+�B������>�z����;��h_��4��������dU�>e�|����~ߛA��1Q_u�L*�Ҹ��s�sR��O>��G���mI�		˩�w4Y��͗(�Urb�w���G#�9t^���Q�+y�E&��g�����c>�<x{��+�s��"g"���Q�!髌޽��f�D���8�*碟�9��
��w��wm��XZ1�ͯ���ǄAgJ<l�W�[i:oj������i��ˠ���V^�o�^UPM�I$Υd0좵�7X��Qn�6��QM�G4:�yg@۫ eq+l �'��&R��
�w�R(��X�f��Hs�}��-�ae��w]���_Α]�ފ�nb�6���%j��*�FP���,���L)�foS�)��\^�X [Zn�Fv �b-&
Fg���N�FZ�Z��ϕo"��@�"z�i,�¤��"���i�7r�#b����-�d�	�p��������سU6�_dY�
��@j��C��Y�칆T8XTn�F��M���y�ګ��Y�GK�{HN��c���|bR�"�,���_x+E΢q!�q����Q�7Y��m��!iYC���e�$9��}�q�i��ẘMW�fW�iP������Y�y.>�_�~d�����+r�g2eqE^)#��m�׉�o�R՝O��КYq�4�!wER��bT�k��'r��̴ ���m�r