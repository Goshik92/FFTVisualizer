��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|۶��-�E��S��;z��Q��8S��fʹ:9�F
L�~Tbr�)	E�+�@|'|�;m�
�K����D��T�J�Y9��n��nw�,����2]�X����y�\V@�L�F�� PG&�O�.vCu$���N����]��\$�Sg�� ٤Ē�����#��ӓ�=xy@g f뀧���>�[k�e� l�`L0jY!�M�sn
��rHo�L*����!U�D��t��8�N3�4�$'X఼Z���%"��� $15�x԰\�i��'�p,�7\dX��K'h�)1��#4 ��7C�U��S��d�Y��ÌV/u^����a��#y��3���z�4.u�x�c�>M|<�s�/�s
��7~�4�%L8��,��_�K�I�3:�|�X*w�~[�)]���F��c����*���&�� ������ Q7�өd�A���!p&��׻
��AFo#;�,*��S��i�E�D�ʋ(�����C�Zn��Y���j�(l���޴�7���6��^U��S�G[L������]�i ��B�M�Z�2��%ί~���r!��+z�0�f��'�����������4�x�1�S�$�'�UA���!j/�AyMZ,��󆠣p5���װ�� �6�u�����e��~[O�[�5����?Ei���.ru�o5����4/�9�נּ�0���"m�+O�©��_^Iz��{ULc�Z�P���8V�����А.��z�������Z>�#��TL��e�8��k��V��g2�#��t�)*D�03[{[�>e?A�����M"B�����-�D�K��=�6`5:�`��<�8�S�7n6B�*��@��*P��6�	�?qH9�����EF�r7�:��ea����.�ڋ�Y	�ϴ��I��~����x�[���k���J��hH��D'2�Z��e�4�_v[�D��Іۙ�ŷ�"��9EFQq��5�K������5�&8��̞3��8h��l�H���`A2Izly/�  ���l�ܕv�:�%�>Z�����U�$D�c�����&�s�Z�/�w�J�n�c}ԅ��>���!�6�kF~��h�2�*��`[Z�n �L\�tu������H�]�0���c>���SyW?��Ǩ�q'�Ą�����T�"�^�)��81���ZjY#���͘����!�RwÃ���۟�W�`��ՂT�1��`����M�?��N'��e��Eb��Y��̯�>>'D9������|�猞�	��[8��w�:�Vd�ok���hb�v���0&_X�<� v}aMɷ����-�-&�&=�9w6�=����Cg��ھ�@�t̉{�����#8�V�f/x��;=D��j@�L���Q\t��s���a��~��G�O ��F=Ŀ��Z��.��A�缔fYZ�&���`]�x=��CRݪO����5�mו��v����e#��l�����2;��KǃV�Ԝ)�s��}Kb�$,ܶ�z��U�j1e~)��49@/{-tƃ}���-��炳WPT�넸W�*��F8m�ܦ����Ճ��H�w�f�7��m�ZM����6�7*LXON%�\���%Ŧ(|�SVÌc���+�;:[��e��%���f,��4��q�;u �C���pO'�A5�Z��g�}�gg0D�1f�/j��}>�:A�����`�+�:�ǏLI3�Xk����WIh��I��y0��dh\O5cB�4�l�2�F��ށ�]�,����z������ l������d�223~�@GL�S��f2���L��m4Ƽ�����?k�Fi8��+~#�M�M���GG�:c��Р�>�7Mf����<�E3v�\�d��d���Rp8Du"�Iwq
=:2*φ�,��lZ).��wXê��f�
����V@N�T\}��a�q2a/�1ɒ�_��Y��pԟs�����R���O�Vz��
jG��R�GZ�����2������l�2�yF���3�ֆ�ч�����[c��r"���i��n�ū���V���
����k���iƷ���o�Bb��#!=����'E��g:)��_��I*����O�h�-|���Ys�I���
;���~/4������Y8\�\��ђ ��ߌ��$t�!:�!͛;�.���v�P�g��ze����7�"��u�Ƣƒ,�ME�0�����/��2w�#��*?�4&�*:��������u��B) �^���_����i �&l��CX�$�ڿ��Wx�/E�u�@8A{
��T��1Sh�HeB]ֺܳX[Ϡ���#�qk�.�G������o���az	�N y4=�U�~b_�s�4:��~yB�gr4I�D'�π��+��J��Ț	�:gy_�_����
�4ʸ��ͨ��}��A5ٍ",���b��x�R��N����OT�)hx2o��Ӊ�<�?��𛳼��%��L�����!�kG ���5G��O������#����>z��P��UOl�څv�%{d����Ǿ�2��I7��:�O���u[�"�K%T�ѐԖ_���1��[|�$���$%w�C��Ƅ���mN��ΚG	0(+���)�,��q��1t���t�+C�������	t���Ĺ���<U|���%���K�����>Մ�9)���"/{�
촧d�����~��:K|Ն�Rk�O�Y�`��U��P.���=��\|��,c�dҎ��
��eTS�E#>
R+��kd,D8�������������pMx���L��3	N��KS
f}���/|w�x�[E�&�����+'�۵�[�V�^#��A���Ry�P��bOntX:B"�|4�ri����	0�|���_�6�ƍ@�!M x��tYR6�W��\���Y�]Jֲ3�Z������H/ە3k�`�C�t{uᙧ�[@}�bkJ�8�����f�TꜴ�*�	W�$
�1,�`�_Z¥�M�bS���0�a�O@mGmf���ש8L@vn����Cq��)!Y��Q"C�q��_t��P�u
S8�Z�ojYw�|i947�i&ow�l�Is��5케���@��� ���f{z�ھ��^W��-�秚��:SK�m�5��D+]����*	�L:�}��A�:�X
U�ێ��SݧE<�Q���Tg����OS^�da���!�9�[�L�s��th�5O5�MM7,t�QR�T�][Ja�X��o|Fį?�8�Gɼ�<f��g�����_�FV	X"F���;b�S�hT��g�f��,��ى�t�;G�ID�su�Sr8�x@*Q��⬷@D�.�nxB��*vs�� �5��G�>C��7�A�Å�q�����O����0P|�X�=əK�ꧻ_�E�Cd��?M(��'�b~ر��7��vWG��\3]�~���u�4誶�e2NB�y�DG��M�@\?
sjŲ�Qz��䭆��{{�t2jJ��s�ݨ���<`���G�\r�^�ng��:�ほr6��w��")��J�U��̓>Ƕ�'�ԩD$Qq�wTw���h���A��y� ��g���O.@W�*;���]����4ɥ��8�!{_����E�B��O���jv���"��y�.P9q{K��P�d�L	�$W7����^K�@��U��3Ҧ�0�E���i��ف�$���D�J�j����ʜ}�A��O�{��	��F�K�s��Z�$7Ӣ~c6`��(�-1�_J�u��W�rm��0��l�����_ΙG?)Ab�n�TnSi�r���a�%�g�E�鵊.�ۥi�����#=}l�(�*v<f���z�Bw~l�������
'���|�����t�'�U�z���`v����Xw���u8�@A��K��*;Q�E	�6��CNZI�U��]��J�՛Q�1WJ~�D�w�dU�V��u�s��)�����(��g�X��7�ȣ���r��ޏw��;8��`�ή6�7ۣ&1xX���+�hfV`��<���_�,?`3X<��_��P���,(�*���*�53�p�4���#|�)���y?�Ǎ�2[�s�]Iّ�ˌv�a@�n∟2$���w�:�%0���������eT���6ި����+d�ǌ�q֗D�.O�>`�nW�nw���׫z���B��8ƛ���(�K��������6��� ��(�7d�x4��3�5Ưe��Is�]	��Rn쩍�ZQ���m�6�}d��Y��?��TQ�M��;s���=O͉b��]�Y���́i3~y��Q���c���Ѱpmh��4��u3eY{*]2��2>9�X����@�Rό�3w�:�*=������کa�<�����Q�d������0K�m�J�z"<�Kr�}mVW'�����i���&M��_i@-":��"25���� ^��|���6�kY�L^�V��j�Ƴ��k���k�����Y�s�V�8Q<6��DDK�C� ��H�yy�� J���0z����ӕx�"x<������F����H�+^-ӡ��_��.n\��J� ��`�g"2����)��9�2L{�¢:��c_iɕ����ߗ�WPJ�x�F�/����R�j4�y��V��U�r�����_+5;��D =}�����n�Z؁o��l�Y8���$m|8�E�&��J����Ԉe]u����;N��W%y�J����fm�����	P��A���:s��-�P_�ǁ<ٻ���BV����BbZ�����t��p:�'�l�V��4c Ζj&x��������2P� z|��V�2S���Ơ�Y2�0آ��Y{;B1�;  ��_zn\J W��'No������M]]�1�G=�㸟u�Z݅ ��4E�RF��/ӭw}������A�X�ii�����������lU:,���(%nX�Sœ�3����K��Ǘ�V��7�����g���u��*E��Ul�Gr���̧d��<���D޴�"�����+ϳ��D�*b$\�;�_C��A���ɈwW�P˨���\��c�'����іӶ/������V����`O��J�B�V��������Ռշ�����cR���s�d�]mʃ,'����=婅"'�m;7i�;0RY���VW��-~��i�ftƛ]����9�ri��ބ����Z��6U��u->E��6"�"�K��xfa�[f\vA*��WT�q�"�}ƶ�����	�S}H+�"^t���
��~Ŧ��.V�-̛��U�d��j�PN�A�I�����
p�j���&�Y�`��Δ9�B{�4�2�R�ǧ��G&[���������A(�xZzQ���Ⱦ�|Y�����ۓtK�ǜ7��.��'�7l0:6xN�B�i=���WG��'����/wO�?�lY �<�����d��8����^k��Zd�,���[)D��+�vϧ��}��Gh��ŔY��,5���La�y���	n%k��
�~��!B@1�L>��p����w���-��'�������Ԩ/.{ ��q���|Qi�E����5@{Gi�&c�+�V�,?�� �פ7g2�)�I��az/�=���s�<��'cR��ʜ_�������w�w呸:�³�@�^4��V�xJ~���ޮ�6��d�q��ߙ�c!?%6���+|����b x�b��|������ď�~��o�G,/�|۫�6�ު>mu��N{b`���X�a�p�@��]z&�Y�A�L·SI�8G���1'��U]���jA�b�Y/~Q�,A�U�z�%�'�-��4������Þ����Y��bJ�o�6FA�S�5�wR��kCG|�9������C��3���HE�1y�,^�g�\��~��)6�^?��s��&O1(��F��Cf�
�ՙ��	n#Xk��]���H��[:�d�H� �Ԋ;��`Τ�M/��z���%�9)NY��[Ta6�W�譵,��,2���hPAe�9܌�Ñ�̘UW�x<���u��D슭1���B�	m�I$[�-TPJ�+�z��u�)d�)Iry-��
�a��|�,Ⱥ�W$qèJ��6��>|%�ĠɂށJ��&�ՙ%M��.���=����Wos%J���,?���ׯR�S��������o�9�9������R��yW0��4��r`jC��\������*Y}��܁���_�R���ηґ$=�\���T��mSȺ5�V .Uߝ��Nܨk�,�&s��8��A��ݞl��ĜZ_|bd$Bʵ��v��f��R��W?iW�VR�&�)�l.���gڗ](�/E�z�f���-$"N��)��`�s<5l\�T��	��o��,�gxh�$�%O�c��q~��c��Z_�p�١���ϡ�2��e�Ab��^7�p��W�6�^��]g�������ㄆ����~�?BwAr)���PK���FR�@o->�Q�Wݽq����{x�n��D��%	1{I0Y�K�-Vڟ� ��	��
�(r�Ub^�E�p�l,SK���fgk�Oe�i� kRP�l�H��u��� �\<�s��rU��N}x�&:v�������
���빏ˣ�G^�y)$�-�\�tΈ*��c�u�����d~zN�7��m��{ʡ7� N�N�=��i���\��?���{���E�L �x-5�*
(f���\���-�1Иx`��4턁� <������	H�S���.��Q�f���6�-���R^��=�?�3�T���<���r�KX�/��ٿx�[�:2Ge�[Q��nw��D-sA���d'��4����� �ZC��T����a�X�1��]��؛d����\�f�B�Y��4�	�+f�Wy�����7�v#"� ������ ����`�"��J(���乏��o	أt����>Bv���
%H�%q*��$�4z�nΧ�B+M=|jd�5�({�����|�o�MR�H�	�K����-��ܚ߈r���r_+y�t|������^�Ϝj8.Q_��#��!JQۏH��bc�_pD%�c�8͵��X�N���2]ia�mݼ����J���S�1<�y�kA�A��,JϏ痷2m����D����c_R豉l[���b7k�z��} SdT�.  ?�X5�K�F�<m����we����5�����r������?���cy�]͐�]gQ��M�L!�5��H��,1pD�~��y�ࣿu�w-�㎋��.�q}����A~���H�����Р-����w	�M�M`�<�ġ���^v��n�pDA�ݱ��)Y+ª@��	3۟�u��}�*V2�j��Ҿ����*�{hb����nJ��1!>��Y_G$�������m�s�;��N��V���<���rClè��"�3���]��%7�-�&�j�Ï�~�<G�����~��L����1η��uV�n�����} �= ����ԨW�i����N`��6�A�n�S ���}��}���D$s���'���Yn����������:�K�X���@ ��S���
H�*�"�5�r=�[�U"`�u҃�Sp����Dm߮|�x����]��\�ܪ�:�I��~��ѯ��p��@M@z�Նʈ�Rn0A�@��}�� ���k���t+�h�������)�Շx��rֺx�Mqo@�mMh��g�*{�C
&�w��Pe}�����%" Y$Ɉ�1޵솲�$C��sS����a"���e�XYQY�)�����^�H�!�Z��I�l@����M�O@$��,�5(m�yP�4>NuO1%q@+KR@N�1W���$�3�):62����J�$�O�ǕK����:D��Fx5D����T�+e��!' �+���yU�ok�nطpU�7��K���j�9�߇�a�
sµ�et��6܀ȼo5��1���Z�C_���'�c�ހ�uw�q�c?L�Nm�D���I{)����-�ΖS��c��N��Y�o�Zu�9������k�Q����.�	�~�(dGH$T|�j��R��z�<�6����A��0��^N�U�-�}Ij(��&�9\|�=R��ΞBX"�j��EF �{8u�΅&�~�3;�%ܚt�x�Rf�/&�ھ��q���1��?r5_��ڭ��D��������<C��d�c�	Vh
�g��LR68��̬���~�:��^����r�������Ys#��j�8�I!�m���U.����v����t�����Cٞ �BAۨ�I^K������?���h�ʀ���Y0� ����#v�q}u��/��s���T0b�O��7w�޳��++�����/a��oD;Wn��.�Le�i[� �S��%:�Id�����Z�c$\	�P�����ep�9�Hc/J���](PA�]؅�R��"c]���ƃ�t_X��%����nP����V�Ȩ#�����E���l�x��\}�ڒ�Dù���2�ݖ�N�B���_�W{�.C���Ϩ޽�Y7�Ǣ3�-"g�8��j�̵i����swV���l�l�gk�%����]Xq�'��0���!k�p��rW]��B#�E�#�KR�Y8n��m]�[p}�7�xw�x�<���C_�<��y:	+9�T_#�C)����I5R���\CL�v,Ń[=�ǳi�u>��I�@W�W�ԟ#K�e�;,��\۝�q"����Ҽ1)�Y`�����mk�V�d��d	HpՓko*�j�9�`���s�=
�R�U
m��d���RO��@eI�i�� ��D���0!��P����O�Jy���-�G��g����u�M��m�n6�=ls�?��������ڵ=s�#Z񁇄��lZ�,��ʙ@u,�1
I��\�I6+Vj����dp,\�4�o�q��:�81�G��:Hnf��$�#
�M�C��(�CT߃�����ݖ'�9�	hgc�W����_xVe�'���-m9�Зl s;��md#��U΂��9;�8N9L��bZ�R�4�%m|f���P��>�K}��.�HW��8�yq~/�X�fIs����SyŊ��K���5Vt;�|I�۲4T.?��^��W���>^8�2�)*�^].�F��� �X��,�T��y�����}	�[����<�K�T�R΃�a���x�O�ʈI'piV�Ql��Ԥ�z��Q�3Hwh	{���
��c��������V*���D1��l�����t�y������B
G�G�F���K��]I�{��1�G:Vk�֋ �UVq>rR	d��NN֮j/�>Cl�ö(墝��C�j�.���O���R�J�^V��%�bvW��˭JH��݌�)U��=/m~��C�\���^q�K��]�4� ��<G���і�gt`����Q0Ux7����h_4�*��W9r���`h��mcml��j�0!�|A�)WzdZ<B>�k�I�\M�q�	�G�UHyڥ٢��[��#b���Ɗ�����I�{c؇�kT��S�o\d��
-���N���Ԭٙ������l�c4юŵb=�iN��hu@
t2Č��=cMrQ��Zɨ���'K爯��1��5��ɔ�?^hk�i�4�wY����I��w�s�-�u�r�?A(��9.h���?�j_Qg J��D�SZ�C���"*&��Z1L� ШkMJ2��(B�Lp-c�[9����6�����-���О��U��i�,�޹I�<*F�@�l+�_1X�҉�ߞ�+�� D�4�ʐ�����f�]��=^d�k2�W ��h����/�X�a��ff��*MQa+�����X#84͒W��y�i�TY�@��)@_��JF��7>����1�t�-^�Z�؍�"��+�)��ssp0��.���ąMX���Ӣ���3B/�,�4ԝ=󉚲������J N�g� �6�h��{S�T��k -�r={�G뷳ݩD���=�Q{�SgLo��l^c��'݆CB��$�#�=!� ��A#���X��<=v/���X=�S�2 W���sZ./�؞��dG1=l�au�AZ)r'����紺��p��[�AK��$Ni�5QH��v� ?�W.b�@ZT^n���N �+���w� ��,y�f�ٌ1S?�ȭ�M���&Dٍ��W�%g	�������~_6RL1���`lV�>&ԙ��x�z2BWx|��.R.s��	V��v� 8P���э!H1r�S��{�/����JL��]o I���i�'�=LE����X ��T2/��N�AO�p��n���c��2T\:��J�D��C������ �v�&E*yU.''��QJ��_�Y�9Cڊ>k�����՛<i^�V���jq��OE��/3CC��h�ʼ"���Aɘh�4�H�_�z-Uc$����"]�,5a�J�l''<��Lr�;u�b�݂��|A��?6��������H�7�u��i*��'�~<��*��$|�6�єi��oZm9GsD;��p_۷E��wP??f�3X��f�g#��J=�ި�{��h�h�U���!+�+�^����C��=��$���^HI�Cԥ,=kܱ��z�ynG��-ƪ��~��ױވ[�I��k�UW{8W�W�L�m���=�2�����|�2s�Q�X�K�|@���O)��@g3qsI:��$�c�](� Ln]F�/�FI	>ȋ'4W��N�~R�Ƅ����{�EU�k�W�ާ�Z�G����"���?��M$(�n�0T.o����Y�{Rᚨ'��P�s��Q��p,�|�)b0�����b�h�./��}5�xM�ab���$��DZ�WJl�X_�����Vj�}%t��L��@7Ͽ}��������yb�Z�Z3t�*;	M0��
)z���:�,���sLYD����o@�G��	=Bt}�Pj!XK�I�}̄�L�|��Nc�ϘM�|����[��ܭ�*�PEߌ��e0��5p񀛏���)9P�s <�2��#6 G��sn�X�;[�>Kh�//�Ħ�̥Z��-��-%�,T䘶 Y���ן%�x�0EHa<�i�%�G�*<iDQ��dI�4,����Dz��鎚�?ܜ�a�i9��K��7K�����"����\�&�/�j�e,)1���ɛo��ߡ��b')�{�Qi���Ĕ�oY�d,. �
�#�p���ނ�w���I�Q9�Gj{Z��Z��{���w��Ή�=����d?�?�ZM`�r���:���;S+0TA/�����I�w]I�fF���j��	�tB�]�|��1�]��G�N�;L���8ҏ�8�q�P����HG�y���>��ZA�۟�"a�!���W��?�rV�����٬щ��0����λ��Z���'���z�(���e8�۩B������<�#����U+0[���n�z��m�K�:�w�N��#��3�;�Q�����>p݅�콍��@�(�W3H�KH�o�?\a��T�~w�2BLׁ�	��c҂zf�;����*��=�L�t[jX��G3�b��}F���.���C��"��a*�Uy�r�' G��#�q���vS��M��8�(�}A�Yz�h������_���ԈD�'l����L�u����]"���+�>�f&[��(\{��՚�"��\�ru9u3i�g��MQ{���k���ŒD�
u�G7�OI'�ؚ�ũ�[9A�N�4v�QV?g!���֬k*|<�l�}*�����P��NR��2��b㯞s���ҡ��F�`p��i\���/~Nç�X�af�k�]@�kY��a[�U�s�ƺ���9��<2h%�e�D;�
�ZW�GKk�X ��x��N�i�ȕ4q��lJ͔�ϯA;�޽n���c�Jp����M��jMh�sK����ֽ�	[��4 R
�=SN�"$���Z��(ӄ3�hw�� ��U�������:/۬����#����aS�];`����C-0��L�R,��^�L� a��._
!�k�d��	wG'N���P��.�����Gv��6^*��V["NV�9�
�K|�s�Pj{Y��v�@O���[/�D���N.�-�%���7�5�P���ru���4G���=a�s�z�_�>��4�x�'���Ʒ���&T�ʋg{��Y�~~��tv�k>@�p�6I�MRRy�kp%Yxh	�����M^!��wnbv�OJW�M�}f�(�=W���I�tO)vh�}���/��=��Jp޽�h��\sR�8��q�����Z���-���s����gY��7���R0�:�k� `��2�`Į7W]Y�̜D&`�H��v� ���>\�Ӑ{�*B��`l[�<J\�b=�`���M�L�%o��fF�DJ���z~a�+�wp	��{w���D��+�o��p�e�������(����,Sn{_+s�}��SBHZ5;)��C��B�@z���I�Nb`v��g ������_�
�[�1�Ib�[�#�����W{7�Y���Z��8CL7���sz��$�vMN�"��J��#�Yf�ė^XN��,��F|׵}Kc��/�mT���/�k�!4� �фs��g��~�Ö�K'Aj������ؘ&�����G�[#K@۠�H���S����vħ� ���(
�@��dWK���j�X���u'g�ͬ�ǁ�Yd���"�N��WVP����M���IM١ۍrv�\�k@h�9GKA�W�(���N�9�4i��`�H� >�Is�����,+�@�g�W���)��7^���x�Q��`��R�
GQM�i��-��:'����P?l��k̳�R�D�Cw�7�H|y��I��Uid�/���Uǐ�4�Hpױuvw�I��Ai��z?���ō��j�UkK��>s�CU�yYG����g�"^0��CVG�K��VC���_�э$������?�*�3�R��m�r�U���W���6����e������<�`Ƃf����_[I��q'��(G5���{4�V�L���!'=Y��Y�bo�JY�1�����?�3��E̕��� g恳��_c�:�nU�v3��p��k��o�ݡ����Q�^���|߅�Sܶ�|y�á鋜e)��]��u��H|�i��-����_�I���F
��x�ק�;'���i�F�[DG�J�n���^�vh���Aڳhd����=������㐚%��r�����qj��w�>�s6��ǓF����r��uX�Dc���PRvn-����qA#�{�b��k2�47��m����3�
�`hԜ'�a�-�S��}/�M�����ja\d��+8�f[�;N�tɆ\f�ޞx�I��\Ш}��1zuX ��*�R�"-H<��)P&+a�2{5�M=���҆Ǯ���H�rZ�����Ä,|�{���֔e�5��5�\����k����ƣ�buxG+$�W�#�km�k���T8�	/O����,��Xv���2T.h8�'j�U�g��\����d�H"��L��H�#,vXY���KE�Q�$j����8��;�#��N��5��:�c���.{��W{��!��LM�c.޾�@��w�*(��(j٣�m��;�F��-�K,����SZ:���&��� ��#1��ۉ��[��T�b����	�cEu���#9�6��m���'�m=t���� �80}0á@_;��g 6���P]{� }E���^��X��,�0��vЉ�9�8���?\)=�s5�I��|�o�-9�	����)52P�Z ��ٸZ}Ջ@�1�&��@��J����@�.;
=���m�.'�DW�>��\�h���`���;�E8^x��a���,(�#8�	�����n8Q���<�K�d��<�x�(��n<£���9��R�~6��}��������j�'�쀼����^,��i���&�2"�s��H��o�-��n�����+�K3�N=sX��P�k[d,X9+3�w�������S���B��u��[M5+>�yF�����Fyo���4���j
έ����>�AO�
(�i���8D���O������S��%�\-�yx��i�8V�.�D����aK+�x��MJ�]���b�>�R�5ޛ�=��c�mr_��|X�Q�Ofo��-�Ȱ�jv�Fu����vN�G��w���f�8�h0�N�Las|N	qE���X�P_%�Ԍ�1�ˀ65?�"�.�ޙ����6��8-�4 �����,�.�r;_�{��	�~#=�A������}�#��U*|�ۿ{@�:�Δ�M�h�(1����4�i��]����!���O�ؼ8��O�x���>���Q�DL����>���r��"����P�4'3n�TV�	�$���jb�"�i��+5��D~l?ɋ�~]	$QqZ!�Ø:��Lx4�kA���r�I��L��Y�2Q���Ϧ���'�~�/�vBh*�^����dl���o|�g����]@yx�c���<�\�z��uiOQ���5���*/qp�#�QZ
��\aip�;�+��,Z�c!����o㏗=K����Ÿ�RÇS%\e�(XgT�D�w��t�C7
dKzҡv��#��
[:�~��N`֍�n-�4�泒��_��K�M��MC�%s(^��,Z��}���y�(��<q#����Sn�={�~�X8�d�l4��#��ĆL �����@w��5��ڐ0(��bW_�� ��#��������Y�T��E���A�}�%���_���I]��H�{yG���1a;e0���>G*�4ڹ���!��fo�BWl]b��h���]3�3C��%K���3$�L�ƍ�y��>����~�z��\[J2
�$��DR���)���prX��1QT��F��N_�`��u����S�'ƛ��Ÿ�'z���/��-�y����Pt�F�n�H����0�志{���\i=���FTk%�����h/h����ߤ85��KI/�&�g0�N���wnyV���K L�Y�5�>\p��
x�հ��s �:x� ��1��O(�A��z��Z]B<�>�@�G�	�C�]��OҘ{X?Z��s5e{�L�w�0�hu.~��&T�-2���E��x�[z�H���s���־��] E�,�G������~�e��?�~�{�8y0�e�5���%]��Թ�CىFw�׌�m͘/}�a�'�ZԢ���
�A.#S�i^�A��$n�QN�z�m�z�!�E��6��͏�z܍�
�E��G.>��ɕ����SaO*�����Q��2�Ǽ���w\��_q�L��xoS�3����}o�P�����Ԕ�� ��d�����gϭ�NԠ������K�L��<p���]���fWnS�$�J i+"g�7:ؠ}�܃-�.<�*bo�cy�O`n���h��v��,B��l/T�t�����*$�+t3(���K�,���pմ*�fjW2��G5k̸��ȉX�}��T3�w꫿%!������.3��\Gr����JE8>{�;Sf�I~Ut�����)i�����-�3�Z6+gg��jB��`���X|��-F��ș��Aǌ�B�K����m'�v��?h���7b�R�����wܛ��*j�'�2�P.y��yh���g~���j�t�}�W��m;�ʻ�q�q�3��|���u9:FF\L���� �_�>P����Z� Po?����N�2��;u���`���0�w���ֿM��?��p�X6�I��b�pK�S�`�mU�ou��c�(t���o		*����(E�ⷥ���c}�HM�0e��k���m'���)��i�C�DnVe��󇰞��������#5R�Z����`��T�avz="qϒ/���@����ħ���Ǵ�I.��B8�t�8�ÆSph�M���	�[3�БN���'6*� %%+��@W�o����*�O0�#F��_�f�Yyi<с���t{Nk��s���UE�a�l_��Y[�.�v�ߎf�{~�!��p&��|�	-�m�9/���m�c(���g�q�.�~�o�,���ɉm��JK��+F�Q>@��*;�}]ӅK���	
V���Ɯ	��F����>�,{1s���d���ٻ����c��1���O׏@q0�`���]A$^K�-*�ty-��%�`+1Bjχs�\ ��IC:ӛy�����?�&���`g�R���zZ�D�k�4������I�A�� ���~"��䭍�[���g�����q�!�=��9��vz��L�ߋ�p�{��p�ǉ�~����Ɍm��5B�XVP�/�ʡ�/J*>O��\eu\���[�|��(z���X�Ӎ�Գ@$������vq�cx�?��~���k>�>���\�\�x�]�U���BAeDG�WB��
�/��>b����� X��h����<y���������X	��f�A;�L\6��)����Hr?��=BOI�WV���޽��."�h&Y�����[&"Ǟ�E�^X���/ҙi�������}�m� ]�2��=�"����H-L6���u��yr�xPJo�M~c�u'�S��"^��j	8��M�a��m��	`�^�0f�h#����i�@�-��e�=z��ݒ����0}�ըM��l$~�S�L֤��<$,YA��Nr�R-���� @�LQ�e"A*����]1K���f��۽�p��m9Su�	壎�"SB���m�	�^#F�SwPm�����[� ��'׽�~V{*g�$)�#����ʊa�����C��+Z��
!��Ȧ��OEF}&�-����ԏ^���Ga����Ť���P��gi�-����>��&�<����~�(jA��*ǜ���q�$��Қ��}��,�4�e|���^v��� Q��3���7����=����Eӽ�-��n�Z�6Jg�ޜ�,�b�qۻ&� �����	X���j�~8{%o������)\��Ǿ�m�n���V5�XA�t%/�B����7!���W}��C�=�2X��e�]� Eb�
T������}u{h^�Qyp�B\Q��D8i�]�C�h%�5˒Ϥ�х�&���&���e���4�~��~�+�ءm�csg
f�G�#Χ<��m+�t�|
�����%j^7`t\&R!LsF��To}k�k8�9��q�U0}�gI��-yɟy�R����Y��z��j�HJ���nX�@�l���Y�w�ic�Qac��2M,���s/��b~M@�>�Ę��qL.���S��|��(uλ���F�'��n=ii�<�<w]�H$��~zgY-c��$٥��4���F��6*��"E��_�ڀ>64���j�l�z�y���-B��x�/ߘqh12�#V��J�}v�8Z����D��PnV>���vZG_���T�˯"�j8d�
�O����ը1@��_���\�6o��ٸOPo'�#�_�ߖ ��J��\�(��������6�?K�W�0�4y��R<1�<���1�'��X����[����8�2���_6����e�l��X��� >�}
n���C��Tr�X��Z�rЙ���%��ƽ���5��A�if��WF����>ť(�����}s퉗S�<{uR����C�3�����;�������s��f��}����"f�A�������������æ����
�	�7P(�'T�z�����ɟb��Ҟm�A{���#�>���w��ķ[�^���g���H�}��6m�+$����	�m�2ʐ�0-�Z��sCGT�eOb�.���Śn�
��꜋'������t�h,��A����4��G�S�"
%�狆kؚZ��̭���k��z��'� ��e>DA��cV��?L<3^�j7�֯hH��K�.Y�zk���KH_D�N �<dMښ�(;��1t4�������6���.�}��l���)V�i�d>�l�����4
r6�Y��:�bEOe�?�����TJ��N\I����5H`�"զK�L�@��I�T�����K�����F@⡾<2�᫩ �a/�j��d*�gi߬ԧu�T�YDb
���'N/��YL�ܙ�ȹѿ������X�s��-��:�^jJt����g��������"� :�)�0@j�Wq:�zp��7��SfRC�����òNI}!���j̓/C˥�Dr�������3"��Tٓ��Fæ�RzOs�9�
Ƚ0��0�h����R�9�_M	��n���q\^5��KN%(;�n���cɽl�7&g�K |������^:Z���(V W��.8y����Vb�k�j�t���a1�.y|Z�컏�À&G8��m�œ��+��Y����H#���
����E�ˣT�ê��ͺ8���A�c�����-�A��*_X�;�9���3���v�����s�Ǌ�R�4�/z�%>9oiw{1��f������qP��0T�Y�ł���U��f��dL)�o�oy��;�MW\���,hS6��~|n����K\Vξ� �p�Y0R<�o��hFi�b��
�]k��n�U�e�l6�V�[N��J}��2a�ρ���/���b������A��sd���k=�+��+Ɔ2N��^�`��z�f�R��S�TO:���������#����I��3�� j�S���i�^����\�Eʞ1�Τ�\ʹv�l2²��#�r�遅�Ȋ�g�ե�"��D��{P���� ���.T�A����-�3�d�sf�e�����j"�Y�b���c����i�r�1E���

:�(�]}�b�r�n��Ĩ�*e_aLT�!ٓv�Yeo�uh숈)d���4_n�jq�"@���؞�?
W.(��cμw�5T2u�p�*���H��6$v-Џe�ʈ?g�_~���1[F���2��pw�_)�]����{�݂�Uk���C�b���)}Ҭ��j�Os^�ed5�`glN��Dp��u �h�޻���=1j"�&�~�A_d.��ٛ94�Z4���!#������sH���-FQ�."f+}���S�4�B��4�R����w�m!�mIlQ�~�-��N)����B������uB(�\U�8��B��%Q�C�r��nJ�?yo�f�d"�-�W��(�j����A�e� )@t�pnB�U%��<�������.fLܠi���o
"��1s�ڔ�s��0ѵ���*�}�pSp�ԝ�sn�+�ʭ�ݵ������Z��A��D�W�1�N�f��m�A�ɼŻ,��{k�Ym7�J�
s:|Sz��������^JB��-T�.�Da"Y�B�o|+��r���+�G�+T@�s���.|���F DSM�֑����|�V����Oh5��&���,S���U^�)c�n��y�)�����X�v��1.��V�}��i��t]�:��xo�4����W�iO�9��=s�׫vhny��c&ue��&�\�;����gB$҆ƽ���2����|����`��(��?k`ޖj�`71���|�8&k�j�͟��^F�GB�PeQL8ɽ�@����5�>ׅPVM�c��c��҃�B��:||���T��Sd��M�S��-B�2�V���R��#�m�g�R�2F0�t����G�r������}���EK�x���O�7����+�E�^٣��$��Xdh1�|l�&����
�+nA]%IG�?/�#6b�|�q+4�Hᡬ�o��u�J>��%)�g�!��3qy�{��*g����"Ƈܜ�y����s='$)��`��aW(��o������߿s��"�LGA��po9���T��H��\8��u��2i�ЕxE���F*C%ׄ)���o������[���8�������z�D`%6W^�@�g�Z��v.�����<�����&�{�G�-�]���|0.�-�^��ΜK
r�س�V�/�N�+��^lA�'�NdT�0�G��H|u ��7z��뼝��)�>����3�7@�}5���^W��q�"�Ax�i6�1�����7�Q���5T�qt%�ͣN-�V�x��޿�^�;�{o��)(�y����oAt�p�b*p���~WXq���Pk0:|rc<��Ї�҅uz����/�Sf_:�|�oa4l'������ȇ`�dQ�N����h��8�Ga�t4�A��$	��)�]�,��)�U�ƌ�N��6 ؈��uX�Eg�L9�U%����	���0`*��=� ���`\p΢g<Q>T�lws9�]ش�P9r�L�j�~�^T�Yh
���b��	�]z�B^w�x����x�.K� ��x%�N���m�f�����}l-?W�V.�`���w�uh޳���~����~���XN��݉1<a��yp^;��,!�!��t��1�*�W���Mu��߰&ӟ�����y����i�(�6�׋�f��2Ef&���m���!y���PX�ͭ�3�Z��U+j���m����t_-���v�c��d��<�vX���U8��Q���ʉ�UKA��Am���d�g�(��������^q`C�^� �+��:�|�s��c5:�2�c�k�c�E��`ꑉ\;�A���J��TI ��+IZ��4���={���tF�K`�YR�3�Lܰ�wͮr_�T*M:`�Z�q2S�0@<��?�@{ ���� �'rs�� .��f�$%$���%�y^UV��=�|<��c@ v
����{�x�v�r`���_m���A���`��!��4%&S��!�`�@�Z�[�U�����*�9:�'�ROv#�S�ZA1I�PƗ\@�ؙSM:��V�G 8���W�P��n�CL}8y�/�z�q*䉯��M:�<�y����~5�	�8N����=��BL�`�s:��\�����4Y|s�ڊ����e�7fy��hSl(����)��C��ڣ�B!1�5�>�Q�֮��D�g���G�k�P�tqWނ��.ol��nZ$��
�#�.H|PXo��d�]�WMZ��r��w\�Aѽ��O�pL��9��T�>Ig���~Z����/�Γ����o�$���g�#L��=h���Y�^9
�VAJG;�w���6O��¬���4�@+
�HŠ��n��%�#�^bٿެ�fa��k���r�^Դ�	�æn���j.����O�� ��.��B�	\O�1����E�f;|I|��B�?9��P��� 3��p�(2��D�j�|:T�m4=��|�O���(F�DtM2�
�1�<�����u��K	dt,�D!�HS���3y��)�`�I�ȕ��󕖜}�	U�;| ;�ݥB3#Ņg��K�54,�l���%�=��Oũv���ke�/Fj��j�*���� �J�b��ڳ�YlJ��,�[ȣ�����V���E���5l���~(����J"�������͇�%@"�� ��}s�jeJ-9ꨉ�x��i�����-&�7�8��c��(���C!"L�&FQ/9���������W���h�y�*BJ<���u�c��ro�n*�Kv�u�A�vMӠ��($͆��F t�'�/fAS,=�M3ԯgQ����Hs�����a֛�|,I�@.)G9oX��گɆ1���藎���E��@��:}_����r�`.� X�$~�)�y�wm�7Jp�[�+�P�Yr z?/.p�|Ur7!V��/O���|�k�7ޙ#bG*��@V�*�[�Q������sk/zs�Wm~�w}��� �� G	[�Ķ���t<���|����)�o8�EN>���DanH�s�Z�M������M�`�������O��o��9r�����pu�qyM��)�9;F���,J�	�����8��Ǎ�٥�͚UD�~��S%��*3#_`�As��D%N[�n���8�B�_9aݙF����� '�+����VU�9nBM>��xƸF�oPﺣ��$�b��M��L�8� �Gj���oS�=z����(Z���s'�]�k9ju�s����S[Vu���;H��i�l���,�j�r,,An�����Xw���
�D�0��"֋�6��Ց���EGO۝��vH�ձ̭����3�W�W�^�A��'Sn���� 7p ^�I�^��pZż�3c
��0����O��D}��
@p�l�ʎ�T�OsD��� �D+��V%�pI� ��%��K7m�x���=)>������~Gؑ�]�HL�:j�f�&��߸�c�i��o{�1QPnC+��L-%uFDZu�Ԩ����m�z+���\'�퐭�ǃޡ Ӗ��$[�Ht�w�Ă����_y�0�M�D����nk�4캪>���5���\N�F�3�"�4��J`�GxS,�J�Z�v���W�qG��6_��)���'qP �D�%��70F}N�tl��}��V"u�p00�7���/���87!��	�L5��N�@��yjqPr>��)6L�H_���^Gݴ�d��AbI�P	Iǆ O4˗���g-�yfxC]�N����\g�6=.~���r�A����$T�ǡv:��V+��-����*�ٗ:����+=4����L3�I��OiX���3X�	�2�{������} ����$//~A��C�/�_4���!�}��+�����.˖\���-�;K� X'�@�6Zz��8&h�TX��Roco!J�I�	h������~�.��|bt�n�p�e/�[]S�z�y�%&e���C�����'Pz��iPx�eԯ�W���/��,�?�j)|ϓ��S��ˣ	tRN��1�Ks㋭��N5'Z��������#�C�2� @�dK�i�=��8[�IE#�,*M��MLv\��Ja�����ę�?;.���¾��)
�S����j��Ѣ���ެMU����j��W�x�ꭼ��W��/\چ_�O2u�I�N����	u����~)m�U��<�ǟ�~<dZ���F!Kk���`��.y�=`��m{�k�Y��|Tmj��"��[��^�<�46n1��/��u��t��I���)d[�I~&x����do9��<�x3J�Lv�>�j"�>����yU���u7W�ig�{?;�*�Pͼ�9Tw@���R��.xK�t��?�� �c��O�i�qq�/���Kv0B��ju�o�nZA����)��Y��B�8�	�!/+'${�B6��z_��-h�N���O�bF|���}��,~T+��r�Q���=	ދ��&�V�i��2�GE���r�<�IASb����n�F˞�_N��%�ǆ�]���Ze�9W�" ��m?�	�����"�����^K�hs�3B,*]����K����.��oO�\���Ȯ�ԏ�����"b�PCM��6��	�)��;��ɋ%pcZ���X�H�����r�{l��z{�dI���nA��D׮�T��dL:*ʐ��v����t3�O���$0Q v�*�oU��wk�Vk�У� ᮀF��:��J:�󵑵s�p��L�L1�Du�C�����GS���F��uw���Mf�tĺ�$2����:b"�~Î4�5Q��r���K}QF���`�B�Y�V�����n�Tr�F|����MF�xd��^u��_�zt'��K6Oy:�F������� ��|��a3.���c�o�PN���#�*�+l;�i�]�����`|
��閉����&\�Ǚ�y%�u�6��Ng���"�.� �~X�N���B�����Y݄�	'h��f+�BE�"��l.�a�>y�J.��`�7�8�i
�"J:�ʩ͂�(B;�H$z%�S�L��(�4����h�<���w}h���4~:k�P��WR��Э������l9�d��lu�(��9���dO/Z�M]���X�ev0;�+��7������������������y5���]y�7G��[�ÏW��ϳ��!8j�Q���3�@'���	x#��qS���9�c�ؔ�e���j�u!\W��[w�\�|p�v�����kvX~A�o�7��?��7������{Q���v�٣(u/�!8j���?mє�eZ���/�{��?����{A`�Q�:l���E������c^�z�ۚp=�?�K��;G4���Rr��=�8�1�I�H7���܇�Ճ/�?��}0ކx܄UNK�����F�@8�5q: =�����GR7�ϣ.����1^:���A-#���_��S%s�C�H��7%�1u��m���_�ڻ���|�IȺWKRFiR�͝��h��z�_�U�@�y���g�XU�d�ÛɎ�	�#�*�h؁{Ҳ>�1%�p�>�h�2M뾶�z�#/�NaoO���i��g�6*K?��Zi�e۳R�E>#����NB�π��U�L^�4�a�^��?�)#t�[%�?��N+2�@����7q������N2a��g&�!_��V��k�vTׇ�@ظ#�����w�e�X��N���
��J��ߏ{����#�3�2�**Q�Ο��9�q}�AONКź����:���e��x7�qJ���K��x?��3�H�gk)#rX,_w���#o�9���7'�8OT� ��^����^�T ����w�Q?��qñ�Bl�l]�1$JM�@d�e~u�K"�������T��P;Kp��!�F�o��$�u�`���!>ac󗜾נ2�A����p$��w��H��+ٱ���č��0{�4�}�M.#wg[�$@
+��D/�Iq��u�03�k}������Np�{�=�v���Ll����^O>_ڇ�2�*ځ}��+8cb��]#pbJ�d�50P���f�̺OOR֧�Z�)����Q�pC6�lC��x_(�Y���H�!��f�I*IBK���`D��?amOV��\��LE�o���/�w���
z�,��G�,u��0g��W���2XS�Sq�o���C�X5\���M'�ٴ��|�o�))�i��U����I�yƲV&��z6[�㘯�[P���1&}<��XpTs#�A���t�ݍ�l���鸿�� ZA�H�pQ�f)٠Jʂ����ܮ�#p/9��������ôrW�UxȮ9��f[�CkΠ'��l����#L�G�9��Q�׿Cх�[�+��5b#�I�)#�/���}3����&@����N��Lg�������²�.��x�ݏ���:�^*��@���t���w�ۑ���/��e?�[��ņg�����ϐ���C5��g�nu~V�gË/�ǭ�D]a��b?0�ϫ5�d���;ڣ�އ([��.1V�(��J�BP;Ź�]�-`(�8�B���I#�ђī��Ì�t��1i���䙒���
?]O�'�D�>YW��`#��+/�۶*�$^!w�r
�+n�rv�_bPt���I|�U�\R�3�.�?2�@�3����[3�����H�K��nZ�q��.��sTunC��bK�q���d��j�kȄ�=M�� �;����]�Y?B,���%�f�r%���-�y(�Fz��}���E܂� �J�z�2�I�Zs��f�E�T���̎�v �Ñ��q���6��mK�3�!�FK\�TԎ7�ܭ&P+�Q��0���:٢hŷ��B��?����g��v"�[B_�g0(�=��ɖ��� �%���#F1F/*�4�=P7������Á4c��.�:���ô$km��������A]ԶBE�ABU�e��9 ���v{uj ~�C���_�W��]�(-�Q�v��*Y�����U�pu���Ç�2�b��j]��k��1+��kT(��&U�&�>�n�*����s�b�,�ױ���K5��I��P�uA�[��O�Y���
W����aj�tn��[&��n ���u���GhK�X_p�2�x�"�}�髹)�A�^��.Q�-I,��9-c�
�ug���fI���Q�߈����-�����ebqV�Ђ+�M{%�s:f����
uм�c��
c����G�+��A�/۟?�e�fN>�i��8�_�"���7��f�g���V�!E1km��LG�W�&�ik�*�?��S���|U��5�~ٙ�;�+�j�u�d���)K�W.)��=?�_@=V����"x��*��o��e�F�t:�Ogc��g������
az���{�E1�T)J�~���R*C�o{��,.�c�P�[7Dʂ�����[��PWf��.�y0��'����6I���[�53��5�dP� ��O����%`Ƿ�m>�q'nC�f�1���M��y<�N�Nm��]�+]��[���тO{�z�e���y���Cp|+&�i��*�X1q�����wt����L-]� ���ؗ���"RÄ́h��N'ش?�s��r&8�`��t���2rߩ��WR_���hE�mx��O���ʅ"�Ify2�q�\'A�}�[�%�Gv�R�>=�Z�9� �`0b���T(dF)I���y��&���O��~�p�swD�~��yg��H�+^�φ�X��K�D�����l�Z�	P���+B����Ɋ��tk.�议�,�k�0�HB�|<{��v��]�ڟ=�N]]MB>ꈁF͋"F����c�8�z����2H�`����S�=ݟa^j6��d����,�pXZ��̖a�R��>�]���e��sخ�$#^H��@�E���Tً9��6������͆�k�$Az~���~!��%+�͟��qf%�Z*�I��C�h7-; �R�.&��.�[��/���~����e���0���࣭eF��r�FV�������U�e���G�j���%^��(�������&ٱ�<<�ʐߧ~t�/�:�ߩ�$��}��Ϲ�̀�}�t���p�W�"7�%G�^&��s�y&-���y�8�cU��G&$�`����M/�x[n�)r�/�_��m ���w\��'xA�^�Ȩ��XV�d$�=�>�\Ȭ��A�񰏊�4K�K��c2zLN
�"6�XA���t��N����8� ����c�����>��k��:Erkd��]�2JX�� �LC �BG$S5u�Ȭ�Ќ5�|��)��q�ٻ�W�X�R���V=0���b�4�ig��%���������r�� {�z{��
D:���]z��,������7�؎U�?H�'WgE�R�ɳ[z�%���1�z�)��'TbkbA d��HL�������7�훴�'8>|�|�}"ێ��8yx#��-j�l?R�4�֎/x��[J<�4tNU	-���T����,s�q�[0�,Yν�B��
Pò��Y�:�R���������i�V#���5�$����Ʒ�jq"+�Ѣl����W�[�ǹ<�Ϛh2U?�+d04u���.�y�Qt��T}�v�U×��Uo��2�ṉMT o���蝧z竤�r�wC�R*0)(���2t��!�ð�{�S����R�Ø�WșFWeEA�BiMP[����,Ϥ�T����մ;-,��� D�;}K�Y�s�Np��h�ۚ?z}�
vs�,�T���UŎX԰E.�W�\�lU݉}����W�ؿ�*��z�b�s��^���-<4V��1��}:CP5w�>]���@�Kk)Xb�#b�����w��+@��b1��8dy������ ;��{N?�GZ^�X�"*����޲\>�i���&j���^f���j&Ev��G�/H@�䷦";�Z�G��$U\5����l�g���?e���V)�ͮO���6^�>�y��Ҥ$\�֔���b���7�K�Q�U�sfLZp�8�������xO���vd�}0��F"6 '�>)@���t�-o��OXO�h4���VL.�/��Z.+��|8u�R���� ������rf�N�")�����+(P��wɟK#��J��rW���@�=*_gK]3MN�n�.�E-0hk�b�<��Q�p���IfR���n<�%̭x
���r+��;+�ϖ�E�OR�M�Dnk�O'����g��[�>.�6IФgBH�� \f4��'�mCD�����vO��O�o���q���:��*��Bw`�Ĕ�O	��UT���e���WC�Q�� &�wk�	[�L������oY&�L�eՌ���P�f�;A$�+�;ff��)�P�&�	w���B���τ�7�I���TiނGDu��>i .8���G��n�@?v=^Fn��ڽ����"��A��*d�H��f�Pɗ�?5�=�2
(���Dۖ�EI��
��z;�Ȳ��1LH,qj���Q��l�8k�U	���Z�:�ջ1��X��߮[��o�F>
Qk&���~���q���v]�=���r:R&{v>*dt�Ŗ1~��#�{A���������mEd�S+��5�����ktx����p�����5I�G<�8�"�s7�l���x9Vy���A�J���}�[7����ӑ��@(Х�]�IC�i	�(������֌=����]�YB�Q�Q��V�(4�r����/�����'c[c�i#�69�s'����#&�j]���/J�@�v�ǯN-�#�"�!�M�R��͍u�]�@�eǛx�W<���z񷦞~e�ӭD�x���1a�=@�'�e�J~�@A	��kO�E���JvP��l�b�G��c.݊��kj�Q��"��=w�[�$Y��Cڟ�m-#��1���T��H�`�.���2��������0i	�A�v�A�Fy�-%z"��NMo��z�FN�%�?�'?�)���(�>���d�{㆖U���	�F�("�V��"��֬��м�؟�;f����.NߡtY[ԯC�I�f�����Yٯ7���k)}�^	"�OZѶiY�>�z��j��#6s�aЦ|o:ך�c5haSiz�-�Hn����Q��7��G]�����f#[�CU�W��Q`��{qe{�����E �['�����Ճ&/�)"x2iᡕ��^h��L)I��(h�VZB���;
�+)�S�y(�e�)�X� :#��A>�ϵ~���������f��efG��u�9�1�E��x{'�z|��kQ ,��]�E��Y�҈WxE��{���YH?�-�����U�BqU�ʨ�u$RȚ��Cd�?p0:K�@f��#��s�&�ꛣ��/�n.5�{↙I����0�` ::�����)F �ě���W�ɩ���(6�����fnHٵ�?;K���2z�M����ai&���4��8�/k��/#�/����Q�#�Fik��g�G�o��tc��3F�,����iv�u@�)%Zz��e�<cy	z�'�UA2w:�SS��:'������?���h{U�+e���.T �����;9���i�"m�Ly���<ҷ�W�_���4��-<uK�� m�l�@8��j�rR��B��a��o:v�C�Л����s��[��g���"YbD���1*r���-I-w)����2���=91g.�����V$i�C@�����E$�B�Y�!��+�ͩg�M������Y�ܹ �wg-6Q�GF	��3fR>�z�����pw���p�=�z%��M�aUH��<901��[�?1P�:����8~��:|yK%�Yq#��O�ؽ�\�o���Y���i�d��L38��!�a��`�H"��̕�5^���̡ܻh���Ey.8��8�\�{Ҝ�	fM�T�����W'��y��wf��$t	�H}V��w�=��o�H�()�<o�L�����׽I�ʁ���Dv�Lՠ�M�R���_Z�������߹c{9�c_��ܭխ�6�89��D�c&������;6d��3p|!�Ao0�9��7&R!JR�x��r��Q�wT��Lj���v۳9x�
]߷O_d-_�z����r�t2�<Vɉ���{��|lS�]9F���w �%����@�Nt�M�1y�(����68��l
:n�� TF�\��mF��mp�YJ�q���])p�Ѫ�����
h���9�rHt�$������&�Z�U^�jn8oǊ\�i����
�!�1���
$��]�1��(�ʳݕf����Q�6�N3�}x>Aq�H8�<�&4�
�+x_�9}�6U��^�i�݇��mO�K�t�7�d�7�i	�4hF)�3|�ƝxG���2Y�Y5���R
,�V��L� �N�l��]���E�
�T�_�#�/��E��in���,�7�*{�^�ڄL�LA!�����3$R��^�r�j�E�Gh�C}<�"���Ɗ�[m�h��}��V���`o`z{�#��P��r�O����Z�HN����K�Xbx\���;Ao朣}g���vZ"-%�&, }Y��H���XK?��<d��B�b���1���ht����S0͆q ����D�jW���j�(�ѭn���>\0�Y��˝�Sc�ZD!Û���.Ҏ��� c~��ih��@a�b9�ߪ�=���jJH���b^n��7��l�s_E
n�ɞ��R�uHF�����"�=�~o�-�4^��%^���R)�~����Ο��P��/�X�y�.� )����.����/�e�
�iawZz�	lO6Q	;���MZO�E��f��gKT��v��r8�ΐf����jlHd���}Jdź\*M0oX ���,5�QȞȁ2���I�{�k����OQ�t�1���]S*H>O/�6�7��v꨿f	�8��˕�[�Uq���s���g,�<��4�����đN�O���*�&�_�-��� �u����@�L������v��T(@o��&��뚟@���>aln{dN�1Œ5�FJm�*j:¯9���܊1�R���5V��r��Կ��=zѐ�F�3����~���
u�@o���C�y'	�o(�s��V]S�(]%_M%��U�^lA�� =������+U��~W/��X!a�:�EOO��J-��؋�e�\�(~@��!T�&�%��v�'�A��Fc�b��VDXn]���o�ӏ���>�Πi�j�$���w���ޢ���Qb$��s�z�x�|�:���� �k�+��:ԩ�].R����1�|C�N�MX������[렕�R%ȍ� ���@����/$r�F��� � p��߳��ӎ�X�E��g�bRݭ�ԝ����n`����R�`4v�+ܝ7��
�&�姻͕�ѓ�[�aP
Y ��r�_�B���~�Q�!.	�FnĊ:��r#��u�gZ��6����Y�D
W��.#��w�gkN.u)r�8(�m�V1K�
���G 9�O���c� N/��[�,Ǣ���%u��VwrP�h��xS/ژ!��|~-j��\����X䋘Le���ZG�_�	BA�]��g4�h9��fS��0�b蓝���U>����Bp��'�Ǽ���̲]�!�/z\u���7���j�fN߬��;���6����qƓ<M"��?��������>�N��A�[Q�1��6x��a�����Z���d���t�҈��V�V��V�Ü1-�����߭�T#1D�M�^����J�0d���}QU�[1��ב�w�i�����"�����`�|@w�����ȧ�P�y�{J%m��'>��v5��Z$�st��+2�z�\��R�K�OJR��F�<����6��)	���2+��U�`��m8�V�z������xUy;&���ƙK~¾��RT�kv�4c��΢� fmRӿ7��z�꣞@�|�n(����<Q(y����T�J�ufC$��W�W�N��)�4���R��ʀi���u�0�Ǝ}s���� ��Ks;>YGR�Y����fx�=�G��V�:s7_���\�c�I����!]���?�s���1�8��(��4eT6�t��&;�Ð[%a���RO���:7�D`�����2|���ͭ�Z)O������|�4X������⧙���ӗ�hn����J�W~a��g{5s=�Ar���Y�쑟�a�f�6�p,���k65�|	�.��4�Xz���S�ZR�?�v�����p �]��ʌ3 �U�v�Hq���$lM6�����UU�Y�9�z�4'�KE׸»�]�+��kF�r*�4�%YNdж7�Ȃ��}ʤj�RC̢��S��Ef��C�U���8�4�Ո����ڠ܍wr���鲝�����#�
UؾУ]���u�}5M��p}ecO��6�ӈ&^�q��L0V��=#5`��ұFYb�ϒc4���k�ct���M��y�l���������m6�!���P����̅+�Z|>��c�ʄ������R��)%�2Z������������JFɀ���c�2N��4����CSGv��87��1\Y�ۈ��(12���{�cJ �b)X�%?�%����><-<K��%�������9n��f�~�~�v�ʃ�s�lV𺛴T��ʱ����;��6n����ʾw��K���!
�K -�|��;�t^�C����Š�!*�B
�{~�B�%�s�X\�$
5���.��Z ���ߙܔ#�E�N�|���^�g�-�;c:�/�%�������l�@bz��J�|a�y(�?s��H��������ˍ[����$��E���Z���~)��Ǳf]��tۂ(]	�{{��F�L�t�[�:>V�R�d��P��4�sO������Y�gv\������l;Q����)��\�����>�a��ɣ����T�!PC �j�g_kr�q.�	1w�D*�'x���&�����<D=.�aTV�������Ub+�������B2�0i[������3P ����Y)?���$?^G\�G��#���[��d6��oo��(�4��W&�-��h�z�X]T�U��V������[�U(���[��zUpk�`$��b������\t��Y��5��hs��hl�{>ȸ�<0XR���;�Q��p�xijV�)��Z8Ȉ2����Ǿ!6b��#��n5��I?ރ>��((%����/��ˁ�趔F�����ڐ�1��!r
pW��Ls�G�1��.�'�_pkaq�M�i$V�����W�'4E��җ�P�K�l$���㤝 ?����M|�d���*��9L��f�H����7��9���AJ$�щ�F?�vrbr�_D���d������Zj��8T�fȐ�=_�Tq�х(b΃i�OP�"����N��!�H?�}�-`5��biP.<����֥�'vM��)�q3m&��4/��2?C'�S��?,��@�դ;ew���%�H���L6� �s���g���r���SɎ�9Z��=�P9�U?���솝���`�Uo-��"ºr �����B��9�:�ℇp޼T�~�C��i�"������>��c흘mfTL����ͣ2'gG�Fs�x��EQ"���O���ƳD���Cua�rE����@Z�c���ji���c�j^򒿟ޕ)�O�V_'K�*%Ŕ�7��h���-)nO{M�����Si�֟��*���6f��Qg��r���	�<(��w[~�8f�2n���/#G����*�%�Ӎ˿l-�Խ���+ŗ��PH�ET���BQO��O�ɋ	Ɲ{Bo&7LX���$��|�o"��c�4f!0Ŭ~�8�F�K�����'}+�;��?O�ؖ�#m�W؄�w����rl�E!EV�8�{&Vt�]@ǋ�ϐ�0���3���"�L��>2�@���&���c�|zC[�z:�d#=ķD�騍�/dה�o�.������՟{�F$v��ަ���Xu�3�������(����s�1�E�뒆�d��8���%k�ӥ��+/�ll��C���mr_)�_ȸ�Z�q�Cp>��� �`F'jQqrLRJ!�n/�V�^��-�5��hJ�w���0�Q��Ǭ^T!k��u*�1�$�����R��HHn9ROl�h��ߞԚ�l�XS0+g�L�m:Uj��2;�Mϰ��?���L>>-�G$�M.)x���Y�8C����U��
븕�j������[�Y��lҠ�Η��8�{�0ߒ�?l�p��No<������[x�����w*�Q�5��Mqx�͒�"�/١���å�o�=����T��hiTxα�t���{2��X��k��fʭ/�ͩ�?�y��
�a��&I�t�s��2��x����#
��]W���M�Mq��]6��}�0:D�G����D��Ļ���h>L��]Q���g���l�։1��?�����cn��4/��Hn���L�C�5�K��.�뚒��Z�=�⣙t,�l�(/.��~Z���t	�̟��&��T<�%P�.�֧L1K~1�TI�\}����&ҴXe����)JR�TaK�m� ���۹_�����r�pE4�%1�I|�I��gޢJQ\|z�ל�Q���;���'�d���W>�T+Wp�2�1������鶾) �)�?� �u���T�w��p�,(}��䶸�C\�YG��N���?PE	z�QkM�ՋC� �j�#�;�W�"�S�}�P+q����6��(։{���6^qd�*�.��3��&1����'T���V��MvYt�M���is&Ң��^�o.�F�7]C�@��܀z�p��z �� ,���;���V�;uG�	)L�m�p�}4#��-�7���Bpg5�vk�ɔ'fe�^��t�S�6_����ӗ:؅���'^���_rTϨ�+Q
9��]Ք01_/�f߁�7�'\���qAL�{Z��G�R4�wF�G}�1�)v2��Y�eݹ8E`���2(ɮ3��<�j�뚥u*"rb��gm��K���MN��a�ʂ�u�~{�7�<	w�ӣbF.
{��tLf�.��zi�r�"|��(��>R��!����J�W��IWǣs�Rÿ�,�F��GC�귆�n���ق�z�+.g�����!��QsI:����}��;3���P���mI�U]���|�ßY�}�9��6�����c�ߥ��xLG���*qAx�F�?dyb�J�%f� ���L���9y����`,W�~%*�?x�~ �cYt�0�d-�Zwᧄ��A<�\��v���,2%�7[˟�/��2�c�P,�b�2Uȁ�%�y'-�}=�Y��"�U� s)�Rώ�X��Ŝ�ұ\�s��9{;~�����&���r�s�}L�r�8��M�:$�K��+��FR0I�KP[�%����-�h�\5��E��n��� 2u�"1�K#��Pl2�c	�.V�F"���#�x�zl^�Y)̥?��g@��ugG�/b|�>��g�_�w�+�ڒw��v�/h_���'r潡�W������l5G8F�������Οׁ�K�������;Խ�|N��|�n�&[���$jTN��Z��N?{I)�et��eZ%6�g$b=b��vc��u9��җO�S��@�^�s��V�Nl� ��]ec��=��:`�vK�/�':.)� �D2���2T�sHͣ^��V�$U0q� �X�х	әCN��X�`� �Z�/�lX/������8�ֶ��
���+f�P��"����S;2Om&c�}ZAq@U���d/=$�R�_�9��J芄-��[�����9"볫㰅f��w��9�2�cj�p9�&Z���PyHI{��ҝ�퐀>��Y�/�MX���c�-Ѥ��=�i#�k�#M��2=�u�2���
�"]U��aa���f_Kض뮗r�ǀ�7bա��:w	�b��l9�!-L+)�p�dl��I���HS&@����L�'�`"N�٪�C�Y.�c�y���~\�� �aۯ�[����m^V����8$��yB�
j�dr����<޴��+I��4�Q���U��e������&���[H�5ş�.�`䄾�l���c�F^ G*[X+���tq������|�dw�Hu��_�,����b��$+��G�?��B:�x����bGm��T����,�q�Y^!�_A��hk ��:�@*�Z������?�T��c��`!�Gdܞ���$���d#��F�Uݒ�kw��,l�utV:y���4D��t������_3����!�h[�E9����T=��$��*+��e�I^j��P��t������~)���*S�òN�KX��YF���Ղd����C�T���U�����"��΋5��tߒ�s�$ �%��>%,鶑ku�/���ӯqK��q��J�d��B�K��?���=�un��S���WP}םM��y�٦�o�x��߷�	��:����F!�C	�iX��g��VS�Q�y^Y�5e�z-�9b�5��^��%�*�UH�iX~����yk�K�@��|y�X�/��=9�Q>��e?���.��P��p����_`e�1�{V)���(:�{Cnӽh��hJ���z���y�[�)���d>����#mF���d<�P�ژ��i��[T�4L�O��nل8��h�=�?���踅��t����گn�����M��'��T� J��N'���8�Ǜ}�����(��ı�~��{I��~3 P�t+��y�A�Z
�RW����,��Fx�٫�w.��Cx��-0__
`.ĈM�\;���m����ĵ

ܤ�F,Z��kGy��v��*l�$��:M���*p��Yy�n���=�P?�4�[aP�F��BD�h�� �9;]-~���U�8f?C�����E0�ks�0�`C/�X'��m��q�,{�"L�-r��<!Q���>A.��~���	�ٗS�:��BTʉEE��E�Ѣ�6b�4]��͸ժ��2��To�:X�I��G��Ud�C��tp^VW�=�L��j�����+�Tp�}}��-9X@j�
�C���{6R	I&Yd�L>N�h%��]�@�8�-p��0C� D����ROY�(R��E�S��4d�Um+�:��w\�C�<�x�E�?0Ҽ��7��Xe�O�y���+Ai�ha�d2P���IAˮ�w�n�}=_��"D���]Tr��n!v���F&id`0��_��N���I�hh~�\<#ѭ�r@���}_H�wp�Y����58��s_Z$����b�qou�ѩ#Q���i삪k�:�1���{���c��ܮn֙�M��xճ�e+��Z���7�{���c�ȕ�Kg��_�sˁ���RC�l�E
.�d,I�ޘ� W��,)���N�����g��i���*�Ii���BJ�52�d}bu�(l��d]W_���:��t�����&+nvYC��Dr`:��}n�����<π_$уlm�U-�M]�:]�_j�n��7l�.�A�|;�|%��~�j
f�}�.�#�LV�K�����_��)�%�9 �7��֪0(C��Ը��]�r�@J��N��|�����H�um��)/~k�-��au���%�/���2�;��S��� dl��7S��1���LHҜ��ܤ��ފ�n�W�=Q<�ӟ��w�����	�&�R�Y�2�!�ڽvH�j\�7ZR�~��&��g�zCPV��6�ǒ���2���aM�G*�c4˺��
PP�]��Iǭͻ��@��m��<��m�¤�"bp� ����8��6dZ:��D�)1n��OڋS-g�nL�V��}Ofp����q���H�ܱl�b�H�}�zl�&FLm1V�U��d�$�]��h��ˮ2ӻg�+5˕g�Şl�+����H��-D����k�c�<��!fMZ�HG��|r[@l��ioHJi��vQ�yv^��&Tp28 ?w� &2�$r���&�[��QW|��-�����Q�Rum����͒HG��N����&-����T���d��[)��+�|�an>���g}�������b�TB��h�/��Oe�����Q��P�?9�[�2��P��ړcfS�U}��~��^�D��c݁TC�#���ⴙalH��1��\П�x���$wz����m�Ln��5�X����:k���	���pQ{�.��c=�1^3�>��~�A�̕�0�},Ȣ�d��}�͛U
��}M$�m$m��!�Vӹ��#ģ�#/<�+(�Nxqn�{>$��ᘽ�����k ٍ���D� ���yP+'h�[��+ϑK�����G�7��,=���fG�  �Va2�B��t���y�P2:z2��w�V��!�H��
<9%�{��HN��/�
����;���P��4�~q��Û�Vt>����x���ӈ���C	 ��F�'�L=��T�=�HL:愍�7A0��O�~�,<����E�G=�n���*����HZw��������o��c������џ�tw�w��K)�|έ3��/l���ܭ��V�;�A�E!2��g�f���_�~_4��z^!�����#��!>&�j���~������V%_���n-�G.+�ڿ:��li�/���n{ro�Re(d���/4���Ȅf���`�*=�:�	-@̄��t�l*�y�L�|*{��\	Yբ�3���^]yM�Ke8X��oV��qt�s"j�o{��hq�1%���m��Y�����ٻъI"���CP(�_C��-��}�c�#G���B�W	nt�xtz�>B���7�qG�{��!��
�M	���A-�#����E��_�T�JN��qo�Ѩ�����},���~�֛�t�1���
Ǫ]7�㬚�������sr�,PpXY�@��&��Riy;&�I�z<��K?�ch�SJv�ٞ�ү��-��:��b/��H�W=ɹ�'����֜wے�;ze���L"T�mv��N]��GK/�-&��������s�4P�5�5����E!f<�b�a�ܻr�(����}���`j��[���ɻ��UMpt<l	\�rA���1�B#?R���yV7M��(kXO7,1��p��n���xL���:5N�S����G�ܸ��cگ�&�\��c$H<�~6�ˉ��tX q��	y�D'�J
�҅?�YS�ߟ��z\ Tک�np񼆙��}�$�њU|pv��~h(W���Ϫn��-
;�����!ݎⰩk��u 
k\n�:<�x�;J�Kgu�NX��V׬�?p�uK����us�1
'z�ܰ�w�Z��r��U���,��O��N>�'�Oh����)�1�Ms��J�d`-������K��V�xv
�7�H��b�7Y��ᵣ"r��I))?sgb^Q�8�e�����b�8J�ĭ���B�u��+7��'���S`�Ե����3ۦ1;2���[��ZHH�?�D�`kt�¬XW��={ܭ��+}�1�������V�/�`���,6�Bokt-L:2��ҙ�W�Z�N�+�����N��U�N��s���/Ld��i�t=V��t7T��GA�ö��=̇0��)�p�)���ll����@�l���xE}�_KT��"��m�z�/����s������m(lb�4~?P7;u�#:�0�.6׈#.<N�b,����~�x�O��Gi�q�r<�ܭ�G�_�r�,PW�+Qr��]&�yz�d��۵�� VgMҏ[5 ��.�pR�O�B��b%gw��8��{
� �yg��E �G�L*c�2G�ĎeȨ�TP�(�rp!��	��W����YJ�~ܟ5�ˉH�<�,�pc&��|Ti8DcE�?��>������U}� �ǲ�*6HW�d-6m����=�в�H���)�/Ł���r�%��K��@-OK� ӿ�%dD�m}s�ST�<c�,���� 
rA;{�g��\�<6�%'�Emؤ/Z5z*:׆��B�5��9 ���N�9Q�ѱZ;� ��;�f��D�Q����t�B��K}@+P���U��L-=�W�C��>�h�`�����{�e�V�y4��* p���]>>� ����nUʵq�@�Pl�1 �0�B��G9�����ox��q	^sز��*�Qi��f�o���)-Aͦ�
x�Htl20�ul � �>��{֞[�fI F���'%����^p�G�ǐ�:�