��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� f
���O�Q��Y.#�d'���J�"����4���d�"�Ŝ9͜����
�~�a�rN�����o]y����1���nJ�]s 3L!��,���zَaw�{,���{�b�[;ҙ�u�\��������.7���}����H��ΰ�&���ے9��y��y����͍2��ё(��7q|U9��1���i��$>�[�G���^#fU����S�"_a[7B��7~ez�#�5��-������>[{Љ�v��G]��Ew4��5`�|x}��4�y�z�f�|#�դ�e��5p���1��L��d=�㺔��y���h����V���Q���t�̿�rբ��6�j�mcP�iT
���c�j��5�j�KL��tlV��d��x�Z��"ks�kCK�|�i(�;�����6��12�XTeP��[��'�0u ����r/X�<��/�]Gȥ���%N��]84����Uwp)
���un(c�Åf��J��f`9Fqv]���+�<�w �N��fѧ�h ˞�C;4��#�i��T6n�Q�T�����ڸ}�rS3�*�x�٨�j���y�~E�s�~+s�G��'��%`+�w+.}��(Jľ�$SL�2-�M�M�W5~���/%��t%���0;��3��G�rq�Ħ@];
!}ˬ � C_3ZjT5�ъ���29L��>ԡ��I�#iDn=*oB'R�؍����v��< 2<���oc�M Yx�R5��ܡ�����2=ړU��oLW9oq��4S�um줂f�X+��t)�a��� R��M�Ć8��,=���LIQxFjg�f�O����ҿ!.j�3�+��G��[c�6��܉Y_���+��9"L(����͗F�CЏ�� 6�vWm}kd�����܍ 	=��U���7:V�Y;��)�h;K؟5`!F~7f�/ *��.}�#0g�e�s �	4+�BR#�'][@VK���f�`���?�s����*�w��>Ъ�3���5�	���']y�?��IFgƮ .U�7q�]U"΁l�ߓ����Ѽ����ӓu�pO�vᫀ	�� 7��.�������^z�%xM��f�*Fl�h�HOl��I^��������	&�d�_��� ��޸�٣6|)�C��;ؐ
J$c��'Ĥڕ��n1n���۱V����t��V,�	k'}q&��5���1$���LP�ov�B��GO6��NE��L� �����k��H��M��&��s��|)����h��k%E]��v1���ş�s7�+ɫw���t#����t/װs�3�l��B�;m�����;�x.u��u����0��VP[n���Jxa�);���)q��|%�����^�1� ���?=���:�0�C����ю���o%՞gXw�(ț��՟�t_��e]Ι��"Pڑ�;�X�>8fE:(?�ȇ��d	��I�8@U�&�g���h�C��q�ݳ�p�^�g�s3%M<�f����Hg@���Ȋ�a��)}�j���$�	�XR�uN~�s�f�n�}�0�]U���u19n�Q�����ď�D�@>���������t܌����3-�T��s��`���,���,Å��"h��$G�[�@�����VYC�$�\��{�˂j�7�Y�^�&����^H�Y�X��3���G�Z���3y6�+-�������*��Nq�Ӯ</���!f����O�F1�h�d0-SQ�o&(��?t:Ş$�
w:ś��*z�1)��z��ұ�P��l]��	H�����/oo}/�����X�^��l�F���Z8,d�؃�b���'w����\�m�)�'q��^$�՚���%z���}v��Bl.)U�$_QD�ԠwW�K�o�ݞ]�>ù;�g���Yu��ت��"�jW��_�3v���XZ�
< �YPH�b����LE$![�p
|w�[ہ�y�d��3�K]�[g[
ŷ�#�F2a ���oU#�i�Z�)��j�90� �qx��6"��6��|[�l�%w!_�A��Hw<�\2a�Qh�Xף�$���.�r��g��k��]��ړc�vP��!�q<Ϻ���2&��W��-U:঳su���%L�I.fs� "����9��-����b�%X�Z�W{F<�:IBؖ�kBr�P��Ų+Z�������g��PK�?� ��$������,(՞�Rf Ka��5�<.F&��o��%�K��xc��\��4�>3	���E�郈��j`6��&Vk�\���H������$�d�2D�(ޮ�gI�C�C4���v.mb�[�˔�T���m����sXt$�*I���-|s�;���0�}CN(��\({��F��8�.�3H�_J@�w�L�d��r�Fn��i,�~(�	��|@ʾ�1[!��#����)G^�b����R��1K[aV�r�O�,����@�"��cF�".w�>�����<x�h���?��~�}�}�=w���ٞ���;�ZL~U��iR"�P�&�ֳ�����9\���^� a�!�7^K|�oJ�{}�B�����kv&U�ĸ!$�qZ�����ô�x�U��g����=^��믹��ic�"Ym�.#�I.�F��)n�ɂԽɗ&F-�e/<\�bgJ�~dc���%�ݯg���C�x�_wU5�V͢�<V{H��mzNp�	3�@`7���j:�qqa��A�,vڥ����/��ә��k@Q)��w��0 uɢ>�.43�)��P<�7W�{��q��/>*�<U'���TbB,�����9���F(�)9�`��J�b�o`Y�q��E]"��O�ݙϛ���ih��z<3������30>Ox�ѓ$�_XzQZnl�}W��p"G]���gPP�{�m�\�V�m����>뭨�W���"����g��~����y2
h �m��G�<�Oa�X�h:w��;u��^P�D�9n�]�����j���X=����io�b���DI��C�wޕ���'��v���sЎ���BŨ&��L61)U"}:�~���ǊF�]n�Yc�D\���¸l�c�=w�~�� �͆[J��~��&ұ�N�\n���ɥi/������s�0��Vj��l�Y�� *�wd7L,T