��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��X�O��v�)�P?,���89#�Kw#�_>&�ȯq,�0��V���߰�+������bߌ/�h���=�
�?�h�A������[��e�6Ǖ�ǒ�I��H:6��2��d�3Ȭ�!5�,~����o����b���ʅ�Sq����8a�,�ȼ����n,L�)���dO�r�l	���HҔ=�!�N�*�-?��Q������U�����7=�N��2����b�������r��o�1�t󊣆�0�O�Vݓ?�,7��u�W���o����Q��#����r�� rv%�MMwmq�;��GL|�ٟPK���'��#�[Y@�W]0����ڵ"ȶn硨YR�5޺S��#��7_���r�l9�S�W�>rD�r����,�{���RC��lI�#;F5bC��`.S�-�$2X����4�.\���?��C��.`e*pӣ����p����6�VW���l�B��.��*���E��<��!b{�tP�0�t.��z����������Z��o�Ny�e�bL`��;Mrӓ�4��xE����U��D(�{�@���cQ���I:a��BڊL��%r��?�\��m(�� [d�<��U�S��Kl��-ظ��X�7cb;��tQ�=r-������ۿ��}b�d���-���i|����)�Z�|���WJ�D��o�Zhhx<�i���
�ړФ�J�tC5����y#i�i�xr�������<RLMW�Bn�n��<T��0�^6����M�"E���S
c�4�HOT3e�#r�U�e�glh�yOV8��BĬ��2�q+ȶʏ�����Ȱ�v�9�r�!;>^<��l�����C>�+�M�BY�Աr�<%=���8I���b�c����)u��;s��i�m-����{����g#�v�vYhna�(���7Ht0sd��|���٣����i�A����(�S��}z;��{���'޹�P�t��L�n�1�g� �~_�X�*uDU���f�9u�K�������!��e8��;�����=��ʭ+��r�-b��?IQ�%���Vu�I���k����P=(i��4�ᨅ\|����Z{Wʛ�w��50W��g��iU�>z1� ���\����X.���Pӕo|,X$���]� ǹܘ�b�J| lܚ�Η'���B�	�yC�X���u����+��v��ٍ�g���p��TҔ�%BJA���K3� EƬ��ĲC�d�M 5E�+������h�3<qM�o7���2 �\Y1��E�J�T��\�t �)a�;NAf�R�:ŰUWi��6J��Z�t7��ǂԝk���;��e�It���7��Z��lg3���]��7����5T6}i2���R����8Ё�mNK\Q,�:���T��`��� �(#)�6�Z�z�M�n�:����g5'��D���k6?�d�:���~��ya�̢X_J�c�k�S�>$���CO\�h�
~�u3��<<3}s~I�VX��3�?��BG��u.�8��-٣[���P�+��Am� ��']R_�>�O�����Z^����ܷl�j�����u9��횽1�P��T^�7�$�Q�G�\8u�<��.��Z��,"v�JZ-�qPs�I�����O��%[�m7e9����D�P�?��
	dZOk���ճ=�̰���D�֩uws7�"1�c^������� r|/���[�mb���l��ӳN?���,<��9�_�F�ھ���>y�Q	�Q�M���O����L��&F�D��*�S.L����Ұ��O	qĵ(I!Ij�R�OmPbj��Ͻ�廠��+Sz{O�!qU8�q�K��Ь����8#25SA��G��$��_&�����e�uC�ݗ�8}�����/w��?w�{, nc�1�=��G�#��M��'7J�a��5�[w�z^��ʾ��7jҼYh�OH�k�	vl�\F��-Z�v ���H��5�޸�yƚ�+˚����7� �n�O�GS{ϭgw�hh+�?n���D��p�xn�ǉ q�G�^@�F�߲�F���D�i39�,��%�۞��@�+(#P�g���A,�t-᧑l(7����,���|2:��b*��ٌU��K���4�r�Wk������$]n���a��?��?e�X!Bk��փ���E|��q�U�x�)8�)?�uj�o��}M�!��{���TƐM	�npc��V��%\�e�&Mdłl����/۷����k+{:��?�m6' +�XC6^0غa�c,{3!U�U'��:p6Q#��/DL#Y.k�j���o7�M5�{@s�����"���D(q/"�㡘��	e8o
i���E)K�v�����'q�X��8ɜD�6�l�M1�~X���Z��}p,2K���ړ
�gw�^��I�<�9�cS��JQy�[�BRÀ��!׌~$�*����*;���loS�����@�n���p�"�f>^�8o4K�m�\��JCL�Vdf6���Bc`�o>��Śਭ�<�����>-ZA1$
�i�"�rI��:�հV�H1Jwѧa��X�+jوh�&dy�W��b�|Ov���$9�f �i\T8k���ѩtl���CAw`*qvs���Κ~��cN�<�u����7#� aټ�z=�<u�YV2�57�#�Z�ь@1Ԯe�iT/T�}�8�|J؏ysC-^Y�nWw&ƇGO�mK����*�hq�8 ���W�rOJdo���9�R9�� ���&�oy̗��)��� �Q���kdY�L�΃Ox'��j+?�5ā���pfj���Vr"��T5��@��¨t�P��b|��nMQ6��U��H�C��$Y�X�8gU�y�N��}��.;ÝX�ΠlCw�	�@vùsy���?�� ��M<2�����j� ^?Ex�aRQ���{+�6��ܨY��*�O�!�E$O��I�R��W�a��T�K\����}���:�����t�U�,��ߩ�'CL���)���_��4�3��y�^�*B41U�"y%`������*¡���� i��)�	���}f��7�(������f2l���v�FAo�� �J�.��������� Q�:�DY���E�a&N�8Ƒ�r�?.�F&R⯾��j �����˧�?�a�C�Z���=ݼg-��yO"���:�*�y�cf�s>Վ������\"�p��D��%R",k����&�!�0�7δ��?�'�Q$��5�،�>q�$��s�U������O)�_�����O���l�k��l���d�+Kcu#u%�ϧ�&����b�C�vp�ʦ��[f�9^���,�>�aʏ���c_z�����va��5�M��Lr�#C��	�U�CN�$M��z�\��6g�G�a�k�-�Һ��ld#��>'(B���cל��²e�ɛ=jK\0)�8���h]�Y@�(�zT8<ˋ���(�� ���7�r	:W2��J�ẫ���lW�����7cd�Sj>�����)v���aլ���� wK�!��u�"׀1`�
J���v�@j��ڳN��'X� 0:W\��n.O؈�gzK�<Զ��b�F'���fIz�Ǥ�y���*w�I�\�|� (�`�R�je/���j�<mM����g�z]jb����5YǺ�䧫 ��]����ux�K�ºMZ?����dzQ���{��X�h]Nה	_C1��J�5�:Q�{���˞
 WS��.B�#�/�l��$�Þ��{[M53P�ZF�k�Q�"أ���|��K�n�G�£J5�dL�3;���7}qh��ߟ<�kRk�=�>�m�>uȤ2��Mk�&]��n�Ci���ŮŻw���v�F�Pdw�)�@K���P�!�$*����u� N��[�|_��&
�mZjC��u��h���'ؙz�9�|�����)�v��Z�FZ~=�S�	���篝l|�q�J7�����Yg4���y�_�4��"�1b��� #
�������� `���ݙ󂺏mn'ˀ� ���K���Iu�hR_��()s�_Y�,d;�NA� ����mb��!��ŧ��A8��~�{]�r�������4ޛ���+��J]ha��۲�jN�Y�v�?��q���X�R��UP{����¿�E.���H����-S�ě�(o��Y�d����`���A�.5�#D�(��{�Ǚ5��}p�m,'Pb�,9C!A���>�
�!�C��Ϟ�
I9���Zֳ��]#D7�~��I!K�I�h?,��=-�d���"=Y����P��Ҕ�$�E)���X������0?�R�Ѫ���
�.KY챺ax�.T��x�����m��H�%��
0�#�������%U����׏,�9/R�y�(��;�m{�&
�z&<�.���L�3��v��m������e:� ?��>��1e/���$Sۚa�S	�u�o�"6[�Z"��*>�� �)��p��%�I�L�%7M;.Y�J���,ө4��(�0K;4���)e�*�>�szQ���-�ȝ�h��_�p�5W��;��j�̱-�����Ehi��>�ɣfl�R]��IS�������@�t%D�ѐ�-�-�b��oMAa��٠�0;+֕�촀K�r�Ԇq��/��Hw��^г��o��ŭ��ۻ���\��gu�����E�'���]���q���
��B�V�W�c�v)�Έ����0t�F!��.�#�3�ؓ���aᆊ7�tyr��Ps��n�O�ch���Ն�R�V^����
j��~P�7��7��O�O�E�A@��K0���,�����vf��q��l�Cp���=G���^�+H
G�3��;Y�pE�f��G�g��m�J\nZ�0e���TKR�)Q���_� �DfQp�?��ms�MUtx��A���ӻ��>����ű:k<$�P:���X^.;�s����s?�A��1XV�RQ�F�:A�����:��z-j����|��[u`�8�c�:Ȱ5q))�菜j�5j�Y�ڇ���<�����(Gp=l@�S�Kmv�X�E>L%P�X�E�Y�n�7��h�����|��L=��d�d�GTK:O��c���N��K$��"�x���O/!�f��%�iW�^����:L!�p6TP�pJp�]�Q6[y=;�ܕ�,@��i�(����?����௉�	~�:������-폡C-�ǻ�X���T~�?���~��&!!�#�������ۂ44O<����G�V�0�*߾+y�����j�v��,yi(.?���LY�&���Q��/�!m7�f~��r>:ՄN����r�t�l�����/���j�����H<���G+;��;hf��F�8k�C�r�$�鋡x{l{��l���$\0�����i���^AC�C�x���x���i�J9FrV�B~�W ����ʳm4k?'H~�CI�ٳcou[w5q1�My�OޫZ�� K3<
��;���s���#\c�-��Tvft&���7T��s�=v�<�@Yb�w-9w�1�l�:N�\�92�n��Ж�􉁠�@�e⟀W����q��2pr<�+m�š���*�&S���)���jX��V���a�z0�Z⭫�h@���L,�V'����/2����5��*%�))b��s��W�C����c�!��d=���a��� ;-�wW,�w�Úr.)O@�Yy�5.����p���wm=�L`�jg9�wY��#�#Q5�qYw_���~��'��-���mx�L
b=�q���A�;�O����\O����l�8�Y�y�}���=qU�J_k��@%h�-mc����(D���2�da��7V$��$��/��8���7N&`q��G�IM�x��>�$C��w���}����-l�������ԕ��(Ƃ������k5ۤs5Z���/���4_γ�z����M(���Ry�'LZNe�C>s���J�/�u��p���x���&�]E<��M�=��2�莮�r䁌x�eE����/�b�X/a��t�~�˩p�K-�I6����7�7�[��L
S���Iy�\wɍ5�cj2lJ�ĠQ [�~¾FqT�e�}d�g�� }��*�Z�E0DJ۶��aۛ_�!���G�a_��X&R�f�Ȳ�~\���������^����ߐ:s���+Z�AK�����	�Ҵ��A?�O��[׹ˎ�%I2os�@lh(��;��K �^���|��d�K7�х�)�G�4�����E���]�V7�^��R�d%l��+Wg��1�����_w`V�(�6�D%m=�.�*V'���U�}�~����]�W,g��vƟ��H@���`w�]f�.�+\*=��^��y'� "�~QR�x�(����0,E��ʹ;"�w4r}�/����3�����Y~ّ$P�J�� �5Qr�\���秉'�լ�Ͳ���`��
�:Ͽ�ݍ�QU�B<w�KY5���%K��|�|�W#��ƅi�c�D�+��tj�<$��@Fh�>+�X��%9��V|��`Q̉����-�rL1��z�[)��-F��n��#i��G(����'�C$�����(�H�>�ci�����8�����f��jNu��aqk uռT<+�d?]�R��i���:���*ؿ墏�N.��.I�(  �6�(�B�Y���V�;�i�KT�2�����ߌp�K�="	�h(Z�N�z�@ 3يM�dC�
�s���Gv��I��`���_�*�ZL�B���6cӖV��*y�QzRĮ�҇Ӽi2	�y��~'AKJx@ ':M90����1����W�U�6���3M��=dO�)��������6�sH-&s+x�}<��R�1���[�#��Y&8���l�,��a(~�&9���hMvt����q�����;��J;�vq]8����:��}��	ǯ$d#1����D�$���&N&���z5$69岖Q֌���B�>�]A�]��<�߹v��5�#��.
�Xv�**���wV'\�B��@�rY�I��^!�M�<'4���[$��U/�����}�щ|��lI��͟Yb��0[���P�M���T���ܚ'�����J�mj]��d��駸nKЉ"���n0�f5���?�E���絛�Zߊ{���U���!���d��H��3R窻	�0=���֒aF<�:$��:\D��w(g�H������1�EX",���W�~��F�le�T�)��{U���)��� �KxN �op�D�`�W�\:�h�b�s��5;��U�ʽXia V(���)䝯�?�~�G��f�֌j1�m������Ê����6�8S�~o����R|�����^���ɖD�f-b�v�E�
2�8��OD��R�vt�NN��������`�o�[��0%�xW�Kg.�Vu�@`�Naa���Kwr�	4��of�fa�jgӚ�'�up�ِO�M�������B���lw������Q�1�E���v")�]���b5���$� X�������Tp��]��q�޸�����+��w=�W����i�����3�nw0v@^����]��		��;�3�yC�ixM��<#'$;�)O�w�ө�*���K�2����F�n�P�I� J1�1�hW T:co��zbS�t`Z�b�5�e�4{�^�I'Z��c}�X ����ʿ*(�)�ĸ�#d���Ԫ%�u��/5��OF���v��l�Cj�$Dz���%�_�m��j+E,Pah9�q*I�[m ��xR#�������"��YLJ)!��h/O\,�k���EsSj��ɑx�M���a�AT������R*��v9���p�p�T�P�f�)uY��w��iж�@��,��΅���XB�Q+��<�ڗI/yg+����L�f��d�i��Ɉ^�Đ���e1PQ��tC,��q\���M������>��W=]'xY���aI��F�ze�5�]i62�k/d^si�R���u���8��������a�jC)g�:=���>z��/l�)������S��9r&;�9�kSkk�j3���Ov�Ѭ�3����Us��e�ԎM����ݘp�i��!>;-�8���ʵ�n�$7����k�(����|��ȧ�Y����B��OgQY��2�?��^_5�aSgs��O��T�,�vS����C�����-̜Z��__�!�c�k�e��]�໒^����a��io�	S�".	�Z�s1�%5:fN�T���¬ǆе��jM��'�%����xUaG@Lf���4!fH&�����=F�eGQ	C��l��]�E^bsɃGH��L +������*<j~6͵8���]��n�?`�c땻�Y�$�R-�7��ut�r9� �Z���[�*~EN�G�E��KA��B�(F|�gF�`<�j�^�EWڝ�®�M�5#B� 1��=?
�X�����i��k�pZZr2�+� o��;"�	�h� f��E&?g�F���4PA;ۣ -~c҃z�bޠn�%�� \�	�2�za8d�\εM
~����қ雥��	�9C�B��`��@�\vm;��>���$�S��/0� Eb�g- d�C��Ixw��S4� Q̆�2���9�Y��?P�\��Y#�yH�L���'�p?�dy�r����8�趌x��W�8������[FI���-\��@/�ȭ��Bd#����o��t��ݽتe�F�)]���?ک�Z
vD��H��sV*��V�Ng|��M#Rq�}g-�@-��/�+mna�ΪΦ��$z_y	�<zy9|g�.��!��MZ��X�0�R�����"w��$gHF	Fo��Mr��$�HG��c�k6��䡭ʉwv**���
"o���^�z�4~�؝
�q�W9ߓ}d������*3��9�Y�Ki��,+4�w�6k�E�/S�w��p*�Q��x��!=)8ï��,a!�f|c:SaH^�xp��Ȱ ;" ϸ��"ҫ�/G��x|�Z\f��$m�|�SQ0��
#�^����%6�5J�N�O��p]U��NTn�H���xߟ��v����y��O�rӉ��� �P軬	�Ժ���>��[�͓m��x�O�_6\[75����z�����/��6d`9��!r�Ր�ٱ�X��3�%��u��&Nv��\:{���L���Nt���= �o�f	�]Z�3�L�A>5|�P74!ס�O��¨��n� `�V�HkuT�y����Z)���]r�.T��"���� �K9֒��a/bz��%��r�u!��u�.�*���1/�K���Ӛl�!� ]J� 4D	��q���0-�+mP�p�%r[2�Mk������WP����74?
=����% w0ӗ}uU���0��*��C�ر�?8~�t�Hu�yL
�c�|;LЫ.b�m��ʹ?}��<ޗ���-2G��Ŋ��fT/��C�ж�	��P\��jG��Lˀ��k�O�o�[�,~�FR�ts��2�D��()?h�8��P�#��ߓY�R��ݶ=����ڄ���W8Gg �f�M#J�E6�Z���Ay�fo������GC�:N�Ɔ��eo�
wI/�I��S\�B��U���R�Th� �f)Su2�/��j2BA���O���o���c����8��z��n�������v#���s}-�k�}�g=)0I�,K�[2�tn:Vj�ن�𩈕ߵ���"�!4��נ��4í��q��j�o[̂������6B*�Xg��qv���Ty��eX�#�����Z�)V�ml��!tw��N���q�D� �� ����4�y?���c�ʄ�]�\1��"�*��}���Zo����>�t�sd5dG��aլ�B��	^�G0��P�?�Y,XMc�ND]6}�R#�i;��٠z��9���k���
�=W;^&b�]tTd-1���"�ۙ{�tj���P� ~�h�,֟��-z �_�Ry���O�^��㑴}0"�\�C_Eh�S��a�`�6��]�lҩ���9���o\�$�N"g�ޚ[�[lD&7z�>Gn'�v HTc&�Ο��n�۸��9ŋ�{��dЋ^�Y���B�<�;�^ �h���굂�g�����L��FK>��sb\OC��M�ۊ����]�u��I��I/�j�]3^�攕�w������z8���ً����2�㪊� 
ٻ1��~y[�	06�(4��±� �UX��ŕ�f�'%�S�5�f}��R-Z�Yd���Ч�]�9d��)L��j$k��~�v��7>�Q�-ԝ�?�JNr(��]H��5^�I��
��'����SM�U�K����E����-�1�_l�@}I_2 �p�xR�-���E�@��ԩ@���v���|8w�ΥВ��4�	�����H<����)KCg�t��`��XPf�WV1��lL������e�S�;�RE"��գV�&�V�9���YD�N&��+]�O����v����q��yR-x�V�*K`\fpŇ&++$�#L/k��*��H��a�Ɲf	�Ʋ��d�㶇O�Q�x�y��X����W$�t��������	P��aε�3�`1��u|��s��2� �y'�e���1�=vy@�6`��D��Aa��!38[ű0��#��b�$�\uw�bi���U�@ja���zV]e��|�'`a��Ѽ~�W-7�紒LI���rj>a',Du@m2}�o�a+�,'��h�Z�����N�R�C�F�����~*�	���U��й�c�����i
X"��ߛ�����c�7��<B1��`C���8��m�����.�C��Y<lr�:���>ߨ ���$��˛�@>
�l� hi9T�!��8onz���'��:OPƅ�3���ZI^���L8(Ht�f�u�3�
p�c��Y�T�o���]�K��N��^G&W�[<�+J�\\S9(ln�z�w	����oKÐ�o��}��{�K� �!s"^���!��