��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�^���x`��������"K����J�=2w3�
e�gƨꮋ5�;��`����I�}�ɱ��N��5�~4��&��@Myl�[�����s�z���ݙ���Y���M�	����>V��k�c�>a����ِr���%���@nΠ��xƦ_�q!�{�/���rP�'cGı&̕��!��Z}��uVe�ғcS���	�텟[�lc�%����xS�ɅLn�q�W[��إ�Ɋ��`H��%x�{�T�^��Tj?�N4O#�Ty �K_��`_�a�}Jشq��c��*��6�+/��L�S2�Ӽ���%+�)�����t`��wG4'd7�(�%�rD��O���`D����T�	�� �Rf�n���Q�"��:1�8H3��A9E��\����f�FՆ� a {�;^ןw{�4stߋɀ�R�X�bS�ӆ.S�����u��cXte��*&��g�^C��5P�� S��-��h�5!�ݲ��/�)�8�g�68!cV��4�@)�ֹ����r�����R���������l�(Ӥ��`OYW�6�p�"&]�;�>�z��Ie�d�@�U��x��i��}�wA�$�����Vt�8pg��Nǹ4��	�����]Gx��k�������U�����8�?�N%u咻b0�����i^��X��/
�%pR.K�P����+JS�o�d�d���:�2I\�zOV���4)�ܐ�v��I�
8	���U����YD����昬�vs�՚�j�)<�!c�@i������1|��*E��<#��?�D�f:@��h��QCm �@�!w�Ց��*j�Q�Tpr�u�p�� hE��g�[�o��U��&̤�7�E���/��-�d����Y���Y��Q�,�`h��u�O��M�9e��>W��_0����},i}�XlOŦ�3�җ�'��/���b�����T�Ƒ���?@���ƕby��5��`}$�#��,�4\��;K4����=�'���p�XK���7���+/fl���n�g��]ɾ�0�m+�<���in�G;= ����l��'ڷ�-�	�hr֊U�S	���YI<��â��}�E��*\~w�*:OA8���UBXo+Ԓ�t�$�_:o�J�z��NIP�bӅ4jTU�Z�X��êÇ�?�"�(�|4�	x�~� i�oU_�S&�Q��({�qe�@��\�F���@��{Z��.�s�~�<nF��aʷH�
�������.Hn�_2nb�l�o�����-Ul�Y9t+ۄH������t���6\u�8T5�5��w�� 7"���M(ov񅩐��m3m�W|���2Ք�{.P����?���8��8$6wr��I���!>��T�(�9��E��K>�AƄ)5YQ�19��I�z��l�A��?��[�@��_��*��!�C�����Hۤ��Y!��ۅY·�=�0����L��g�����ط*S�L%����"k{��¨�bs粧f����ht��[:Ӑ�k�D�$Jh!�(i����ъ-����@;>yҤ7c��w�<~�s�5�fYN֤�"�E}e��k�biN��m]1�
�\y���T�TX�4��`�=�RV��HG���N��2/Q˞��|�+�@������2q��8��!��Dڠ��_0?u9���>wӽ���T2��
p��
2��~��J��UdOu{a��sKz'�3]�@ǝ��G)�Oa�<�= �{�)r�P���4���Gԗ��8�t���R����R�kxP��U>I%*�>�:�FS~�@����fI&Y�
�����(�;2n��m��;��"1���G!�g�x����c�\�;��Pfˈ�R�n��,��Cʌ�IS�塗�L+�Ĉ�b���Ͱ�ڗ�����xp���(jɲ��e:�R[�Ț���ٺ�c1.�����W%���
���u=���ej�.�ې9�Qa�[���o՜�J&��?lO��Y]�6�י�<���@�R�Bl=����O�bJ�S9�`1{Y��A���M4c�� x!W��3X���+G�T��2W�%��a��A~�P���e8�����'qVNr� *_w�I�U<t�{l�-�ޥ\;�8�G }Fn���#)���_a�.�U����rd#�ܤ�+�e�ݨ��� �s�2T��O��-��܀k[;�J̏fZ��)\>����0�;&��:���m]8��s�w�_ҿ���j<=�3K���9�FE��]#��ۜ�2���� ��fw"`N~�Qꤟ^�Nx.�?(�W��r��h��e�i�����a̿��j@>�*8:r/�ա���h�6t��4G,��f�Ə��sk�#��[n=𥑰� }=:� ��	�����ڣC���G%�`��i��|8۽��K"��Z��bBy�n��۩l���ܔ:��Q^C��N�N��OQ��t�b��q�Kk+�] a'Z����:��r��P�"���A}8�y�YORq4>)�}6Mᣔ�d���U�"��Avf=��kڒ�9��ݪ�)� ��B#;��X���qF6�k�?�r�R�$�6�'���Ti*	�p.����&&u�qg�?Ը}�*_X2ߛO�\�jq�Ve)���^�FZ%�(�'.��:?:����z�Q����� IC����Y a�eins���\�Fn�-|od�GS�'WO�٬���)Y�\�y\��ѫ��QG񆭪 �F�M�V+N��du������#Z)'�Ʃ��n ���@[m���' ��B�����e:��af(�]���W���6��~&Z~�G�B��n��-���*����(��&z-. ��2�)�׼s5HՓ�ZhH�94\kSaE�T8$��&���@<{��\{Τ����ش,Zfbه���P�4Q��,���و3�_�wƊ\X]��sfz}��I�C�����0��]���_������蟟J/�R�8+�![t�j�S:  �.6N�`����u����N�'�"�ϣ������o��Z/�\���@�\I�X�0�����S�[@4����J�q����̒�9�_0�֏����q�SR7�5���c� ���I�%
l�g�;��ig�,A{ȼ��$	�RI&,�pa�jb�D:\}�C�%n��n`be�'�9�W��J�[�L��?hE��0p��=T�Τ`�!�]�#�Wm|��7i:��lw�8�hf���֞T24+�I�[A�Ð���G��{e0��z��1��BK����~1��
�p/O�T:������=��3}^k���=���5�����gʶ�^�g�u?������h��|T�Hߤ���^��,A<x���y��%�P����N�%���$��2שR�r��̼�j�j c�4g޻�K�
*��[�-;�d��"n1�c���6Q6��s7���2Yck���|5���R��r�Z&Md1����V�+H�(�;���p��Y�<� �GmK��5��s��75n�374���Ja���N�e�=�X/-��it��3ilL�#V���J� ;�	!,��}s�*�;�8�]*�D-�z(_���
-yE�׽�"E����mQi�u\kgo��d�q����ac.���D�#�S<�D����?��H�_�%��r�,���I����F�g�e��M����Xn�@̪�#�*|®\��y[�b����r�#�댈�*���įq�`k���g�3��kr<����5�8J�)��(��IN��8,���BC�ح1�Ǭ3=�%�{R�0�r��2��w}��X�I�;J�ٿK��϶3�̜�(b�^Ǎ���<��r�^�,��j�60L��D�NL<[ɑU��s7�Q�m���>�8ȇr��bs�m# ֟}D�`�2�ݢcch��Ν`�B;�l�6���o��[� ��3��׀����8si�g%�8�l��NԽ-��<�t�US�H��#E�&�B�����[�RJ���9�CJV��):�������d���	�b�K'�����zy c�Y3�X�ٰ��:I��KdrޝƬ�	V�,ק���WxJ����o{n.׆��O��	Ƶ=h��X�^r�mE�n�z2P�p�a�hk�=�2G)�˭)�x����a?��,��9&�JhН�Ͷ^%�MϮ��ޔ;}<�rMX��*qA���'�]z�G�[��Zs�b��+)����V1~���o@\�%�.ypl�@<@ �ozY	CH�,�U�Y��@쵞fV�RTu�� �-��Q�$�@��Tc��n��(T���r�����-c�d�+s�@��/�=�v��4��Z>�������J�VK1����KP<��d��嗫�0���i=߼�k,|;XsK��{�}��"�ʶf��<�xs����M92��I3
�?�)c��)�ي�Oň�"��t��$K̔Ӆ�f�G�~��c��8!�x��	�Y W�Qf�@^k��MOTф_��F�rKB�48��D?��]��z���N�-{�isDސ���*�\�%��D-=��^�(�5q�-d��ك��P��W�l�A�ݲ11(�="��n�=�#w��L��u{��Y-�o�x�F����OkW�T��ؑ���s�$����բ��0�����;6d�PL�K;'%Ѩ�:8B~����zݒ���P��6�f)�0g�rF3g����w�%K��.���M��N�����-�i{��ሹ���Q��J{�2��~$֓a!l����y�H{.��DjULū�!<5�.����?��L����z���� ����O��@]S���S�Z�d���r�nl�&ab�4���L/vpQVD�5=�=�DZ{l7�=��p/�BX�q�?�C�!Ia���/xd�Wɺ~~A�7ȏ��}��aq2�G�8�B�k��BS2���y���<uDc��dP�Q���2����>L?eBa,��4Y֣��^{�1��
�B��}�k5e>�LR�4ݢV�������:B50�qcѤ��y���{��q���N�Z ���!DO�ԧk�U��	@jL�\Q	�r�G�4����r���x|�a� �N����:b�}9V=#$X�b!�+�\V�`����_��Ig�%�	~�m%& �9�g���ϝ�<�� �qe��eT;ƥ�u�E���6mɤ����t�������v��F��kZ�;|$�Q�f/_�AS��w��B� �M
���*q�z���RMlo�~��u�?7�T{����@��'5���($3S6[}V6��9��\���M����Oduy�l���\�����%mW9�b�b�V!��\TPZ �eŇq��x�����DP�j�x�Ǝ�q�7`�ڋ�PL���G��� �<����Xe����~�����emA����M����_ǿE� K�M���K1+)��L��PvY�L�?�*�ʍWmQ}�e�u�޲@-��;m��ÜL��K�G4o�� 0qֶ>���g$b��b��~/�M��7���t���� ��}�Y�ų�v��m�q�]Ŭt�ظ^Զ��?\үm���o{����s�@�����R]���4�*I�d`FA��?EW�-�,6��522L{�9�~�Ozj�[��E�H,�xA��U+�<�ߥ���*>9�K��|��T�ޔ�+�O��6Zv�(6P��Q����L�S�����a~ڱާQ?��|�/(Z��@��M�������
BR_-9z3��2,&�����s�+y[mw:1y\'�mR��-Y��]�?i�]�9��!�H�sk�9����i�>�F��o[���V��YE�f!%n�@ț�=ߞ����ջ�[F."9��b��k�u�+F�����.��(��/��u^��]Еw��&&��&ɥ�"f�q�V�-S��uD�)�6t�@A���0�Rn&��gQZ�Ea&-f����M����Y;��W�#��5����m��\ ��Ѣ�9�(�=��Z�vl.�P����{��U�b�K�*G��a�o�����ӑ?"�5V� ���zm��=�±�ѸN�@
Qf�+*n�a����_�k(OZ���4����Db�kF�	hڷ�z�¡�K�<�~�uo��]v�+��c�ZR�H{!����EpI.��%�+ʦ��p��è�m6t\Pe:G��r�08�/���������R�EB�^��;���G���<0�m�B��Fޘ~~)�{�i�K�9�Q2b�&^��<��ږ�W�TBq)� ֿ�x��@��n�ď�-ϊ|��H"v �L����׳�M./[�_>hR���p���� 	ݝ��bz�E��Rl!e1�,�E����[n��5d��􉎒����S(�jθ��_M`~�]v"ِHw���\&k��hK�t���y��M��w��� �Uǲ�e�+>x����Ҁg���Y�$���ţ�u��\
%h����8�"�i���#z�29E�$�B.��R��Km�;�O� ��N1��c3ư"��8�׳��N���PO�5�>cw�yA�>��T�9�+��; ,E�U�xqps�.�]�[3��r����L�>z1����"��,�}R{^�&��kvN�I?��B�%���n=�e����?�����!$3�|!�x�˲S�<�Zj�<(�$�X� �8^E{�=7|@�邪֎��:��h���-[Ve�n�ڛ��ֺ�;M��W���j������K�TO�"�q\�MH������U���~�M��#f��K��d�-��_�p�b뿾ٕ�T�gc�ӕ�sm�=�cF�Ʀ��)fX_��$U�Z�M�F!�A�&*rlؕ�����|�qLٰ|�?�/��Ũ���@�{�HX5
_����R⃈i+��bO!��jn���OG���@q�ѵ����Vٸ��sD�Cl���E�Q���HEL�E�je\�Qw��5rԨ����d��i�WTb���.�Z�,���˥�)P5�c�A\ж����f�����z�	��&��b�}���<eM0[��*��1�vA��i@��m>�F̫���M��\�i- �q�J��)�0,��XF��wT$y}��k7�5�t3in�+��s�SNE�{�%�\���(�pa����-\E�)�Y�v؉2r"��G�J�����U�Ǖ���)¼2���]9�s�MX�.��J���OSYB�]
�a|C�Z��"� �[���%��ۘ��		��.9Bu+�1�:#����I��-���K�<�q	Gv�`eg=_E�C¨ԍf�*�W����*lK�ꗢ�ytfv4� T1(uԎ��Sc}�L6�2���ր���ڮ���`<I�-�a[<h7i*���ѐ��b�EM�.�2�|5��9FO2"��'ĳ�|�Zy�V��qc%M��ҟHQ˻�4�o���R��G������\f4ߘ1P��/�/p�y�q)�Og��aר�O�F�ʝ]�^N�<�r���fA8��g��UQ���xw5��z��N0Q]"��(���	��0<�dE|�,���� [s/�л�t�c�Ȇ�n �ԙoQ1��1���a	
y�Շj�pi%�l3%��,}<z|"�yڌ�p\�.�9�x�Op���֘=][^)��ƌt��C�����?/QHĥ$񆢟eB�XH���qaN<m譵c2)ny�*Pe#b��ײ��^5�AY15Lw}�a����I��� �%�,:�|rt����:�Cy�F����?b�IՎ2�]&F��p���X��Fc�S���;��%+kU��@���j��\d�G4N�.�@��W���	:֭D+&D���lD��]��{�I^��T_������'Z^px���*:��QBjn<K0ܥ���Z�-���g0%��ı�K�{��{Q_���S���,G�o>sY��ӛ�(���ֶUt����z�m���u�3(�~�1\��:W帺[e���}����j��N�p�J�2�)y<I޷p�H7�����H��$�᪠��2k�H��-k����}����^�욏o6��|�UB�1��.���:�}}W|�i��� �_�3�	��PÅ0�Ă��t��� m���!N6&���/�%��c͐1�����_d�o����nU��!%�s�,v:6��K潸�i�ȳ)'~Ȋ��$��[p@���>�zh����ǋ1�ז#��z��[��w����`EUa�-��ppt�Fa	�"�����Rѷ���20����v��r"�8��ֽ:�0|��Ѭ��i���i�U��D��b��e�K0VcZP�u�+K��Nn�4�)���柹sB�;;7Q1v`&b��(�����"\�u)&���9�|l&����(��`_k�s�1'CP���e�Sҟ��Gd�JL�$��b�"dt{:�8P"��T����Me���Ɲ�o��2{�H����e��*I������$;#&���{���B�F����P ����:��� S��Ϊ ��P�l���BrA�뗸���ȗ����=ؔ�І�YA��r ����~]�����8e�5#��� I��7�!�����~ُ�t�7��Y}��3�p$(A�l�vY�g�$�J~Oe&��:��5���0��G?]�T��b�O|���HxM>٤ )�w�,1_���S�ͺ�,��q��KA�gN�NPU��-���X�I��h\�i���g!F������R&qFՙ�k��Y����ؔ���T��G�)�aM�������n������<,:�e�|�Z���:�٬�r9X�ajV��n�jXﰓt�'�sT~+`v�������Y�	�XEZC����r4���	x�n�!���=�uD��
(��\�X��ӄ��h�Yj��~�j������Ԣ����F~����ڶ44u�w��r8^��l �iɗ�0��3��|�ġ����S+̗ ���H2�Dn候z�,��]l�'lx������Ms�iې!1+��{�,5S� �V��pGH~�\@��F�"�48��K}L�S�|��o�!��f�6W�x骷C�H[�Ak(�~GMi=Ɔ�87Ā��=��bwH!M�^	�m� A�M���zX��.jS��7�����Ĝ�?�8l���1�e�do���N�\aV�xh͆RBZڠ� ��+�U��7KRb��[]��9̭���$��ތ�ԣr
��΃0��	/2@�M�V&�ye �*�naDPM��;u��K�|����P��ؚy�;�<I#s ���{hW�+��LU�����f)��%����*?�j���s�����5^�3�o]�n�N�V�������{1���V��q	��\G��5E^���}Jv`Q-/_�Bᓋs��UG��_��P��&���w>5I1�k0݁̈́��3'K��[̕������lp&�Bs�4w.1_w^��.r7s�Ō�n���∨� Pf%�ۿ��ZO�������=�Х���xAwM��d-�^�=E+��zS5f�G��/q�d�YAJ��CD�&�%خ5��K��I�O>Z`���l���ޗV�b֯l�i�]6���gjaѹ�aA>N�K-�cHL)�:�-r�w�c ��1x$���M�Yp�<)!7�G ЌK�o:}V�A��?i�I�Ǐl��e������z}"�XZ�=�Å;d��y���jơ5�
z�H�]�d��%$�C�F�q#����EZzl0��^xĂ��LF�+b���,OEYGhM�}���i��a�!x@4�S�ݵ]�m���h����a�7E�HѸ��P�t�y�|rj	V]�I�����2Cl%�1�V�7�np"��=zip�[2ѽ��N��|ɟ'4�#a�?����j��3�	����./����HI3�xbAZ�E���2�A��2)SE�(t}c�VU�#�V`"<��K�<��pTA���	��a��wA~d�W��f�:%�a��z�F|�y  ي-�; q�}����D�-!�tP��7�A=�?�A�+�����3c��A�@��&F7x��3!a`ղw̖���#�����s�q�)�~=Cd�#��y3r�|�h���E�,�D���}{6���~�C�t�Rc7v����5��n�h��a\J-9����+:Pmsβk��{J@[0���jK=4���Qࠈ; �S �_�GF�d�۹j�G�$�'(U���.-��`z@��~�7�)|�Y��s�����o�
К;W���v�g���;���;�i�pi!-!�쟪!7n N�8{��8#	���Ka�_��x���g��3Hm�?Pd������=^c��q�9���j ��=�T�^:�wl(Vi��)�#��@嶥@���掏�G��C`�n���w�|��]����rv	�SÐY0XԳ8+�i	�|�� ֘��[�y+�߹)��H+���hw9���~%m�� 
֝�a
��@&�,?%m�2�,�:�+�7J{7�^�`����+�%��z�X� $K�vg0��k�u3��Lv�-wX�y�E�� ef�x�=
3��oI��i��s�*PܹBրb<�:�RZV�;3���WN�j��P`���n�R
v�����q!���$�C�Yݒt�\�x{�N=hi��%��K�-�#�YX��"�$=�uwl�Y�����_���O4��-��!��7�
kh�65��ըB�l�5���@ p~$
����>E2� N,;�Q
P�l�ЭVt����m`:o�wC�5Xe^@`�K���c��g��:V���lnT��?�x0Q͐��k:In�g�{��
5�`�n�`6E>b"M8�s�O)i������s�=WU�^JB{��V���6f�/���@�J�j���V7�|� #�v��FV�Pn
�T�����FY
�&(�}���	�Sjf��Mm���(e��c������a}7��o��ȮCD�C��ݓSJ�V��<��#�������-��@�y�>�Wگخ�S��%-gv<��aƍ"���[`�99i%}]���5g�!��e;����q��*~�	�m�����A�1a�ذ�5f�F_�oe7*���H�%����`0]�ܾ�8�ul͈˦��M��r���rڍ���"�R]�<�C1*�$G2�,�O�꼘z��s";1�+{_���^U��$~ 67Do�JjOR��B�G,���sE�i#,���Z�V��k��̢E%�n���g��.0��"ϙ$.fEd�؋���SĤ�����Yƻ��e��%��bU�/�8/����+P�V�8��NO���d�2/��h�� �x�P��o��$�٢���_��wc<��`��"J����+�s;�9�k����c��dv�u��2���4���n��f3�4��vg����ޠH�{���4�J�!ft��Ǖ�Ad��K���"`$8�c~?��rͶ���.��Í�H�ˇ F�k9�;0���A�0%�"FFX"F�=sHz2�\����2ܾ�2�C�ăU�q��s����m|ɱ�m����X�W���\e{���j���Q�ƛBs�1Ae ,2d�1�7��t �H��ҴJ�P�W���X��z��Õ�b5�*�H+�_ 4�t��ܫ�;an��	\{w�!�M����ς��rqz�l�������-���L'�>eC�ыކ��P^��c���Oub����� �NƸ��u����qpF/��%m��YҤ 
�Y�Q�݅�t(���?f�O*W��K><�T�aB�ò1�)#� �*@x���H��n %�����:D�F�N�~�x<4;�s�U�>�ω�f�%���ఒ���R�wr��
�07$�x�+�𙣖�����2�&F}c���(����a{�$mTٖ.r#5�&����2��Ŋ@?�|��\�q� Z�&�nܧ�xn �&7<�l�u`���]�rvDp"q�<Y?�6\�/� !g��}���Y;�K"Ei���;�ɉ�0��i%��yk=W���ȓ=~�ܲX��9�|D!/(,���e��vz���!t�6�f&��5� ڈs�+>��d:l�"ъËr&��ݟS]�%��I���8�?ӭW�H���v���$c?E���K����3��m���i�UR�(z!G鋟Ϫ�&G�ߪ
?�1~G�
�9�e�V1���c��^U�-��'��\��x���B���ĸc���j�kHX���bG����D���4�(�D�XQ���	�3��f�4�+7F��eq�c΂�7���� �=��P:8�ōLf��)��#	=U�P(+ӹ:v&}��l�&�-_'ѭ�!a)-�p^F�N$T%pՓ�������Pc�t�Q���N�]cB��Z�I]Q+#�V?�8�c�$�-��>��hw�G	�}��;�*O6����k��[G���.�����H�'/�FE�4���ᬞǸo�0�49�&�zP�M\�������߅��Q��s���|f�9��"~�Pj7�+ob<<��=�ƁZ��Cjj���S��aĠ� �R`�-�f G�a}��[^ZO��Q*�Q�l+e�H�b{b�)�T��pպ<`�\x�x��At��M�=���,��B�r�0���L���t���d��Y���oo���񷲃�9u��w%��O+�9����8�����h��p +���{��֐�z�ixˉ9a����d�C���l{?:���,$?����-͝4FN�B��X�H�Y^�+���?�Vљ�H@��q-X��a"ə#�޾�ſ �%�t�4�a����E牟0���Խz2��D�w\�s��Fvp�d�^���z�5?�'Z?�u��L� �}eb�@%I�\�E���^��޴ԫ� Hq�}Ѹ�Z5�]UWg@W!�:�H c�(�.�`��)f������!:�]�������?=Ԁ\��U������"(�MB$c��SPe4��\:y�B����~��4�3�����i��+Ӯ�;��+GR���RbY~	`q>����	��ڂ��G�(�K���Դ.�Թ���(
�F�e�ʮ����&jv�|뤞2<]k��p�L��a#^7�ߨ���P� ZV�ۯD��^j{��ta"���2u;.�d�i8��0�0U�'IIд.���D�TO�qX?u�v�ԛ��4`
�ގ�zΞQ����e�W��'��X:|\c�#t�I�x��aDr�1x\p�*|G��;����qX�TCƎ����k-�޾<!`��%�S��	����
f�y���+�F������l�=Oi/ϼ٪�� �;��QIsT���0X�|Ӧ*��RQ�����?�L�ݻN��}n&�S���Y$���.�줼D����j�ߛ�U&�V�ۣ����Sq��B��b:��
*��\Н7�'I�{��6[X��*�VS���[�\��u��jw֨�d�bQ�Io���
�d��˥���T㟋�z[V�Ӹ�n��|�~��E�eg�^�%��3o����Vh�џфM|Ro�����8bG��?g�UE4>cA�{h�M�D�	?f0�pu��t��h��Q�{��i�T�?U���r{A��g�H�f�f:��i�0i��h\�2ʪ�>������4PBc�Y�r�W0���?�9�6聗��&���1�vV=��P����b��u����V5��?����Q)pɪ���1�!O|��8gRi6l�i��LK��k�r�t��F�QEPkļʻ�?�\p���{�6�m���y;b	�H��=kQ��j|�ƾ�Љ�10�wKy�'�\ Q�E�p��2�*џ�4T����/�[�v�؈�
�b�t\���%��?@�f���`
����y��a�TCm5�rn��[��ڡ�������G���2�A���=KRf͒��ml�/YYpZ|�M5i�6����tTa��L�04�ܙֳ7ԪX�[
ߠ���*,K����i�>���z����JI:�����+�(�W�I��u?!�� �^�:vOVm����α����ެ}�Vf�B�]O�oN��8��ls&DF�(���5V�����j�I�D�5�^Z%�z#ϛ��Ą>Lt8]����u�>�)|�콜y� px��	A���
V�DO�}]%���mZ�B�<�4�F�݀s�W� ,9&�Z��!"½_��!AŴo|
I?H-,˟�A��z��g����P.R%&�R�ˬW��Q�z�����w�g�(gZ�g�~��5T�=d'��hs-е��F<)�7�g�z�S�wnQ:�Њ�p���k���j�tt&	���F�qH��,�(�{n+m����D�P�H�x�E�i�����^\�<���T�q>׽(4wOڿ}y��Mg�� �H*iِ�^ew��g�^�OE�&��Oh!��]��g�b��9+f.�:�1G�{a1"z���z��ri���o� �O����v �#C�9r����D"��#(g瀸�LT�`:/�����
/��l>�L�[�2��;�h��,��]A� '�.w�-)�:�(����A�Z֛�	���D�-/�P����>��l2�)mbh���Uf���V����5W��(����}��wTd
������c�@7��:��%�%_��5��K�5YгQ���2^�Y�\���B��A�
����8����t���\��}�Yϕ��uL�J���(z��Saobz2l3r�R(q���E�j֔<�D���G�����k*
�A(�1���J�H{��᭏4��'#�~�����@�?��"�<�NMB���q�v.��.A"F�c�ь��X�J��`d(-��x�]F���b�!�� ��z¦��F#���n,��B0a<����߁�7���M};+��N3ܘR��I���b��Q
C���?��$c�g���H���e��q��WȲI9{�]���'Ζ�	��6cK��O��<����'��o���WӍ�W��t"`�a�э%��H)�i;}�����U�y�^��K��������R�^�(��r΀���ww_W�ht�_�bX��O8�$I���kv�(IT�W[}�b��_޾t��&=�}�����\�M��>�%������z!����2�l��S��e��O��@wh4R�U����
�x�B�#Ύ{���l� ��?�1���Ut&�F�Ц�� �k�D7��b"wa=568P���K,<@�SW�D�� t;�C�x0[�\��X�~g'�멥{�nE�0�8f�Dw,jp��S�7ZӶv�ۉV��֜HU5��b�3X�֮f;�����gC��a�'F�H��.,����G\��A��X�Oܑ�8�{�A�,�%���V��,!5�cc�&D�b�6�8�vt�rX{Ѡ[gV��^.���z���<ZP5Z{L�)�p�f,���T@��.�?�%�WO[q��w�j8�X��IA�"o���@W�'K�����}&���Į�*^�.
U�I���D��!j8.*�g?ƓL��˘�g3�R��,���M��v���֩�c�R��
(<N���~!??�Q�	O�z��'�s��M*@K�,`H89<5Q;�^D��[I���>��C�W��=�LH����1Y�ca�T���~�|",i˽�B��X{���g�؈K��{��0'�٭����C�����o男���[=e����X�\�L�'��N��84�忘 � �j�l����j�ҲK��;+R�ׂ|H��J;���n	�>�����Y���+D>*����	�eoJ:�Z�������6?��� @�����G����#� ʲ\�d������"��0�Q��ϔ�$��c&�r�l�.�J��U�*�Լ�ە9��X��t�����0N\�x�}����"�c+g|�R!{.��D�[s=����3�#���(	��O�-�J(��FΊ�B.y[������a�gC&3D����(��H�L�ۈ�!��Л��D�����������4��N���~���O`�N����������/��eU\�j6Z	�~H�������yk���Z)S������'@)҇b���sQ�VJL���o%�G�z�G��qb�� {�y<���w,Ώ9Mέ�:E�\���{�7��}�:I+�+��r��6�l�H�����eom�=��YEe�i��	dA��:���%x'hT� �N��%�3?\V?�y� �2R��0�chә�Ӳ~|���QS�K�ۉ�5��'�b�o$UI���|h@�#.3SPX|��$������F��n���:�����E)�D(̮��[���t�Fʣ3�fpEzI���t=3���cB �=���?�������_���`p�;�k�	�A��n,�G�,0���+��AC�E�9(5DW�o^l�PaD?���R<�bTq�vg���tO�;Qfl8����N5�r��=�p14��'���sˇ`�0T���s�Ip�ә���2� �[`_�8+	i�!�9��SG��@����d��n��l��%�bg"Ƚ+�ѫJ�y_(��Wq� R e�5�\�x����b���ԅw���*��+�rhj�_��m����m7嵠Ϗq��,�Ꮙ=}��#n�8�k���PG%Мn�P����|�v�J��`�a�Rn�����c�<����v��<��t�]�û�3�z!��]\f��帅l���MαC1qX)�S|��d�kM���IaB� �7:�񋆞d5W.�Xx[bk�N�jIƕY���ݾd?�� �C�yAZˋV	O/χ�:�6>[��R�����c,c]݊��a���8�����_�U�޾���Jw�Þ��khf�E ���=ma��5\�/�gҤ΅R(!T0B�DK�
�[�"��C$����e���]��"����- Z�S!�m+y� �{�㑘Y��w��'������� 0�����4�^˳FP�騮iD�-Ky�w�[�}�찑܊[��]M��)����l�{ι�/��u���M��7�ɬ����Bn�ӽM���=T�&�|SO	�dCd�+y��m,���g~������PQ7�����Ҟ����%F*OW�x�Ë>��wx�T�@�[Ԧ����'���$H�u>J�=y�-#pkS�;�e����\Wuf��Yr�84<���6�d�qȒ��4W���&D5D*������^� |$i�Oyw�Kg_��v��en���E��\$<RU��ͽ�L�{`���U�I�6����f��հ�ũӾ+�l�j*��~���O�[zWkA����Ѫ�Iu�f�9�:}��4r��yfp���#?_�']�"s7��A C8�`��l��d5���@��_0��+��Fy��m�Q>9}��1�]������DQӷ9�f**Ֆ�*W[wVط�ְ��<�;�c=�%{mRehjWa��E�>�Q�1i��Z����*C��{^�f�{�N�����ʡ`<W���|(�ɷ�Db�׬=oC�x*Ŀ�������Ő��IÈ��l%+�!��S'꭭q8o��$X��0��ﲨ�o�U��@�E��*�W�* �1���'T���f��^E���M>B�w�΢y`"��S�vGE·������n��*�&	6����������E��Tg�2%y�*!���E�n����Rq��T����w�����QQ��P���ң�S�]5����j,8��=g,�JZ�TA-����Y.�n�.Zcb����#�K> U�)�������>��y簑)�I�mg��b�}H����N�ӳӛ��bR�葙Ġ�f�þ<d��
L�-���=p�_8Mc��5�����^E���&m��(hL��73�T����ݾ7u���BC?��v�Ɋ��3�?vo��v=�N�w�Sy GI�!_S�n�=:�#���oŬK�(������B�4��:�m0DQ��	�:�л���t]�c���O���`����^R�,���o@W�^�`�1P�����B��`~�A���~E�[F��������G��ش+ds���a��-��TL��l����Y�_!��/
D^�f����_6,Mtn�i�/��hۨ�
�^��9��4g9Ov���͐A�Xe��"K�:+c�ȶ,��@�F�5���yH3Y�KC��W/5��Sv!%��1���j<�-�8������Bo.^x�A�H���O@�=��kTG�ybHɴS��C+$�4ԮB{?4��M`���lM�S�N �����H{��I^�0�䐦Z�s��[���Eh�h̲:h.���%