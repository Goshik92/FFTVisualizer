��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��?x�?��Q��'��Ot�뙿�l��Qu����*��4O��P*�<����s))�(����0�)D���a/�J��Q�X~�a���Pa�OF���,�9��&~�/`��*V�~	�i	JJB	������n���X�w�Չ�����De3=%!�z=8�cڌ�ibq|��>�^����W��L߈x�_��G�4	�8'o܈�ߕ����@-�EӸkJ̣�w�d*2�\_=��Y(�MR��������*�K��b!U	�a��yw����Wd�G�H�6Y��O�,��I$�5�=x�F�(X3+���b��`����WO�Q��a���"�U�rX$�Fp�#A��J�<*���6ZZko��ĭ�w��x{mɤe�6��T�cx�4����K�U[�`X(�@'݉?�-���_ת�(�{����p}�'�鞞���,'`;�@o��0I+"�]����;��N*���Y�F(�X��a�������p8��
%-	�S^��[�`�q1����Y�LB���������G���Sj�����HeC�v�R�){�����RC;��M��-��|��˽*��yD�� �,��,�/���QJoO�jwu�+�����-�*�5�(F-�Q6�<�޵sI���v?,myj�v�7H]T�P;\M����v��j93�����ԙ��o4��a��iKO~攞7gI'��C��5�M�;^zP��!��z=��+z�o�p�K�qr���*4�A�n�_Q���{�9�H����ߑBA����3F�>�m�`Is�cUZD�v�����Ny�b9�:�6���8�5ӽ���r�s��<>q	��<E��Ɏ;_ǋ�XI�8���z 3	X�"(�U�����0ub�,���u���Я�2��,[�uR�7l9��ցF\)/�󯎤6�T��?�@�A�����`�����7�Z�J:�u^9"Q���:���n"��8��v�GR�	n,���S��>LPebT�:&��VO+?6w�j�����:�G�z�ilj�}=Y?L�z�����"�<ha�<|��z�=j����PY���.R�8T�,o{�g����?;�5A����Ͻ%t�lQ�E�c l+�{�P�@��:����T��p�;ϖ��du��Jd�J�H�����HB�Sw[�������?�㮮���������=�'e�f6����j�X�na҈q�$/[���T|��+�\��c����Y�� �RW���S=�X����S��A�*��Ɉł�(��`�9MV����c;"���CUd>��g`�+u�n.]��a��y���l���Yф3F�
)�S؞����l�`��%�@ �WUΑ�{VfI�J�<��=�t�	Q��6��q�:�<O�ߏ�Xl��9rhjr^Oy
2A��7��2A�@���v	Tc����K8�4��LK��ZlG7��ٻ�Ex�Co.(ҵ�w)����"]_<��ew�6mA�5�}�y(?���Z����|���UҜz��R��V��q�t���y�I�N"e3>�Q�ap�1���r�����|Z4I�b��� �����%���f	�2�B�RV�ъ%�cd_�ї��QvL���~f�|�М/��T6�;*�A뀏�����g�F�&{늵,�E��h\�0�(m�z��1T�0��Ϧ���2u�)V �I�)�l��Q��oQE[��9�,�N��+a'�7Sf�/M<.�����L���Vn�P�!�5�����H��̪a��5�ծ�sM��>wd���>�H`��T<r��/���#�ċ�8 ��n�����Ta{�L����BB���	��d������P�%��,3�%�ئ�%�m�n��q�n:SXw�S/,�]��@��<SH��b<�f;{��%|�t���(��c2�ɗ��VU��������v5l�<4.�\����c�q�j8�Ϲ}Kyid wS�p^o�@xM�WuR�u��GK����^�Zc���A�E�$@[�����>_8���"��胲�5槀�%��f�-d( �E�x�+m+s��%�ZQ�C���"y���?@�VM9}�8��cB3=:~���uf'�K�K��.A�A��H\�zv%�R����oI��V&V��g?�ݻ��{�i)0 �������ʼ�<��!�7����p�18���I�m2���l��|L��&�R-�����D�����?��^IRx��M��gZb�d�ԅs� �	b`���Z%����A�S~��{�XT�+"	�l�s�"0���	���?�Ċ��Z�C�e��ΩO�'}���q�� �Ot��/���ϻy��}F��t��#B�
��W9.>F�Cd(0ɥq9|���Oe�	�o���[��b����<�|��5�DJ���|���Wm��� e'���lq[�R�����������c�������Fӿ����8+�P����G��q«GW�ŵ�GdL���7S2�G|�Iw*���LR�����f=#���%f��]�IS]�zl��ʞ<������Y2[��ڳ�MR����OH�\��= �����XXo�[�u�D~�h��]S)�0�x9p��7�`Z�RuBj[�u�m����}��D����I��eot�c�Z>ۤ �u������R�� �'��)�L�r� �B1��5�ǐ�Գn��ӗb���^Ő��q&��X�V��hꎄ�l���9[�W �>��$q
���MZ���d���5���:�@����{P���2Ǩ�WG�b��C�������7��8�WeF���9�L��pHJ�H�'�	J���_l��-��{�2���G_o>�^#���kNg���_(�Z�����\z|���~�g����^T	i`��/��)X�t@���	��#x���Z3�t>��f��*f5���U�̙���/"�<��S������x���~06冃���-�oκ�/M�zHXg�irakNd���a�`'~4�EYZ6���j�#ʜ\W��3ݗ.S���>*J$�B4)�@�IK^4dBA��~���⸒?[��)�|��͓'����b�@�7��B
K���'[4A�.��U��q_m�� ���V9��1jm0��']ls��������K��.s����>��I`����a0k�S%�@a���6b���X�w����]3��<Z"�����ʆX���ť�{�92a�X�����Y��|@rS�q���&L���L�����	�yf@ ���>d~�:U��8S)}b"Br�H�p�S��@��������eY6ڛ\�q9��H��/�(w"��R� P[��[N����d?�3V����Z�G�X_1$K��-16�DĽ2��k����"q�碾�̡چ���{K � o�,Ϛ�y}�,-�!��`��ޭ��?y��L��^Z�r�!l���f�ٴ2[��Է3W�SE�@�Ybǝ`R�Q��5�p$���fC1�%�O.�Mi�oɎΨ�0n�cJ�:�C|�JG'bբ���rn6�\	�H�Xܗuo�*������aC�Z�ӲC%��I�A�"5T)��LW���~�_���"���Jχ�1�L��m�F�|��v��l�D��;���׳8=��-#W�,�]m�G Xc��-3x�c��_��޸X�r.��t -m�S��s�**���(��˂E�6�?� |�#�~��0:���%m�+E/��fWD�h�|���Z Q'���C����ś��
�ᇢp��>�AΎ5�����V����Zu3v��+;��3�w�.�{��߷//�Ao�u�T��2�;�2rS^��~N�����E���5v�q	-�<�ABt�}�k�J�;1��y��&$r���/��V�����3r�F�ߒ4|�:n��҈r��RgD�(}3GA'�pPI��Q�T��*�0� �*DOX�������;�G�ƍ���)Y@9�������$�oP�Ȼ|se��N����x�.Q��3$���������T��/�A,2'��X,]����%bAP�o<�3P��IJێ��ԡ}�_WF}<$��+��7rh;�@������2^_�$E��J��"e쵲!�i"3�$s�{YN�Õ!F��_���ֶ�Sq� ?I���.�l��,�S�wq��O:���);��/�c�;��w�b�Ĥh��02��H�-�`���������,j8�|�βг�򾶕%?���o)^ƺaM��5F;���ZTuM�rh��J�,���lG�z�#uV���݉x�Y���!���+��8�0�|(��V��I7���>���b{ձr�B6�K�# ��
l��d�$4>C�x�	�PK�mGY<U+�*��՞�"�>u�**�<t��ʌؾ�)5���
�|��\
�ɺ��7�[yV/�A��N�#'{� ����aM��� >x�ˤ���!�=�H��ߴ*7A@�}lxJ���giG�%�D�:z8F�`������	�(�vL����1���S���&�Ȉ��X��Z~lJdF#Uv��e�Q��3��ꩬ�LAG���҂)?�l��`�u5�-��u�"��}���Og^�7/����)��(E-Om� �F@HjK�f�/2�sBL/x>�|T*�F��e���C56[���ء� +uհo�qڗ���C(��~�e�!�&�#=���{�oP�K0�_o:��;�3.RX�
���w��3 ��6ܬ\?�&m�s�W`�|���l�35Z�o�p����B}�!ÖyƦ�5��^��	��E���7Uu�J0�\Q�u�b�a� �6R�����kR�m1�h G��"��J�z�ԐʈS���ߡ�.o�ģξ� v���$�bہ\߼ao��ϩ��<���d.�H�u�G����I�dI�<�Vj��ߞ��&Ub�N����c��5�xK)%E�)�J"��RQ1�E�]w�S^�f��O�|D��Y^�Rd�Ri�o�ҕ��Q��k��o�jye��=��\{'�v�œ`�%�|�7xf�]�v��t�Գ��KY���6����#UV;���/�o#N����ߓ� ��.+�''A�%e����<T���}�X@���ei�L��D8�Y�:�I�7ig�B/F��Sm���Sv�L�y"�Dv��h(�o�K2,��	O��!^7�Rٽ=OIv`����B�}����c�ME��Re:7�i����;��/�|bcNha�
8�p�26c��J�K*&����XМ��9 �G)����g�z4��\�Hˠ ?2�w�
�i=<H4ԓ�0�O\������/k��߮�(U��II���~�\��D�j���#�RP5=5v���cNvyn�E@
S�-�� gTC��59u4+$]4DLZd^6]���}���r=�Ue���Y}�$��{�y�C���!(+#U�Ն����{����kN����x�6U���Ia�!��5���kf�4�e�<@�y;9yF�U@��B�s���?���\��U�I����T�>���˞R'�_̇��kx��P���򝃁jZ�/�;��k:8���dgd�4�w��A�_���/*��	��W��Mw�$$���r�#�X�����J�� g�ᎌ���?k݉4Y"B�|�.�F��eB,��FqY���Zad?L}��ٹ�&�a�r9����@�Qv{Q|/4��7���AKE�pښ�i����M�`<�<a���̘���3F�	�R�ʆ���絽��I���g�`�D T�q̃�ҡP#@���s�	�}���;+-
��J�e]J��R��AZ��xg>ՉZ̪M	�6�*��3j��]`�ےn������p��^0B�����C]�j�T�(r��s%7������Y�#��(�ڹP�p|5��-��$��lEDbV6�r.�b{���5���t�{���(C]�����O2��WP�v�b䯝�wZ����ZT�5
;_"�3�G>ƳP@9�ʟ��Q�">zD�#��$��oؘU�*�Ƶ̤��� ����'E>�j�8
�&WJ�Po�m��tp�_.������i@~�.�����ږ����/��܇��`���Ĳb)����Q����v�.Ky�(!Bq٪����쟟��G�����d�W8_�8\�������;�'��N�:H��(�x�~���Hh��$����!���
Sm��N�I�6�0 �]Ή<nxu���}@T�+?|���*[�"l�~��yHFZ�}�F,��ͳM���6��g�S����Y�Ga�R��3E}촫~�7�d�VBYŭbۗŰ�9d�ߣ�P�CV�3=���xH�B��sJR��Ǔ�M,M4q6���UDl�ąf���W�H�ѽ�m���}��x�P��ǙU�$ǜ�.���x�?�߸�C�q[�G��
�2݂�W�G=VQ�q��k��Z��MK
��jp�8��Ȑ@�DwL��������B2R�x�v3GeE��Vg@��ף�κ�(T'Z��ߢ#���B��aJ�H��7zܳ�o�(���ҧ��{n��&�Z����e�=�j��<��.��E{�_���,�%Q��i�?={�Z�d�qj_P#���騒Wj�=�(�˩	�v��@���뵄TPC��~S�4����NƁ
x@$���=������g��Y�i+�<�Y���J^wxR�/����^`"�8�g�̽I����!~���T��y�#��}�?���s��v��]�^ŗ��bo��R�'AG@r��z�Y��Y�6�Te��X�]�՗�yw����'.��[���`܈��B����]p�e*&}��|+��lÐ��Q���[��7Ǫ%r%��T�2�29��+�\���9`�wk���]Ō5ؕ�`��#�6�A�]�H�C���ɒ�B��1p�RrK@�S��X�@f�c�h�Q���X�>t�$��*Cy:����b4�:u�ݫb��]�H�6֬rUuiR�����Ҟ2;t�9F�Uol���^�72~!�۬L_j��D;mH���F�+]���r�i�=�98��[�Iş���l+�M{pTc��w���J0y����D�|��4���	�m�:��`�.�6M�E���	"NpX���|ڇr�G��r��}�X:�u{��	�V���u��U~G�m
�P����N�K
��0�� 7w��a��f^
]��[³�?Z��^���i�H�N.����>t�T�m���Kx�2��i�G�5/t��X#`�t�i�� �����θ�fT�Jq,ś�H��!qJ�����X�iEbrti�×[T��\�����m~1[׮n�{�ʕ�b�O�����np��t�#̙u��Z�����
i���o���>�wƔ�ݐH�P+���7yx�=�;���N�)�@.���\{�0��2�ԇw��Pa�!z�(�OLf+�RӠsB�y��8rrc�1��Ӎ=z�x�=��ɥ�0或��.dpR�Mgr���>��ڋd)vKw�g�]`�_��]݌�)B��;�B�i+������Q��,�ANo#��j�����OL�x{A�c�-�NQ��%�����=5"���C�H�R9��\�|.,��AJlP�I�p�R�m7���=��!�{�:�W�@8��W������]g���x�b$;՛�)�ST�ힵE���W��^��Z�r����Rr�P�����5�rI�����-��h�^T|��xZqx-N𿏠[��6����2�#'�id-���@׈��	�am���ޘ�Ja���،�{��z{���Mo�CJEaKhm�hoؚ�0߸xF��ճZƷ��_qՓVKݾd�<M�9<ţ}���]PZ��<*���Zdp_Ӯ"��w0`	x2}� ���Hf��b� ��F�d����^,Uw�@�� u���23)H�>��b��G1������w����UZ���j�i�ܒ~˳R�V�@1{�͑-O�j��a�����D��j�������l��[�ԂN6��(����Hg�I��E��)с�����3K���-�@����"�[���:��:oe?qbϚ��܈��k��7�N���R�Ҥ��y�.�A�V.��<��>��?saS����5�=��*|\#v��Ò����� ��E��H8>�-hO>�[CX�7������ Ț�X��l�����n��J5c��"�4w����*l�=�E�����P8�Fw��u?j[���㸨%�m�3��QyI9(b�s�����<��	Ҋ� TxB��Q�� �O��ц �BeKF��/ܼ��X����>��I���2J�lv�ECQ�X^h�_��1#j���V�4��
�'���9�d�b5q��Y������O�E��e�/$d�D�!�6_���2���̞��9ú>Ǥ�������v}���\\^F���ﳄ~*�M�4��w(�e�7��Gؐ�Y8Q0Z�)y,2�`(�\�V�5U$����(���{%V4�����
9��r��"�,��迋�*0Y��&�@A�v�/.���/͵��k��Nc}83-}�U���`_	����M��.�)VgR@XQ���P�F�-|b��%�Gjҙ@[]>wo���jw��K@��|v}�}Qv�{R�ۗU�&�H�0zڻ�5|�(hS��<3�e
x��B����;�+'�x|��\Fe��v�d���]���Q�Vn�̤��g��Ο�4R�"Y�Ro"vh�_���Ef�G�����4��)���m�֓��La��i N�����mN�XL��4>c�ո"^bH��6�}!2a���M	����0ۚ�9Q�d��
/���}澕D���e�ɱG��N[P�{��]���	�0���}z��5QcD> �V��S���?�p��rr�1�����1~t��*�HD�]�
�2�s碯���;i5E��m8r���v&��j�zF�I�3�+��S\+t΋����V�'5���z�P����/�06��oQ�f2f�;C�Tޕ����L�����y���I~�]��B�	 R����CM����%�]e+7�X���:��/@ê����B�;W����/��5p����R�^#i$l���}�Ե��"x�_G^H�y`H@-X6���e3R�Oԙ:���٦�w��(��!-����v�Ŗ�d�>]��}0_�-ݸ\��6@w�1K�:�(�]�D'�V�\���O��6;��.����/jw�Pk~K�.�Uaq
�_�/77��G���a+W��7�d؛��U��8ie�Z2fG�ȗ���^����w�R����`�_��#H0O��D���I����H��"d5�B�|���Z�1��ȩpv�*hG�`�����"}�i��Ƭ��.^�7���5~I�A��Kb�C�~���`��v!�B���5�U������5��A��B���q���ë��S'���O��6��v9[Ј��w6VQT���烿gr� u���t^��Z&]([���N�X�<��ٯe���X�G�x~}�5-)D֬:��0�#ʮ��n��>�x��j��	 ���a�[�Ĝ�F��м00���w2}weP4����Eȡ�k��[���j1����9�z�>cW �[v\7ٷ���d�5���7I�����_7�4Y��9_���.(�B��3(9��.l�Ր�������M��^�ڈ��O��'Q��������{��p�[�I�F�Ii�8R���L���U�[p�ZK7�z���a�0�>f]?��M��PkV�2��4�w�!%6�l�v`i�`&�BxkN�\��P��d�ңފ�Y������*W���H�W�__x��˹Ѻj����LXCK� <a�|�����L�	���T�q8�8E�7�֠�s���2[?/y�g��[�((�����ҋ��ʤ�W�}�C}Ɍu��OK��G[T� $�Y�N9�iוSN�]H�-{6oϝu?L����/�&"n�~���!jR�����p��[���A�w�[Z�xe��кR��6�v<�0�j�:z?�ƶR����"��o� DG�ȡ�m�L(L��Z�̇7OC:[`n['�(=�,��{�uk�w�ͯ @�+ktC��΅�"!.�ON��q(�y�H˧c|�����ׂy3W�S:���n�j���5��A�DT���s0
v��	I���4�3�XūZ�{$jgs��%Tncw�{���E����C�t4%�����eS��8p��^x|��UDP��ئ���C�09;uK��Nt��XD�a�9]�
E���� �CD�l	�r�@��tIG���h*(t�(�z" W�ց�1�4xR��͟c��C㐯��q>��MqO�հl�Y~��z^�Y�M�P|��G��^Nc;�쓒�R
,�1��L�D�O��l\Z
+jX�7�,T���e("4��������z�)i��5��m�(��۔��"�����غ!����B���|GS&����?����p���U���FQ��M���Wv�#��x*��?�H`��Z����~~�<�A��\˸�������|�B��QI���!��4j��VI��X�p�w̱�Z��U��$r��4t�
G/��7�p���R�X&4@�a�f�p�,�og���B)�v:�G� ���{�4��|)Y9���GUVG,�UB�my��#X�g��+�����ō+^�1b�=��F:��YT��f(�¦���8.�4^�$��ȑp&0YSTf�V?�a}��I�h4�����*GxI�ob`D�,f�i{H�賶��S�.�;(S)4��}�����K�H�W��g`�ϼ��n����o
����k��&��q#��c̋.��ռr��=}h�N��rX��</R:c�t녥�f��i�K����3Z��Ʃ5u��Q�^��c>���F^��Xp��%*|!���������]D�aA��n����M4
e.��3�1d��s
���;:6׫���	��x�n̮aw'�3�>B<��>���k*ѷx�HwD�Y56a$�-2�EUߏ����d�	d4%��� ��|�v&�	��X��,�מ|qX�K$G̜�:�1ь\7�k����}���(� x_y7x�U����d/CX�	�����<twͤ�Ҥ�Df�b՝
f4��2�q$�[cI��b�W\,�2��י�*=O�e6����[�	��L��{R�\�_���6�r�$[�୳��w��H$���w��v��E<�Yѡ�9���4P��S�zp�L�1�S���B����Hpf����������z��YMڦ��H����,hrǜ�ۡ�ۊ��񝺚��K�[���؄G���9�?B�4���ODF�2�Y�Ѻ��l*��ܼ0osB�Ve�����G`���%2e*�1�'#D�	����7[_��1�qh
�sP�M���^��hb��@�U�n3	yLG�N����(��|e����G*��,���	H��R��t,��J���o��Z�v�n�6���e�_�^9�!\�H�y~~��*���}�$�T0>i�4qHbT`����.�G�!N�!��&.��Q�	4)ȭ#���-m��Vs.~mpE�$\F�}�TH6=3b� 6���۹��/Z��!Q�L�%�J��W�6�֮v�l��]Y���	���CDtsGcՁ�[�b�\�
$Y��)�-�0y�I'�x���(57��d����k �fZF���W�ո:����	|QE[n��o�'���X�{�ս�v�]jx�8S�9i>h����A�ݬ��Ήk��4����a9�9g�d�<�?wg�h�$+�Y�P�η�u�y��Y�\���5j꧷Z���2�����k��q7�l�7`���2+�0��_�K��"k��#YZ|�f9|�O��ɧ쾟��ך
�{P�7���I��3p6dj���i>2�z���`�[�"������wp����Z�eM�f�E\���B�p�{W���J�M�o����m/c�E���*x,څʓ����5 �Q�%{\�|�C@��籝��b�� $b���%��f9 `	�8�q�Cϭ�����0�y����!�ݮJ)�'����h�����Dģ�i��6����
g���Д�����T^f&/ZIB�8��Uf]tO����_����g�v�kU;b�G٬Jj?`��x���������tD�b!��2��7�D�O�o6����[��Ӻ�o)*ܽE����CI���N�� ��r˸c���G����� �E�FFczW|3ݠy���}�SKe��k/ܑ�>�7fG|��B��Rf�|��Aȳg!��Q4	[<���&�"�}"^A�z§�A����=t��~������Ǎ��f��� 
��9F���F�oT~){�E��ܷ?$u�l��m{�97N��O��JxɎ�l��̗*q�R壔g8gۮ��0ŞCDhI����zݟm߆�q�W|�M�s��P`�Ȩ�IXQ��⯎�]��Óm��R�o�`�#�-%o��g�Iۃ��ŞOq����Dw�l2��-��q�'� ]�#|�tel�����Rģ�RXџQS��D�i8�ӏ��M�t�����R "c�����~ֲ�ʌ��;�D9&�g@C8t��%�X�K��ېr���T�i�)��{Sx���X�&�.i��,�٨��ii*��$\ϥ�$|�Э�u�_]�"\����Kx��d�\1)�䑳25t�@���w���� �S��tt��g�S,�8��%O!|s������&*!O���K�1@�tQ���v��^�#I/E�NON8��Y/`DE�=y^G�9�:k�i�\N������I0n����'a1O�Ч~#>/�.�Y0J3i�P����ÍF�D��YAOS��A�$��Y.B��H=c*Ƥ0ݥ>u�oBK� �כ�%�5w±��X@4y��9`W�<�8���)��W���6g{����ɿ���d�
z��w[B��m�0�	n�I,����}k�?���q�� 4�K�%1$�:e��J1X(�#�?�=���̰�sv�Z��K�0<�*��b�-ڀ ���Ђt���� ��UP��J@A�/E��~��5�>
���� 	k��A񖶗�j�~T�ܶl\��I�{ɇ�"�	�C���*���|�4����Sxϝ��G�D�f>��BB'�4���͡�`>L�}d�WAT �5V���KC[d��O�����ħ�Vo��t3V����C�Y	��d�H����D��"�����ӗj�I$�b�I�8��c��F���~2v���?�,��3 G{���P��y��"3!�כ f
z�/����d���>�yd�"OM�'.�D�G��:��=_�t���y��T5���t��Ѿ�_S��B��r7aay�k!kξl��ۻ��/S��-�+[� x��m��ٚ	�'�cs�pS�B0����Øm��q;F�E�O��E�x�a�/�; 26��&.s�Im3>��?��k���u�?iZ���[-�6� 
�ʉ�<sPp ,���1���^%�x�֡	����gD%?B����JTf7��"Y��i�#��1$�<��SF·�S�퉕�/���R�}�+�%��t���}�>-|�f�0��4���^�H7j�4>?^�:n��U���f�� �y!���
��g6�Mqe�3�h�~�k셂�v(n��
]�`32���ZO�C�ʚ�dB��>=�"���z�[�����9�\6CQap� M���WK��*�T�i
����Rm	�k����<~:C��b�_��V�Q�1ŞHŌ�e�dYZ��b�G*�*
�;���6�y%���2�hո���.��.zڌEr���a�^̍(�5���PQ���ym7���&�ǈ�VE���16����>��]������L��_�r5��nOֆr#I�
i{H˒5b���_k@��qLS��M�4���W�x��UlO]�������+	/I���p�7Y��S�Qa�,�r�n�ir�S�Քo���_�ul�խsĘ�<qhR�P	(���1��>�K��� ����7͇�^��d��%��~kV����e��q��z1���������H<FTH7��F�fp��a�2+���4�Z���k�Y�`�KE�d��ܿ]NF3���)�|�[�� ���^�lWZ��ך�k�mϨ(�!�{�xq�u.H6j5�璥�,��mT@���`���|ۻ8�<�L��A�\��l�=��5�
H�N���b��Qv��g/�l��l\ˋ�޿!�m�l�����f��.f�&}��,^��Bh�X�(�a��k�8�>bvRƎ��Myu�,���ׂ�~u�s5��Ӹ?ُw��0�Is;�C�5*88�SY�ȃ+������^xKlG��Ԃ�>��y��� J�g"�4^�!����k�cH���>�-��f8�j����<�51���w%�୏�rCd�xE��U��ņ7�£�8&��ڏ��"��c���F��S�����x��_�3�NpQ'_;���['���y=�o�u�Ҩ���q:L��+a��cW[#s�OV������T�^.���E ��Up�,�ԇ��I�f ��N㓊,^�v�Y��	/��Eko��4�M)U��<h���>��n��� 6���m�k��O�z�&zʺrp�Y_!���;���OJ��?�.���\:�x�5�T���Nb�� ����~1��4��hc x�$�~&����� ��BT$�?��G�ޫ1�&���G�F��ԂU�r�26d|Z7����e��t\�I����q��L�q�w�ӷA�=��]O\rh�_ßt���
{\/Ee�N��_/$әF�u0�[��M�-�9u֢��h6�|f���^���*"�����t��/&�X[^��P�Y�u`I�Ce?G�wM��o�B���M�rh�D��Z2�H[�;&��<g�^D��riҞ�50e}�>�;%
���R�]�(ċd2�.�L�B+|��g�����U+�;�\��;=I�i�{���[��S�c���i�gE2��c��z�RH_\{=|�ڰQ��$��K\Hi�7�GN��a?��K�D@�����{l�͝ބ�1��s��VY���R�~�}���7c7�y���K�vl'�lh���v.㮿	+~��x��xay��������*�����@DZ�ř|ٗ����k��u�K2�/�P��|��P	OH��b*ib��(kbJ�`�؝�(E1� M��I\��6�M��%�.0���a��zxDB��@��6N)��[T��L�k�S�T$��ZF硚ٟ^�MA�HH^C���8Ʉ+�<*�zr����u���Ԇ�r�{��|�0;1R�1Z�]�8'Q�A�!����bJ���'�y��$�۩�YA��R��Ҟ���&H��)�[7D��B"<nB���y�롅\�41H��a~����ʷ8�y���6^R\�ļĵ��w����9���)P����}g�A3��i[]�L�-��'rj����&D�P�נ�Z%�>�e���r7���#d�Iu�qm_�?��18	�q��d`a��X��֑	�}��uW�����)��!gw��i���^��Ai�QF>��Ihh�t��HR�VPru�syFJm��ӟm�o��Vǁ��V�+��7���c�c�Ra���EMd<tj(˺�[B�x� pl?H �ea�-���aȘ\(�W�� �L�V��4wo�� K��e��� &Zd�Zv�jm�V�)��XR�f�T"a_�0Z15��R�w �x'=���AZ	hW�!-5y���Hѹ�C�r��_sN�����?1�,�vQ1���o<����cs�y���K��IgB��C��L�e ��(�n¢�@O��x4{?S� s_Y���^�(�f�r���Iߟf�q�o���4rvd���P�5~���j�8͊�_�*%d�D�ءF2W��`���$}}�y��$-��4�!�Rp�U�n�zN��k 6���.�DC��D���ӜXP��=Th��� ٕ� l�`m��Zg�*��}�#���c ��aЄ��]��[4N��s��E�,��4��+AE$]�%ݤ�_�;8��44JH�)�2��5�ӕ�q�L_�pf��QݦYѸ����f�]�La�ُ��TnP�3m��� �b��t�;E�ũ�=��N�-�i�;<���}KXWd��s�p"���0���g�M�WX,ab1GB��F;��[�@%�_Η��, �J9��Qx�Q��yga��C�� ���Cy��*�~��Wk��D��M��L��hģ`�锁E��U�*��ؚ�{H}}P� ��Q��NI��0]r���*K�`9��ep��p��-=���W���p�T?g#Nx�PR^�a�>ݎ�Yn�H��T��
I�Z2����6Fyt�7k��.�-�)�R��Q˿/N��I�y���F�yh�e���!��w����Ztz8��Y,�7�+!��d%Q+�`z�Q��IhI»��*l:��Ҍ�)��Y�N�`�(��8��=湽KM�%�O�^�N��.k����X@�Gp�^���<���r�Q�P�k��|�����0e{�����Gʱ�{�1�ვ���>�O9ll�Q�W��q�g`�=*ٶ�Y��p�Sj��/<Z؛���Hԃ���Y��NI?H�*���ξ�% ��ڸ���q���qC��Բ��7�_����=Yr��yV�✑�=�`9�8�C?-C��k���)T#w�F�lM�O��@����	�ކ�ʿ�)M��9�rdf�S6@��WA�2���(��~y�P",D�- p���.�8ޠ�aV��h5/�f���x�u�N�G�(�B�?�*�i]i��~
	#��QUn�=T��űކ���@"�
us�5�g7��a@\�t�]�e��t�_׾ ��W(6ך�/&�t�-D��-@�� ��)'�*���]c������\��<�-�F�0A�a8�����KFk]�D����RVn�|�I]]����e��-��h��9�_�����?j�Ջ6+yF�i;�B��&��-�����-0�Qiׇ�D���/ݥe����A����˗���$t�er��c�$���(���d��b9E�.>O�D7|T�Y.6�y�72��u(qC=��[���y�Ow(5 Zk��/K�B<�����~�.�*�X�?#�⊰�V��-f� F���t��j%�N��,_X�7�fʼ�8x_=�����:�,&�M:�l�����:��<b�(�������4A�56Ӣ��멮�_W_�Q���M���ߴ�=]��Ō�'H�F"�=(�6W.�������{��U|7�$է�wc�J�|�5*�Qڢ���O<ZY������j�����:�5L�>���;�-|�J!���ˈ���**&J�5�4��bo�,�� ���k���SI��V��@��G;�́N{��2��򄟹/1���;
3X� s���^��'�կ�?R;��>���B��a�{GJ�X��
G�Yԁ�Xo�B~���w�Cn�et�5��C��+�,WlKk��A�0���H���3��c�^��c��~E[6Nܽ��n��lbN�xv��}A���{� N{ǉz���n-ʬkmgh�KD3�e��k�o���y���<����Nzɮ����lU%zҫl=hc͖`�����2�}l�P�rM���q0ӄg���Ǚ$8ǿ�Q:����]�B��M��ժ��J�"�k�f�^"͂GW�8�Y|l�6�=����;�EE,�n툙���M+Y���G^�k���ٺa��c���$���֩w��+*�Y)LCL��jړ�f=��o1�%2S�X�I$=�q_bJ+h �cH����U*F�}I �qD�*��b �y 8����.U��SA����C"
���K�cQ��~Y1�P�$��bB83� V�6t�VՂ�����}�ط��G�&;���]1F]����,^�.������-�<a����n�{ִ�A�VX�8�AQE��q���t��k�"�&2�� �p���S8o1���աx���
#p1�JY�w�x~N�u���	Te��Q-P�0��$�@�,��fdq�wq4��,�ǂM��~�O;�%C�����Q�Mc���q\0����PM�s�-Q�E�ℂ�θ����ׅ(~��H�����dG�B*���Q����`5��dq��5rY�Ys�w��T�n�[C`h��S᪛ a�e.u*ۢ�g��H1��QT�,�V֛�'�`�ݦk���t��>���ɒ>�m�I��BIX��٪����"�F�t+�|��h��=+��c�����tD0�)�4L�OΥ�C�sߦ"K��@K:����l�uN�bCb��묥����I)!�= �{7]BHt?Y��.c�p��[N��d�T"h,* �@�Շ��U�}�60H��ߚ�)�b�p�3�75��0�Ihm꩙�3�cƩ3ۛQ(>܌`&�.���o���>���%άtK�ڶ&^�B\Y�W%8Ѡ���0��z�N w^�Wy�eB�1�=�:0���z�φOSǎ^WV���4�`�ձ߮Ͷ�ڄt�^�[�Ε�������S�H4�nlAj:ȷ��`]�s�.<��[Q�%/�`4R�d�Fė��b���@O�&��A�:^T���|H] �o�Th��߷�S��{.#�@��Ö��<R���~fxb�h,��gX��������X��Ŗ�&��|�Z��3cYlC� ��|*�(�Ч��u�儳U������)�ta���.f�ktE3���<84��Ce�.��J"�_G����4�p/��������ĳ�>��\+{��	v����G.рJj*�74+���DK��c�䑂 0?=wv�'&!��6�&ׁ����gmLW�Kۀ}�:��k�WԾ�ͯʀ�BU>>E#���h|�,��yn��8��)�~��� ��V�qA9+r8�s�\����%D@d4��!
3��P��g~�ب��B����Ta#۽�8J��������2{��:���Yq�D�̜� H9��w�����	k���Iy�j�H�\@.4�X(��Ll�������O����M8��Y}a}R���<��ܥQ �A��׮��1=���sM�rXK( ��\�+��b�������K�(��ŉN}�Ҧv��}���%������  ���[Q��b�������ap��u�F�pEʸ�xJ�~��i�t�[�����/�� �2@����I��U����^��R��^?�)��#~7�D��4.]Oq����{�b�~
�����Q��Ƅ�p�tb�Nú�����;�%������En��[���RU�J���[��?Fi"t�����yY�嚦CeUAm�iKi�C!�A�y	"��`!�̮���)�`zJpOnLN���8M�l>틒C���%�G������r�tG�`'�*9���a�e �1�G�Z���7��rOd��!��O�T����W�
&��T��	N���ȓ����XI�V7�@����l��k��1Ĵ�!K���޾a��}��^5��������p^&�}�ͳĈ�t�>7�HX�"�f%2RY$�M��ւ�y[��#eya�K�)ɺ���������F��v��w@ύI�����1l4��M���xa`�8B50O`x�'��`$l����Ř�:��Q�����]1��q0�v����x����2�gB(t�u��ړ���e-w�TΕ�2��?�����_�H���/�����/�}'%C�0��#�Y����>{�˽�.�1���p�� �ltIP�v7�h��jX�����b�{��Ha�E�2P�s�ŗć\���o�?�-��(Y���vi�-��T��Oۂ�\�����I�(/�-��D��}��x������Ip�1G;�$��\=�ιj��U�$�@��T'!P�̋ �`�6a<Z�9�a�fP��<*;J�qӤ�R1��l�)��'�䴦yi�"h�a�5vfY�z#���
��*|�esW�^��S���x�! R�S�B�d����!���Oy���uN�{R�t��c��g�k��~�~Jf��wW�`�<�8�k��TD���P�f~E�������u����T��@�Ö�[��`nh7*�����V;�$5j�n�����7��%�g�<3�A��tor#�*�� ��r����Q h�Hd66��h:ctk��6ƒPv����h����؍��*�嫪+��[v���\�5��t��
�:C0 ������Q�!`�r�����cb
g޻I��ɼ����d��������v(���z���ז]ɺπ�����C�esT㓩4�BVݽ5{t���p����!la�gO>�_���L��W����{�_LĮQ8�A�H2[��{�x����l1�`���=�>Y8��jg�X$�y�3��;`-5Wn��69)�OL���nO؝�Q"���y���.r�)���qd�q�j%9D��͘��g�򔒪!@���+HT�b~,� x����ưAl|��ec���^�|�|�i2<�{�h�MX�A�m�������&�:��~F
&]���S�-	E�9F"@;eut�Q��Tpx�HU���@��FDn���k��\��9�d���@�FpH������!yY[ (�Mn��e8\�1h�<�����m�F>ģ�/�'|!��)x\7 ���R���u�M������"��䘛����ń��FMړ��z�<��Ǽ��J.S>�Ɓ��3Y�`�kn>��U���$Rj;��{��K.2g�2����B�_��������V:�e���+M�� ��[�};4@���5{B)��)�t�HA_C����Wq�U�MfP��&׍�#@V�ρ_3� ��Y�a�AuD�	�þ��w8m�Nu������=�]s֍��\���e���<�H�2���%��51e�
�R�
B�����-(��(H�9��)yu��*����|��h�'8�n����d�)|Fdyuɕ*��ў��B���C�ŃЀt�'g��֚�A�P���ʟ_Lce���8��K���h�%�; cBR�{咂Eu�sîu�t�e���s���T�1�d�濿5kҶ�CN8���NzH�p�������Af�r`��7��HK<�+��#�M@P�͇����a�X����^�7½�a>���egd�N*}����6�X�MkH,��|yɸ�N'Ud�F��z�:�p*�Q�uQ3y#$�C�Ȉ!����k��]eh���1��ް������#^����cB�i&��х�Y)`ٻxi��W���~���s�MV*2E,��ռ����Ȣ'j�`G�����?�?��J��mۻ&��;�@��<v�W���W_�*F�V9�Q<mDLޭX��H b�͍y��ͪ,z�g|晓bĶj;�8����N�*|�y[��kz�^.z�5@H4��ӝ+���$x>�k��m(3��(�,J�_��U��_�D��UC#��Ǭ<g1;(=�T���	 bT�����	�'�+\���M����r���&�_��M3n�&����oO(ǭ�u�!)��A���t�q��)s�w�n$܆�*ʝ��?i��[�m���i�d:�L��0�w�늹�L�T{J�AQDƃ���ӝ>����Y>��3�4� �r����a�7B��eM��Xw� �ȡ�g)�+�Xg`%�j�cؚ�t�?m�pB��,�b�� �����gB���Q,zy�70�s���R6��U@R�5��Ծg���_$���;�5��E�L�Q��-Y���\����T��L�C���2�e!�0^w(pO{W�7��J@����������ޜ��aU)�e�\B;7�U����R��4j$!�`%��iq�s�G�F�5�dX|xZu����|�l��e�T���
L�dZ��؀���B�!t_FtV��m���Z��j���0�1+~�T7F�~9��Y�N����`V"�e�Y3:��o�>B͂UH�����eި����\=R��w������,u\:c��Zss!S���f��'쥯x0�6ѴY{�p�D%���}B���W�6K��l@6z6=��fh�=Ȃ~z{cB�5o_M�>�P��$Ɲi���Y ��g�I��k� /�q4��
ޑ�=۬��� �{Ao�n���Э�J���E�Sv�O�Wy�N��O���.6��n�ҸL�]#���T�M~���O�n`�O����R)�]$y������W��A��$����.�/I�(�.����f���A?�! �fzt�x��Ļ���S�|�e�|Y�n�ig��pݟ��,��s7�λn��W*oP�GH笯D��F����'ʻ<��pIX�VEI'����)������
�F�li�+��Ʈ �4���pݎ8�c���՞A�c�O�J|�6��H���N`��;xm�|��N�D��^�b�:u��'k����
�o���BUQyR��_5Ր`l[Aa��$���?F�cg���PrP�ݙ�R�`�[F�Iv����7X�O�e�t�ϲ��TF�ЕH��-�A��07mpG�������P�/9�-�]?��9R���'��]8�sU�aY�`خ��v����H疴Ut���Г,���C#���5���&%M�{h(�:�ft��$��,k Q����Y�ۉ�'~v�q竻�6��i0�2N)�����+�7Ҏ��JR�L��ӗ�h��:�[�p��ц�Q�d���� m��sJȃg�Y6�(�18U�/��5� �+�87W@� mp�� R[�dަNP
u�!��40D;N����#
��gtk�V��>=��V�F��z���LS�aԈ1�;DX)�1k[	�N{�.��Zg�Z���E�~0���_�(��=A�5��L������숼��uS�(�o���XW7�S�hK����ԧN�`�=S��6��;���h8��6u��h�[� �L��~��@�Vՠ+=]���S�P,i0!`���̊��\C��%���v\r���ct�5o�!D��w�`QQ|/�x3��Ђio����
~��H��x8g.�*��t�#��7����>�H��4��M�C3ᗭ�&�%gLF��|嶫2�z�_V���h�Ԫ
5^��4�8XN�2�!�/w?���7�(gd�����n�c�[�^�1iY0C}K@0�}��o�g��w�
Ei��	 �7k���`ͥ�B��1q��3֩�L,O��&�0g��؏�@�+|`�mm�/G���Y�}�v�#I��J{?�8�f5�9j8�
Gt���1t� ˕���S�:�u��8Oa�h���9>�ӿ}�4To�.���&W�ƀAͤF� �ԅI����ESȸc��AZ��_�K�sҌ[B�u���<�3���3�����p�	�G�r]�r��JO]�]=ɪL�-���o?��4�g2hq%O��^�[�#�~�3u��({�{�:�g+0���՟/.��qj,c'��ew��Ԉ��z����$���bwI8�ۄ���pp�������ď��0e<g�Q>Β�}n#��c����QZ�;��(z�Ҟ�ҥETv�/ϣ� [v7������X��
� DNđO��
6�,���3/��%u�2YQ�tp���г��	t +k��&��&�Қ�����i�+�,F;BO:��p���L����g�v3�5kĘ�(�$ԭ��K�[��]��<�x�󼎡�M�=�L⥐I��*�Eɒ�A�ֈa�Ȅ��MC�������#9�̎y,�������*��P�𧻓խ�+n��;������İ(g�a|�,�O|��_��VFC5��u`�gԎ%��?i�'j�4�p�cP�ɨVO��BGZY8�x�HL(:z��}�*�tC��d�!%'�dx��	�)���41�9O�>���es�?צ�ޥ_���/j�?ѳa(�P������l�]ϑN�ڳ]j�OЂ�o�PH�f�s���;�e�M2����tx?w���q�JN�9�*=�;@u� �T��gΑ�I��O�������C����'@�(q�w}\c�����Q��ݹ����J#�(��V���>�"���=G�2��l����f�Pܢ���e.�ߗa��ZG�e�˰�Lӫ
�g@g�b�2:�xݾ�iS��Bj�"���Q���w�$NӸ}*�<P���烦�:��>������%B�R��H:��_��ƍY�G@�u�O�N{��d���y���K+���A̎�G�<�ɹu6A�ֈ��:��z�J���6� ��m���]�/�6��*G6f�hH�z᧚���W���(���O�[�z�0�"�w����� X����}-�E�h��h�&���t+b����Ln�2��^����\�pXm�3���ڒ9d���-G�A�we�4�'G?"]�ȃ~��ے$A�A�m��LG���#������å���pW�u����<�6msX�5��
����Q��u�9�S;��sL`��|��j�i�����4���� K!�b:�x}��$(��a�qpc�kj�������o�m���$r����CP �<H_G��5������u	I�*Y��"}�Ա�����b�F�c���ó��N�}t�`(��Si!X��V*�P׷���xk«�+�f�ZlN`�M�B��v���R�}�_d��n�]�s�oG8[5	}�{zJ�zVWH�ĺ�QrZ��o'�m,
[.�,��H��SS��1Ha��Iy"	s�K��
��-dC�!��f'q��� 䝲j�Z�<�P����ml��"��O�fj��UfvME�ձ�<���
�6=��]*[ʶee�u./tV@dsl)� 4j��ü�`"�wW��ו�f�[\%����CX�0�`j�B�Q'�")iV���~���)+L�q2İ��'V��5�ֱ�%����/2�=TsL~��;g�W��!,n�����t��_�W5zБ'�,�C�89�J����0bo�D3�vI���ZϦ͟EN�(T�~��QU4X�4��I��� �k �1&��%dT���D �,�fspt��{#o:v��?���i�bX�7N3s�Y�K��5��IQ���q��C@�����u|�_(� i�qA��y�3�g[����B̻��;�y�1�Ħc����s�[�~��!Oi����]���梫<�vb��7j��~n�g�9�d�_���/��qLQ�td`�K�W<MS���#�5�����S��P}��5�5�f��ƿ.5��~�C]�89p�M�꧸3�bdk�RN��R'{��C�c����Ꟊ�j��3-�# � a׳��dB�k"T��ՀJ���؎2d�G����r�$��c�?���.����s��D�4haEp� 3���t^�ޖ^�q����-h��e����~.SS�B�O��"�Ƥ�������䊈��)��ȝ���Rh|���̙�|ԖGհ٨j��D)��W������8�V�m���@�� ����̩R��Y(~���}E����r�e������,#a�%p)"�_÷:}5 u�Ǌ҅A�&�ul�{��"����&����׌޽��;CQ����Aݯ�7L��ֳ#��9(�.7Z4S	�{����t�	�������*��[�;cH�s�[ ?�wTF���S�i�i
%n��q�i��no_��1|��Y-��h��h��*C3��S��� Ʀv4vE$�&�q��μo\��|볙/(Y�;�_�s���ma]�����}��T@3e�C,7<�%�#v�c#@Qa#mV�I*у9����>ä�nn�H�^�h��ֱ�KE���[�́�9�ڴ��0�x����f���7[�U�.�n]]-�[>������,�� m��jŪvy�_���G�26��@u��-���[��<���=�#��5��[ɍW0
�e4��uԖͣ*X��!�Z��ՠՍ��4H�?nK".m�m�Se����pw��k񅸕�68�xF�����mo����-O6p5�K[@>-�!;S�77+��o��) m�U��E}�ʞr:�q��Q��p&�N�l������e�N�T����.>�ݠ����,Z~�U<`5S��r��`Q��B�e��V[��îZ�z8�����u�*�P��?�r����r�ʊo1UXQ����C/�����	�yk�n:�Mľ4+�}�R���?��vc� ��lm�dǚr��va�BA�d�e���ή��N�R�3 ��vظYY�{�$�aX���p�^��)0Ob�J��3���(�R��qπ��1���)
vU�@��$��CC�;���!IbJ�A�ֺ�/�.�!Aegl���U��Ï��Q!V��u��ˤ�"L��3\<"�3�=�9#�Ղ��I�5��V�����(�%͗4�ᨐM2)�j���Èӳ��y[��Y� ��b��^��T	���#M�Ο[*�@�f �3���((�6Sb[�w<�Ƞ�P��|,�e�"¦w	�q��;�k���ׂ�3�K19�[�w�IT����꿥юi�֚���Y�uvH	%iD�b�o�B?�U��1v�}�/�<_%��/P�A�vL`��u����٬L�v��xc;���U���%.lT���������M�b�`�q��ti�;�+��b0������^�zD���dԎ�(�?��jh�쓘�7k`\�XS<�Ba7([��i��[;��3�bpTb6�mk"���s�d�,y7�,���{u�Q�A�;K�x�!H.f�{?��g0��w�3
�L���L�S��7I��B�N)k,ri��3���~�s6/dv��Ui��K���� �:�_t��-6x���9�Lo:<_%�.m�)�i^/��t���O��	�/}�6���r=B���(���^Y�@�!��l5�w�(�8�#��Z�N|�gvΐ抧�c.�ć��]^�GǑޱ�3�w�uga�|�Z,J[`�D���>~}g����*!E��pX�f~������p#>�mV��	�_�M���;j�0��|�0 ��u{�,7�̍�f&�IU=Ka�_鲌�a�Y���g�㬑9c�~g�����עd����EK�%�˺�l�0�Ћ���I|te�a,��j4����P���2ꐒ`0z�����x��OP��$���f��x�
v��@ѲqG%J�xk��	Ȯ��M��߭�ibO
2aFTHA���2����+b^6���l݀���ѧ|�)��<� ڻm�؆��(C��@֍��X�`��