��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�����9p��s���v���	a���y�A��n�M�1%�P��Jl���� �k�
:�q(T�F��l�F�j��;*Sc�e�op'Ho��$��'�*>��e���y������@�%X�9��o@����&RY/�~f�C��31�qĄ�J� ���2��:<��-��q*J�����>+e�!1��]4q§ �]m�ԫZ����v�����F�q�S��8�00�F�ړ� ��<��T�@d�Gu�!�h�����j~���C��P�Rc���FfxXs�� PC��԰�O����p32iXA�t�"�Q��&?,P#̓�*eA�9T�x��0�8nVHAG8A��J	��c���G܂y��S7AC����&� �?�,�	�B�Ũ��aU�P�̧Θ꾸^�����\�(+��F�I�j�z	�Ϩ��y�g�8!�2���%Q���_�m�$�x���b3,B�6����9�@fZ{�G?֔H���R ���o�;��Hd�����������O��3�m.��]k<�B��I_"Z�L2��:*p:߶����aȈuJ�L�_&�݋�w�����j3�����:6���Ɋ=�����e������0|)
m�N�|[d�)��H���ڵE��Jq�)Tꗓ&�^`kC��O bC������h�j<��+�E�v�)��G�i�SN�p��x��Ǔ,�z1��@��t�ܕ돹S��Iເ��8�^x�)�=��V�fE�s��a�3c�e �ɢ5xE�'�fr&��W`��r�E�m�_R�W�(�|1��hR�%�O��p�ʼvkn��I���T;6�<���d�Gt����d��qkcR��H�5=�E�zD�YX�k���B��&+8�w�}��3V��Cbk�9G��3�����h���7�#���J���j���d�]�O�x�kk�J�1�A_��,�&�:�C����+S+�p�R�^4fN���U81�{^��_!�R�q�Da\��p��{��Ox�o��,ȕ����
J��wܡ�V �p~�P�l�}8���KP��שX���B֬ȼ���_�R_�?Pٷ�x��4TZU
�4E[vS���J(R�v��3��C
=�(�?�0*���p�
	v/��}91�v#��kܙ)ͭ��2�^�t���m[_\ �u�hz(�\r�=��fG�?�5v<	���+yvK噘�c���%�#F��&#�̡�9���;�l���r�-;�����WA��6U���6�()i��曧���ߍ#���]�sI9���a\*��tН�}�okI7���U�� m�X�P�w����3��N�7�C���m�ĉ�)p!,1�"J���4�'�mm��g�Ԥ7����@��;��M`�Q�>aJk���������ee�6JSH����0u��%�dY�4���;
<˪)�XN˳l{z�y=��W�쾗�&����}Fj��>���G��\�}Yj�����.ݼg^�ee����i��>�H�����f�^��g@V�.׍8��'ȩ�Һ�M3�cQ�&�LhL_���YyBt�Da`�G�#�u�`j������ʁ0C�m!�ƞ^���s,N/)�&c��5� ׏�w�} ���=�v�l�fH��C���<d��l\wb,��(h��,G෌���6&*�F�<��o��f�H��"���XgϨI?�[�-�'B<O:)����E��򌵱��]��dno�B�$�4CN�]�=u��n�o��<S��C�a!�ŗ`[�yD�n�<��!�Q�G����Ĺ5s��&\��
ޭ,h�������]��y:�%��w1�<�J�vo����c4��	=cΌ����1����8�Wˬ	.���j��?	Wg9�Я��d�,E��A�9��s���y���}��<�Ș�2I��������:9띩ۓS�9�{��{w�_�7��qt�RP�г�������cr�1�.`�� �u2�ڵ+,K
H��cHiN:*�$�7z߸�M���~��i�O#�N(�CK~j\+l��,2�(W�q�<+P��)����#mD܅�൳<��^C��s�vgOH�pB��ݜ�0��/�IoG{�-��co�΃'ܓ�E�<7J����#�?�^�*�����BH��8Xk��QQ'�r�m��C�e��qm����ٚ���{����<���\�I��ԫ��\�\3H�m�8�S���^�ȣ������	��6������^��L,6���Χ׿���h�
��?p��(�81����hc:Frc���C���\����/W��_�e�4������_�u��lԗE�oE��=N\�v�f	Kg��	C���,�@�4�nL���ʇ�����o|��g��F�� �K�A_��qǜ�"ӣ�?��+!��JAɖ���J�'j���sT&����[x;�����A�%g&�1�;��Ҷdc*]:�wih­����P���o���8��*��U�D�)��G~p',���=�_��83"���L4������ں��#J �4�z�(C�Rp�s�o���g�Ǳ%Q��u���A�ٖO�c��tBT[DӆM`��IY�x�+r��on�ȉ���d�ds�d��O�k��~6�F��֊������������.^hA+=��Kм%��H ��-�IޞC�I���)��K���&��L��@p��P�U��[���A��w��xT*U�@ �)9(�k0ݜ�	���(����w�̒l(�W��,�X�[�t���`/��<����R��(��ѣ��]��=!�ܦ�Lv���s�.<{=��У[�����`�|o��MX��ȣ��T�ĥ��Ӿ��[ØټKʼ�V�������l�Honѓ���2�m�''�0�8�cw^T��လX�4y��;+5��L_��@��G���b�5d�GG�~n�]4�: �U�2Ŋ�4���}�X�n\���F�cq(]�-���C�6nT:t��8!�?��/�_*�bf��aE�k�3����Z�a�`�w���������*Sǯ$RoG{]f#_��I����;"�[�S6�{�Gl>��)?X����h��WWh7d�	.,�9��M.�k&��]�3&�j�����9�9ȤP"[����hZ'��0��n@5N%I4E�n����As|sr�:8N��!&�B���^,�X�Wk�Cg�_�2a��6��C2v>��m2�e:���<��$��"v���<JI�Ij���Lh"�o0��P����6��l�����5� ��6w˙��Ef��]��q��Y~S��B��3��l\�͊��U	�s�/� �;�]+W��hI	~IX�9�Onu$ا��wzg�#ZC�Jm�Z�(�B����y 0)ugQ� 0�N*n���h/,�p]@�1	��3� ��m7�
�����5�ԓ�+B'0�qW�Tژ�������}ۉc����Xϧ��Dv�;�"z���c.��R��AMY��(yM�"��Py���;P
<��A�aS���o�f7�!�,�r��`I�sG��Hx�ĥ9�+�pR}p�:����b�M�Ǳ1p��;�$�9~�:%�N`ׯ�|�n�;�!�m���)j���{t�ˬ�d�!�`�.R�(OWH���G��O���1� Jӓ]{1^�67�"�6ol��y���h�W1�}�*$�%p��A���P9�#G*�쓘��b5ٵ{�u�Z��zwwB�|(�ťj�5([!�ݡ3;U���('�*�8�� );�l/�F����Gs���?\�/d�O������y|Y���b(��j�C�d+�G3��gf�6�E��q_�z����N�l����s�.0���=�Wh��I�� ��ϧ�ϫ�':��i2�-+����O���r]񿾕�ޭ�V{�MX)�w�T�q��I�4�-%�^̓�N�G�1�
[=BR�J�6�4]����@�5=6���Ė5�4U?G�p�s��Ʀ�V�>s@��3����+J���#o���ۡ��(��Q�S�$>��3Vg �m�%1����O���oL��x��v��t���K��VI�_�h����m�[���?+�6��:,�n��%�j4�Ǜ&]}��j�f��"�f�1$�J�qK=
��	�=��%�5�������G< -n��5�BX,>ĿT��������(,_���9E�i
0�M;w�t_�	�gv�1c����
��p$����F5>�S�`L��Z��p�١[G���S~�����#�>#�l����dKrzy�,v}���I^�3#6��Z?�|�PH�H���T��q>0�Xw$չe+R���ē�����Z���o|�8�E�՗���� %���m*X(�^G���i;���h��:V�gY��R5[��w�0��7�U��7��2�`�E���Ԑ.�����?2�40�u����Y��е��1��zך��b��y�F'M�#�f��@m��`$����]Ȑ��3l�Or�*�~�_���� ���e���� /����F��[L����Gp([�g�n��Z͸�Һ��B��b>0,�D��h4�SZZw#p ����E��1���6�~�(�b��D[Z���=��e�8����c]:2E's�A�m�_it��Q��W���C�d:1r)��~
��ΐ+��c�+>����.)��j��"R�BP��r����SvD���f�U{!O:J��z��M�"���p�G��۳��t� 3��`E0O�U�l����Nz���˚��ut5�'�1���z �l��@�X� c��4fMA��W	��3�g��$�W!�<o��S<��h�$���C��;�FD+?p�G��N,�����po��+5�.ï]!��d��ڇ�_��㌢dD�X�<�Zx%\� ��yv{>�-�B>
�7=W٦�(��Y��D�0�G�Ґ*��9.gn�E�/Ϩ�,n0(�/D�(��$"
S�[�J/�]�jl��x%y��N�	���	����%���I�t�Ě�`�~����z�J������-S�
��U�j-ܒ��g+y<����,^ږ�LU5��\��u� ��g���C���K$�վ�Q�-�u�Eޗ�Rsd���8�����H�J`����%f%O�A�{1�[�lTK�H ��Tq���W��j*�$j<�^���ȇY������A,��f`+�.�#PBg;���� 8�:������~;i�%<��BF2nW�ነbi�gSʭ�����-`X��r����+pK0p+�'�D�ers�"h^��[>������^�Նp5�r"J���%xٿ3�ٜH '��Zf5����u�A�PE�,���� V$6z��H��)e�_�;t��éA#X� >�O8��;�A�	"2�!��7��'�۩�C��/�/�lr7�4ڑu	cQ-��9�T�bh
�*C7��:����e��9Lɾ���3#`����k���D�p�A��Z.��D���ݞi�Iz�u9��d)9����# ��}oSٰ%� #OV�*��EۍQI��s��cy�Z�$sV��I�t�g[Iu�0�u�BG�Vxt8���M�u=772�/�4"s����k$�����X��,�V�6�����%�V5\�o����U�T0���KZ���L�����L,�5���~���zq�{� �5�Ab��������^�-�#�Z��s�/B���Ɵ��݃�����w�R
	T�	U1M$��&IoۚpPĶ5)��ʍ]�k�{�H�������f��M o���|:(�+�(� ���/VE'NO#���Є ZiU˝D$�쬿d+{,I���%)�Ӟˮg��T��d�lϼ�
b�LeȨ+ܛ��黜�w԰>^�@qX�*�}��݆>��f��^��+@�C��F�}剳�)/�lc�8����n%�
�g��S}6c�~�����"��s�m��vR�|��kH[�"O/�<kn��7�	��@%>�n�#���/��.����� �T3A0��Hjڙ7�	�c��ȱ�&=�눢��tC�����GcP��|.��\*�7� r�>���_�{�m�G��¥̅s�z�x*csW����W�����@)��-�Kr8)gO!p[�aɠ�j�o�Y1-��Q��E� >�͙�w����8K�#V#�)T�B
�l�� Ɣm��W����CBZ^�۝ns���8��Õ����#��4'؍�,�%�?�r`i�X�}�Fg9�'��:5S�Y�H	�PPv�������)����f�	͌��25�-��K�a�_�)�SX�/����<�(��MQ�^AE>��h��M$�6w�G�+�t��yC�|�I�[����%�vK�u��ul"�+�oI���_�3M7~���h���z����pΕn㭗�;�0-~,ϊ�õA�*+�R��+2p"�Sx��Z!���&��ܱz �I^-�mS��Y�P�r�0fw�e�K	e��w<�x�7=��0^��;(�����ۂ���^V`"{�/�rw%?dx �'T���,G���0�˷�o�j�8!�CfHA�Z6�U���:�lM����e!l�^:؂4<�Θ�����k�����m�FH��k3��B`]ā��\pq���fK��DQ'���ģd�P����KZ�H��F�>������{�m���}H���hY,��Չ��u���V�+�W�b�b�w�W��x��s'�	!��\f��!�9�k�ܿK�d������e�L���&��{xos;MS��Nd=�HX����Y� ����P��
�q�x��,w#���~<��@��fƏМJ�tַ��6�V��;��Q'�OG�s8ui^z��L�2M%���:}w�"����i���!9Z˒K�g�C�� b ��uB�>H�<�_�#�����VJ��a�$RH��ƥe¶pc��j��#�ۉ��z���w'�c�����CY�brC�W����l=g&�#�����.�N(�\��HS�ד��,	wS5�|a������t-E�-[��`А���{�%X~V��_�EdP���K|k��1�6v�Bm�����p��5u?xux���L��/��[�Ea�����3%}y0g�����b�.����'A�>2ApD|=�J�����wȓ��
������:� �:�C9�6`�Y#��\� ��n�-�!Z��v�͝�����]i� ;�M��T�z]�u��r�Q�4�����!՞P)c��Vi�Ae\'�R�0����_��������z�%c�D۶V��|=~]WAw�hf Kyi�/�,��m�ܛI�o`��õ���!�C�=�M(UH��=�� W ���U�)Q�D�\ QTh"!��|�e%4C���R��ckf����DEbpa#M�\�E�ͯ�'�8�i�Z��|�#�z�-�>,���1Y�z��㠦id��Z���q����ꚣ0����ؽ�"RHf�^Xx��� �w܋�	Iy��(�M�3�U�_?`�AǮ�0ֻ�ޥl���˼p��%i���9V�v����8��ْm��w"�ȕ@��7I��.���x�^�vݫT�ߔkn��� ��H��|���F�2g���=��3����U٠���k>�;/@=v��݇�6�hJqq�hu��}@��`/�/�VgT8��.���I���bv@?��5�S S݊	I�!��g��
/P�D�:.��
⻇]��G��{�U�n���+�(�1��MlɅx�*<��Qn�*�G=���'������ ;Y#��p��`p��L�ҽ���W[��!8�sS0�]�+��Xӥ� :Ã�*3Z�����^�'���Y��(��#�o[�p/��?����H6�Mh�Ѵ �'�4���ɲ�D��d[(�qwy�u�����z4Fy�8[.gd���n-o,�Y�Bo�5U^�������-W�g&}�n�N ���C�垌zΌԙ�������=^�?N7d�!�+��^�k���A�F6���Og��}bo13F{0���AR�W� o�U![ӃJxƥl�jQp�3�\t�c@�V�_��߲(	8Q�a[�K �qG���dX�Dbs��EH=~C�M�vTm���?������͇�љ\�I.ǖ�ņ������m�B_	�c�`[wo�e�6x�o�� !Yk����/E^7&o}dw�d���X.�P��5�:A�����B0��wƝ�r�v�at 6�(�I�Y�C�&���`UC0���w�}3oۅ�!���
2�����xA�/�sQ�� j'����ײ)j�@	�=���L]��y�"�j�Ɇǀ�X��[8��cv!$4��6�Ō�r�ႆ辏����R0�"Wū�%�ս�(�RVl�SW&$m���g*
��JE!�J���Z{�5]��Ӊb+	�Tݚ{c3%-A��;Ȓ86�C�9�`&��n�ܧ�8\E�?����2|vՓ�1�46�1�D\�d�߯(�J�Y	��9��&���J�b7�y���/��~�dSqB"+-
ٍt��I7"yV�3��j�5<����Z��Ӱ��}X�����8����GlJQ���� ��ʗy�[�ܽ`j4�]z��|w��u�c�4��l5���!Ο.ERm�Lk�:{���&��X$�6Y�\�kqn|ic����(x��U��Oy*�2���y��h#צD��T�Ty�L��Zj����z����?׿��0x>�&J����Z�@�Ք�y�B% ޳p(����|WV'��Hgb��H���6� ��L^H�e��Y��b�!Ȭ7a)B�d'�����ˑ����r����(qn4|��?�4V�0fU�����R�)9�?ҹ7�jQa�|/���l�t�g�b6���'T�i��-��[�.2��iR�ۏq�U�V�&�PW,���Q����R?=�Uz~���8�B�ں/����=S�'���Z��-����-�Y�,�j_w�vE\�St�
����/�d~�h�z�q>!��!��;���;��ܕ�߀��Q�$oi޶�΄ҍ�$,�� ��uk�sv����"1�xM�����m�1^�9��#�"�ӝ���틋�1�i&u�H}���D�Qvd�~����!�����&v�r�^�X�W�L=e��.B�����R�r�`Փ�߰w`�q�  G��%�XFYĦ�GK���22t4/��G���!
Ӻ�E%�8r��`���2��ڷ�דꫧ��P�~ z?A&K�x��.[����*^w8�����(���1v\�B|���?tiL����!��O(N�����"�zS��+A5�@�g�n������1тr��v����k�m�R!+ 5*���O�`�f(��h�4��{��Ed��-An����
&Wb�̏��>�^.����C��F�=�C����\��g�nW��eM+"�s��}���?�d�s�[�b�W�E� ]r�*�쓦%X�n��	��VY�Ku�d�����R�F�R"��{�\n\��I����L�椝8��|�0����2�/��'2��2�qW�k���,�^l:�/w�G�Pe	�����XDQ�GR���L�az�-����ge%kɓ~�ȿ*K�$3�
���
��/�� J�S���-cY*zAw�"վ�N�A>T����\੼a�\������M�ev�)�D��nU�Q�&5�ë�.�Gb}	�EYN@	���L'�)�'Jp��Ǆ��3�$T%�X7zX��	~Td�����7Kx z)&���J�%j��s�%�;�H��MY��犵9��j�z�6�M���rh�[�@�RfR�%^'�L�Q�啝��&h������۱�7o�b�dB��|��e�U�c�@B;��~.�0�+K \}DF@T=�)�>���9��I�Ąaa����LW�������s��XI�O��O��6�!���ڜ͊$̙�!
��^5*~�h�����I��UƷ�I-ʷ�zW�B�k���}�g�P��$�XɅ� �	�
!���sۺ���e��K�:�āBn�ALRf�.��z��+�"�����K����WJź�ȥ\y?�R$h��T؛8�'3M.L�k�L�}q���~��x>i�����ȷF�^�S��s��3ʎ��u����#�L^���?Y�����FG�b�漖��]b!�N/q~s�0�)��1��b�;$�:O-I�4���L������E��-Qt%�7��!A�>�Ϩ@�>J1���L��*�ծV��0�U��b���Ešv��(p	����Z��h�����X%	���5�bh�"�=<K�enJ�]#�3�;���yL�
rҞ�S�����P��e��L����hh�e���:˞�e4��`��<\1ļ�$��,�*:ß�)�AH,�����	L�[�Of��|`��k&�F#fF����7����]���9د�36:?��S�R���s�bV�f�b,�*��T@��_��Ӧ8?���4�����1(yɜ����$z��	���u���-*��������x��'U����*[0u4����K����j����\v7p�\��u��733����pؐ�Ώ
@k�n&�mQ���0P�};^!A�� D���X����M������ׄ�
H���NUR	�@ ����q����]���A�����:���d��^�TY8��%m���Uk�]/� 	�={8��E����Mp�BM��72�vʕ��[ 4��Q�~j�Fl�O��l�i��Sb�bq�_J7w:<C���k7���!cpV�<on���-���V�����������jCi�waUѫnq���+ۗy��L�?�`ô�J��`Zu���JK剘�e�z8P���T����ct?���,S|��	�������!W��g�_�!�r�r�{CD��\�y�7�<ߑDiE�h�pUèf�s�7 �m����~E��P[N�Z
��6T�5zat�ۼ8;�;7�p����(�(�S*�y�HB������b�=�D�K��/��L����w:�
h�K��N	�I�d���{��%P��	Ƈt�c;'Fց�b��-QS��n�����]�����x:
G
���!*XO˱����B���O
w�������	�Ja�����	<��C�м���1��밎��2$w6�R|���@��z��ft�K$�y��u�tѹkH�+��tug$��X�յ��>Kޟ�'`}ح5 �N����bj�����R,��n�e��R�E�9d��^.ӷꋃqx�%ڐ<��`�"N�5/C�;:y�W��5_�h.�i,�o��6֮
�>I�f�p�`�} H��ޠ���iʞ�O��`M�����B���g��T��g�)ssw�,�k��X)�!�ĩ�jB�{�<�ڒu�t��V�#@�.�tv������5�������s	���a�b�b-^W��������+���R����Z#/p˭���ɞv��R�CU��|�u�
�)����m7R�漹H�"�T�t�i��ܓ1J�^#m��U֖H/,�#ึ_�BZ���P���:�\F�%��~Ia.�N��<�D�^F{�}� O���p�bkՆ���������4C���x��[Y�OX�s�g�G��*�5�����G��5��\D�F�z[�*N%˒-<�a�����@<uxq�p�W�0�4(��V�n3&$ �����ۗ�n ,g����rc��˺R=J�"��.�B�֕w�����)!��)C��0$=AA��vU��V�h�M, ��Bn�C=;ִFSwje�МʪZc. S��$�)E<gi������7�]�:,�S�{f�˪7YMJ�n���猪�͎��K�
���\������oB��9����l�ɿ��.��4%#;���t����v��ŀ������h��sP����t���c�I�/��m�	�~�!�i6H7oO�Y}'�oϗ��X�M3�ŋQ�G��|/�d�����U����=u�Jj壍��,�8
7�4&���|�������.���(�H��L?Xs*�`^�(t��}%A���K��`�# ���}#�����E��yG��{@�"��<j0^�]��?eo$��>�D�t7�V��d	t��������bWM�V�&)��E�Ή a��&�*� %C�%��[��yH�Z7�z�H�A" �OA�"���"�bʹ[�ݚ�����.u��y��%�i�[�"�Z�k�%r�"O�%�W���Ik7�����9d:��>*�o��L4)$�%�x�����)�ɗeV�4�fw}q�љ��%{���fT�����jVnv�����/�,��
�y��Iý%�ea/�/\%�rw��7n�V��M���<z���b,(���a	Xoc�������AZ1�n���K>���a�lA5[�zD����q�@��>a�=m6d��8�(�ρ�6c��p�G�Yv�v��8�{_4֋IJY��F�ʥ��UP��օ����F
�7�-p
~��A������Ͷ�$k�	(�A�:/P�涎�]~����z*�۫�e@���'q2��DL5&����D�z���U+����%>�R�aB"�u�E�!>eO�b�)�)��u���xBBI��$�W�E�������uҾ�������:X_�6nūNS=x���ݭ}��[������U�^GC�	�-smP�
�FO�$��%���\g$�F2���Au�I��s� Ǩt���%Ov(�W�5��{�<��B����(�A!)N����|qցX�ik�W�Y��/�;�
-�^�b	���F5�z��f8��Hq�Ƚ��1��x\F;�J��o�%l�P�z��3Ts��6�����2��cxۨ��ڟ�8���c$Ӓ��=�,�a×ͥ�h����^%�V�Ð���H����X,�����=;�nn{S�)�ǎ���(mg��<��	�>V̀Y��<��$��$=�~�z��K�zW�sٹ�;K��p��~f�B'���V��P�3�vH+r`�?��Խ�4<3|!:�2��b�=�\�N�K�7?PI�#�Đ�%9��py�t�؏J�.,�U}68)-#�/�:����M��v�:�{�������s5��Y�(ʃ=%P�NI���O�������J����N���?�9��`��t��^4�s��r��k���m�����"���h��o��>����E�8W=�]��m1~���R50��΂|+�UE,U��M~]�N%&2����B�-?�<�6vs_[m�d�v�i�H@~�=S��}�������_�6��C�1��ܔG��Bq[R�ן�����t-�y�X���A����r�����3���_�N=N� '����#>��[���ݏg�T%����<	��{����nJ�P��E!�e��>׺/Ч�S��Kv]#3��'e�i���z���Z�B��V���}F�B�Y �*�y���o�� �9UYa�Y� y����=hF+k?�@�ވC%�90:���y��$���{,1p�*�
 b)�#�zy�*��=PԨ���� �S��^:���6z���.}z4��t�)��Ľ�{�5�>D,ww*0�2���g����%}[��WQ��q���d���6�V�*eNxA��EjZ&%�~h�R���1FF��%ZL^��3b�SK����6�CPE�u]3$�~�9ؤ��)$�)���Z�'1��a��E�C�5_չGH 9hm�:�Y�Ҙ�`��iX��b�mAHy4<��$ߖ��j�2��U[3�(����@q6M6��1"�b�i��7��&<���b�����T�9OC����5�y?]v�#(���3�V���ʉwh;���<?FfYI��[4�ci�J�Y|y��T�D-t���h�jej�#�D�e|�&�ӫg	g����r�'6r�~���6�p�5l-�/#�j�_)Kc�xd�eA%���b|�%��ʀC�f�e��xV7Gg�N	�z�P�6�K��,�/�\h\���ڑ͘�#����Zu�z�s$��# �Qq5D���R��� ��4���&ۺo:K�	��0�ĘG�T�[�� 1x�Z��K4q��Ѩ��������(P���k����lA��yt~�ڈ�e:��=��=֡"i�J,G���*e �&��qz{��c�F��̓���^p:	����د��X���_@���6��=���w��.�m&�����9A!>��mT�g6�Z+f���q��)����7R��U�@���?����ٹV(3��CŌ�OW�l��N!p��]���BȞ�R(��GG{Q��97e�@��:���"�m9�Zߋ!�s�
�����D�g��\tr�
������*1~1=�J	c��U3��+���V�,��4���ʖ9���!�d7�8ٔ��+F�t>"w��ꪣ
��$��zK�$��MVh��ϵ��l�N��s4�����É9%��꠿&T9�S2��j��-R�E���^H��J��Ѡ�Ĥ@�@����h.�bdhc�7FX�ôvM�U�������6�ǊaP\*�����Qҝ�{�$dh���Tk�;��b��mob�H��A�^PXr\̳I���T���#��lf�-��Vso��0~Uw,�ZI_L�f��F��ڇM6��fVw{����34ƌ�̽�c.���gzwBت�pGś�3�QK��23Y�'Y?-��o�}�����H����,�|��6+��<���%d[-#��Ѳ��Cx�`O\���ń�H�2�WI"ްatO��3�(�z+�kA�ߧ��E1<�=�Fm�J)��;�Z��Ѹ��F�W�ȓX`ża�d��bK)=_w�Χ����<գ�~3>�6�UDKsS�w������#�Vϳp�>�9C7r�91@���0�]N9�����/K���&M��\�:�31��]�{��y?�0�Үt�P�[�Pa=89V_`�<�/�둆JS���H�
�l�i�7����՛�c=:r���T��{�|+���_r��[�<�Gc�p�w��f�TXOluG��T �!�Mz=�Y�9�%���.-@26�e| ���m�f���]u��ps�^���w�B���.�	�(�a�{w�i�	��+i�y#Z�t-�z��e���������ĭ�t�W� �x��>��U*�eB����Ox�Vg�s0��$Z�.�T��/�F-���-a�-���wm��W�~y�<n��t&�����r[�~��G|.���b?JK�iU#�
��M���rb:�)[j�7$�t%q��=�;�o�!*οi�C\��>:�d����eUy�t�=a_�N�GO�p룲z)Q����ZE�**�Q���^u[/�[d���L S}nF3˩��>�o��������׵w�4���!���m��jdӊq����N�EO��t�g3*���hF��_KM4�A�:#��R��+6 �߲��P���,>���;�טAz���h�Q���ɫʙBu���Z/� ��fL�=�GJ92�)S��!�#~S�np���y�����0y:�n��v�����^��EZ>��0 蠴��#���;;�Sã�K�U��R빺ӵL$��Tm|OI���O���|�p��R��������I�KD���:�c<Y�W@���h��������7;���UPd��<��%�BXv�ͮ'K{{fi�����!�vD-��"�.A ��� �~�fi{uBB}LfOS�d���_�(��͠ ��if���{22�������T��ej+GdT���53��gz2v�s���x����Spղ���<fz�4�:]m�`5��&��]\!W��KO��h���XMVqg��;��~����+�6 �g��6=�Q_�d��+�Ts嵞��Zү#b8�sJ
�(�v���J���d����$u9a���s����u�|L�'�9���p�Is��<�u��]Bsc5p9�n��S�u��V*��4��a��gi��ʠ]_叉��/��.��sv����oTf�4@IM1#&<���N$9#֢B�`��ɇP��R<���C}�������~ ��z��p p-���~抂 ���ֿ���;�Njg�ְ��*�W6���&�nZөU�Q�90U�ZA�D^�Qd��I�9o�7FD�荊aa@�me��	]sw�,!��]����&D{?�IL��;_��A�ڒ91\��83���@M���Jy���"���3��*�`�T�s��Ֆ%� ]�kh�U�9�W��ی���� Uzb�]�c�a���C��G%���`�7_%�^������-�Ǝ��E�X��l�fy��W��z��¯h�e`��QNu��w�|@/��z�X麟-ˬ�=���:d��^3�j�!o�	�ǥ-�%�e�Z�,]mE�r�� &lz;J�@
F�$�I��R�n��u;s3T���X󷐫-M�e2NMjex4,���@{�8V�.{�Ͱ;'uNF���Ⱥ�|%�z��ӜB��E�J�Ʒ�@�M�@��m����ìʰ>��0��G���E�x$5��taU�-z�(���S�|��m>�ZvvZ�	l�g�DֶЊ��.�6QȨQ���2�Rå��Cnc�`ܔe��JK�]w>[Z������{Ԯ��cʗ���ܜI��)��T�mB��n�g��)>�B�@�"c���#O�Y�@Za3xK@2e��vGSGB+p��G���\4t������)���Y���Ewm�5Ƣ�|�V����٦�� �8w�b[�<�I�:}%����l9����ɽ [�".y�ޯ�$�_[�ҹ5���ڂ�q�0_έ��~�[��D!�-7\~7�G$@0gO0j��a7Hl��j*�qz���T8RG p��:�Ndu���~o?����4֠�n��o�̢v�Z�Q�	�M��h�8�I�G���8K[9R�}��C6���&8�8�w�,o�/v�lP��u��aܷZ�vz��M=���[R�\76b����r�*L�!sT	�|n}����!a��\�U�;������,ŉ��0���󞵳��0	*`�.R�LK�gi@P�H9�2���>;�x�p3�^�p T�íU]L��UD�M�.���a�Iu��ղm$
8a;j���ܨ�9�rj��&��[Cw�Cl0+�k|!��QOX��^����2'2�%�mLW����=��9�c\X*[���YU�(O��ݩk�lwҟ��ȷ��SB�%b�Q
�pr���p'��W���QB��`���S.�m���COqX/d�uU�{h@�V�K�?�<�a��o�*��&�iWaƎY�4USN��僌�N�:���\�7�F�} ]Qsy}n�K�U���	��'�!�K�_ϰe�����8�+��uM�K�!���=�����zifz�	���iP	V<���闳8�^�?w�D3��G�����8/x��P�S���m���1�����~�My�jQ���t�K"(z���@�q�7j��qY�@*k�Y.dق�n�-��h �7B��gҁ��/p�,Ity4��mD���C5�=Lj0*�zh���?��7�ܶɟ�W��0.~J���v"z��<� �S�?���n�VC���C��a�8�����F���bG�
4�b��ݷb��ђU!>ZSL�h�g�`ܨ��'`ܠ��řŴ�h�x-4KB��E�:H��Fk�?��h�|<�Uo{xE��.����Vg�#\�HNY��֗ã�� !���ߔ+��?$�f�=��XR��RȬ.d[,^��w��[_}��)+��85�}��{!�F�X�Hz=�x�c<FF���P)�Js#�ᰓ�>��<4&	�!F3�ڛ�����G�620��$V 2����}TJlV��w1�����6�ި	�aH�6�w*�*K˼,X���&Z�X���a �C�L���* �÷Z���b���&߮�}G�Ϋ�q��q��]C����'F<����������y7/���̙�l��W#T����.�?#��>��H�w�q��Ww5zk�g�1z�5�h�L�VB����U��l�}!��,R��0ˀ����T��x�˵�w��������L�t�sA�-nt��m�K�Oh&niە��M�6���C<`�"��6�����Bì��ҞM*���V���F@�V��U'�m!��4A��^!8ѻD�9m�x����HE���V�7�1�@��������A��q�zH��-+�W���u�zgkLb�a[x�\��b��x620SO�rޣ��!�5	���+���<�`��^W�[�E(�#K���R�o�z�Χ��G�cH�:^�O��:!F�yl{���M5R���<���˪�h�D�N#���9os9 Q�=�5� ��g)&r۫�'�B��1P;vk��T��@' ~L���8i���m��Z�#�;���;ɾ����YKSsy�}i`T�>`��W��X;Ɛ��f.2rA##f���w筌�()�PLWe g�����!SWS�g���﹂ �x��Ч��h��r��W�+�yل��M�~��,�v3��&�����C����'t�[���:�D��m��XM4�5ǹ:^ߨ'���oM�%��������KnD��y9�ʳ%�m�0��r�.�\�OZxQ�^��"��~0�`��^0���%w�ۨ:����F�����ꘫ��H�O�� )Qy�(�h������Hg:n�z��Yv�@�5Ή�sD��H�����[�O�ުk��2tw��  Zn�7�y>��ކ@�"�n?HI�5�Q[))L�x�(^�����K�&����e���}W��~�>	
�z5�O��O�VB�]�����]�)�9�D�MX�x�3�ѥ��7S\z��C�J�z1
�[���� 'yCZ���n>���=Қ�����Z�H�f&�bƟ~e�w���gv�{	�[N{C\�Q�p<��^;�[բ����7�������T1 �U���u�W��=Slڶx���X�G%r�y˯���N�.�<�O�[���L0����ܲ����Ը3����N^�Gv^p�@��@ێ�/\���p���J���nB[��(m���Ev\�#����錊��$�!j�b�D�Y���������/�e` #ھ_ߌ~�JL���_v���7LY��:��8��a�J'���n��]B���j�
GjP-�:���۔�򢶩��ִ~�Yx@D$���0��S���D����]N�������p�m�k�d�Q{M�ƪ�ɘ���5�9ϰf��M�V�@"��B�b��w�۞JC�M�l�"��*=�K?@n���*�~�ݽNbo�?����*��(4��T��c�	@��7�(N�^fe�(���'�F�RЍ�I>���YߦY�DJqgd8�p�
#f�H���&=�QgV
��O���fmp��* R��8��&n+���+��W^	;k��xq(����c������P��|�a���-VGll�2��C>(�9�;rm-�bj��S[a�,��D�����y��.`���At���N�� ��/��'�'V���s�zN�5B~��xa����L����=<T"�,,t�%Z��Wl�����8�|<���|�i����%Yĕ:$Z�|��&�+��ѿ�yi��	A�(��4�Pb[����ዟ�H.Qu>��1a6Ga�z�#�?���g�>��,82r�`�'m�Kk�����q6I|3�>�]�ÑW���K����(j&�ơ�l�*�H��b{��P$���0!x<^�c�
���_������SE1*�GS���ؕ���㚫�݋0���]�5-�w6����17�9p���m�~[��~n,�P���
��5AY�`�f�6�f�{���k|��J�_�@<��Z~��ר���͵�B�֯ڪ��4VLМ�g��#U3d1�E2c/у�p���/���I5�z/��:��c-�_j��6��q!dϖ��!r$���t�<i���.N����随��f�b�Z��ta�i([��V}PHv�d���cd