��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���2�U�z�[B`�#�� 3�����E��R�=R��1��TH�G��N�����` �۠���<q��c}�޼Y%�(�"�sڙ�AӛXG�{|��AT��x�PL(�]������r�@�h=n�O�^����	�{K�*�q�a�T�FV���:`��Q�օ�H�m�Z<A�=p�Y3������ϭ�;�jHz�#D(-������Γ�Qk��c����{p������y�q�K�Ʌ&�o՗Vy��P�N�*��}f�G��g��&�W��$�R
����a��㯅�Z^<9:�G��S�kUZ($�%��]&�A��Q_�+�\�~�4�Z�:��iI��`I���E�G�&d;���;u�A���|����"n���П�d��D��+Bӏ�}��r4:җ��	���OR�|�t����֙�;Ԑ������j���3Ң��V�iw
����G�u������Ax�:^Wa��U�7�w�٘����܍TS	%(��!���A/�C�mD7�S�/˭n�7���f�N%I�8�z� Frw�Nêp���Rm��{�����OL��t��:�K�d���d��xC5	V��
�+����,[+�ZLz�ݹ�1�Ђ��d- ͇e���<Ph����XeH_xȱ�+NM#�n�%e�u�Bq};{��I������m�w���� � ���T;�GI3?1��T
�3�(�c�'5���lX T7-����ٺ��̝Ixb�xݛ>!g@OY<?��X`�cߗPTf�$D��I�e��z\�@��~ڜ���HfT"���*Rn�r!�9_e�:-�>�����ekLRe�dό��O�ԧ�P� Y<�y��������~"�(��������QU>%����O�zp��p�������uu�Q��e1��	��ºRq[TU�o��Za���GWy���:���MbF���|)�bݫ�ϵ��pf���qUN�6i���6�KOH������]����ì��ʧ�&���Qv.�1��x�S������(�n�?z[Ha�����BV�(Z��?"���b�c��^»r��q <��	W��̽՛��{v@r��g9������;`�t����Y�Y)���F��wc�	>	9�D˳�'�H9����c����UE����{$���/L�W_�G���v����}��ޤ�Z��z�)��IgАA�sWN���Ȯ>�]� f.\H����w�K�j��O��p�	
5f��x��Gb]嫎���aV���,QG�+��j�F��H/��t=E�e ��5��/����cU9�:����h�W� �̏��^���Z�s΢�J�<�����l_��&4�A��׼|ld����X�#���f�Ζ.MB�s�kj�����η��Q��װnm��}T�x3�e���g�Y%az�5��G�X:al�o߲�"��=,��<c\�R�B�6~����63ޞH���Z��k�6�s�	�e�~�1򨣣�oeB�$�)���r�5���&�zp4|i0��;\�+����x�R�fh��jm����L��E��8Iz�`��!<>C�x1�������}��Z���-�b�A�I��q	����A�q�W�9��g��e�hp��&�=�]2�K�{��1`��4���ޜ�������}2s��٪�&����)�9t�fF-��⨖�Ƣds�C�J;���Ҳ���'�y_t?����0�%#!�����U����/�u#K�����w��n���m"$�����������+��IYQ��f~�|����U�l/�(��zV�n�:X��Nt����mc3�@ʂ�Ј�*�#�>�^U�/��CqyՄu��!�d�w)�О؞��Ú�����0�^�U�??�Gvy|�����c�e.�{Vt։���ÿ���v�Mߡv8�8Ƕq`I0y�n5sn���P*�N�:�kgn\I:�g|~��5�D�^��5� ��.(��Y� b��uh�c���6�y0���e�q�&P"	��Mi�3�	H���H
S�ͱ�D��"�?��o-I3ܝ=U^a��%���6�0W[	}3whY1��m��Ȯ�82�x����
<���rMp�6n���~a�	��Y1ϻS9^`�t |:i*V�qފt��+Xm�=�
p5����M))��-�����#��~�Ε��t��e��꿗�.la������y:�K�VƷ���,%q�I��\^�d�je�s�"H������n�o+�ӽ�5���ՙ�b]�K; ���8����-�l�:�~lӅ_,�
N�6�G#�ph�ƪ4�?�mn�*��=��;�W�/F��7A�ڈ�T_��w��ȧQ���o���}��T�}X�hW�u5���x��T�:Fe{	�q���~Z��Je��s�<Bu��y�A���L��1�i�jq�_�v~���(�zށ�FR��,��0�$a��m����$?��B�*���7�d��J�g�ZPxخMI��iìѹ�fG�6��Η޸�PXvl����]�yD9���GK���DB�k/�"�vr�Я�vi���13��1 5��l��z�9rh]��u��Wxnu�T�3��y��/�6E�%>lM��i�^���ڪ7y��RXZ�3f�v�݋��N,�*E�U�����l&?�q�e1@$+ʥ�F+�D��Mz�`��W0M�S���~�d��4�C���5CW�@nW���;���R�z��ә�y��( M�⎂�ɝVe0��Q�6u�a�8a��S�b�t�ܵ�r嬚G���Pq�FI����� 6�{4X�
�#���Xv	��j0����]��GP������GbNؓ�ƞ�xe3q�
���W3�!EGI��&�^L��-6�o.Y8��OC]�V���f�L8�wó����[�1A���M���	���1"��	_����ĮD��>�&%|�ͭ�*�;�Q��d�1-%J<{�)���M��
e���Y��������Nͭ
/$W��|Eۡ���z�IXX�����0@��"#\�u�J�Yu
������g�$Z���YŞ�T�/��%n�hM��L��xKJ��x��
`�,Г��M?��T�'�R�"h6�ѡ/��Y�ڋk,*Y��D��ӑ[��y�⦱�;hgKjA�ĕ�50X�KC7�P*�'��Kc�ఢ��(>��� �d���'�sw�
;�Hqr��s�I��b�Mc��jd	'G`I<v�5͝810]H���{�,֎�M(����g;G�7dm� \Sf��, 󃹰Z0m,�XCw&zs;t�Ǿ[�}�'�D̚�eL���E�4w��)M�^w'v����񦿠���Bmz CO%�e�Ґ�&x>̶��ʉ�ó�6N�"�b������v��zV޸h$���3��_�~d bq��{C�+��.��A��}���&��nn�k��r���aU��8q��D���ɲۆb/\k��/]��l�}CYȖ@ö�\������B�-��D�%�c�7���5�R+`+Єp��K���c��(�}c�1�
����s�;�DM��2ɹ�Ş�M;��K��)��>/H+�)���7��|'�E" D���^������%[t17C���������0��d
�G��4?EY2�Qd~?�g5n�ۙv�=�4�~F��\[(�(�;�Y	<rBYM4ЄÌE`",/ڿ���e�3���!�K&#pX�5�����r,��X.�#���W�^h3 #L}�
u�7�p0�_O�Q�c|��a����fA�/K���٤��4�Z@E"6c:�����<�a�z@찐1!L�^+�\E7��x�B�{��8h�>�}�J�Gm��؁Z9�H�i���gw�{��z�HK��?�� �gO:�zr�@<Z������G��=�VE��A2]vVU���^�<��
�����ks���J+�������iE+&BC�ą�����;���>�Ov�c�������Y�A]?W]K���4f�z�}6SB̕H	Y���gDYd�+&�9������%��*���A�a���8.W��J���D��eS~�W�է�3�i�GosS'�
��w_��+hH��"#�� r�Uv_��v��%[J%����1\�]t��b��!5.��R�I4�O����ZXH�ld�Z�iu�<�z�J�Z�}&٭�p!����n��T&0�s�����L�_��η����םޒ�tW�����U�)A-��(R~��74W9o*�� ��������s^��dΜề֡�|�+���w*��m�\�Y����#��@E:�8?�P�S�G&�jɈ�Q���ثOGb3.��5�^2j�h�����D���ҽ�*���:b���B��S�42#���P�w���e_��߶����V��Y���7�'0(��<���Cߚ�+��K�Q'��[����tK׳�QlYvΔ&���\ٖmE�^n��D2�&�r ��tv!��,j��m��t�4 ZK�%��V�RJ��*�
'��^��z�j+�x��k{g�k/u�f��x9��"�����W.�c4�LWB�3�tY�AR_��(�Ζ������_?~q>L�UR�\���]P�mWD%��Wg?3,�Es^�������п�})���+���p��XxID;d��SG;j�8(mYLO�<,28�3ϝ+'0o!|�O�fr_L�7>��O��yuR/2�0��'�"z(�Ej��m���	��c�ε�ɋ�+���XU�Ph�="?M�b��}��Ē��`��%��ݘe�e���3�߭wYE/@c����9�������� �?��>��\���4���͔����7���izBJ��=�bMp*3V~3�_h>��+����L���Ɛz�PJ�M�:���6� �bD�k5)���b�OZ��f�E��t�4I��#�4��W����;�e@ei��Q�Q�m��&�K���js��^u�Ͱ��>J����#���`+�`�-��z���7֨$䢉o-��#O��>C�ވr���:\C;�U�c'�0w�O9,�O�o6�"�3H_f�n�-In�q�ڶ�/���k���{b�ktbY�ކ4Ĥ����3+���be Wf�C{���3�K�$�{��:9�h�R�J��#2u�ֈXc��g�X��;��m>��ALK9޺��j�x�vܐ[|ɦ}s���E��B���k��<����cC��q�Z�
�����/Z|(%��t�l�� �%*F�ҁ��X�gz�2!��N��y�H�ˋ�\���t-|��oP�g �Or8�/��c�AHHTH��K���;!3Ty� F	�AK�:O/7�߁�� W�ɔ�^��(�^�\%�wŐMYr��pʏrbϮ/2�1�	��MA�G+�9�+�:��N)HC��s$`�"��҄z�۪_�Py�Q]Z��qZ��
!����^W./2�c�P��%~��E��d�K�.x��d����S.�BP�ϰ��h�N�a)�n�ޤ�L-�r(���Nơ��/A����3��G���{��M�f�o]��N���ʠۙ\����1IuDV��e!k2.j��_�tJ�y��˴ fΔ��~D�oL��]���i9�2��׈��.�`t�#O3��۹Ѩ_e���ׯX1~c2�Q6�B�E��f����z1TqNdX��
�l�@���H&���~H��ڗ�W\�'}<
����k��z��+�/��m��m��\��^U'��8��$��$�-׉�D��:�)���+�Q��)�3,T���Q��
؋�lz��ú�m'��r�ĝ��|�C�a+_q� w��8m"������Q��!L�Q�3�ޟA���ko>y������|4������N����k��c�Hۉ�95���B*��}㣁��/��[��,!F-K���,���R3���f����hܤ�{��}V&�����X::?c��."�]�].k����雋����Sq����6���}b/ଷ0��-}X���ɉ�4;�w�D�ےV�S;Ԣp47Xq7(#�����$O�Su���.�9��a�{�i{�Z0�m�a�k�B�aT�r��c�<�\��ِ��@*`2A��x���6vIy��b�w%��.�\%)�*r��\�8´ۨ+�oj=����S�4"¸&�J�e������p�I�4~��ɶ�.�B2���:z�|�?����z�(Q�*V8�Bk�yL��p�ܗ�p)zQ�J͆Y0?��������o�ӂ���d�R4U��q��i��ߋGxFMǁU�X�>2�F^c��@q~$�" �m;���Xd񇞄�a�b�+2�Ghu�:;��*�������f�]����Nx�"�4��Z�� ���e�	�ϯ�*'���`{Wa&�k��[�p�
�(0��H����R�)�������[d��^>�(x]�oET�'#W�Mٓ|�{�s�.�,\��'T�z�av���U�1�Ƈעn��&��!�
N����:4� @��}���~���s<��F��4&�4d�L4T�m�0�M� �0�/�p��eg�u��:��O(��0s=&՝�k�J���>��Eϧ��5�q��۽rR��4lwC;��׳��:�zpώ��D�!h�E���Rx��UB����[I5��{������<�Δ�Xt(�աUĊ��Q�!S�/�L�i��͒��$/J蜎;�5�M�����!-�0�R��ZT�p~uwW��2�����ŏ�)iw����st����d%�s�I�Ϸ����������)-`�<Y����O(�py�](U���\/ˮb�ʴ�����OW��έ��ӣ��k؆Ys̉�o�Q�$~�G# �+0o���;s���Q�P�s1��-�ևBD�-��uԓf�n�,�6['յÑ�0�pO��DH$=���2Q��Q!)�`x��44��ƃ�m�cS��2I�nWL:F�����#�LE�ٺ2��8�x�@H��wuzo2C�{�*�с�#��k���O����`�%�x��c��k��A�d���@���$���B*�x�ju�����	}�!һ�_l#+G��t� ���D'9�]������F���*(�O�����j�qB@�&��U��C�"Kص��Ȁ)���O}�~�N�6@A��dX�`��K�d��]��O���$&��Qؑ��`�k�8���Q���La�����x���+�`i�fW��d�g���8�ܽ8�߳~�%'�lm�⨑t�H }�R�!b�iV�(0�v8:�elbJ ���k<Y��w_;��KoQ-�!ͳ���W@��к��?��@B������܊���=>���|8��:��g���=�I�����ܐ�Xߦ�,��VFݛId%����䳱�&Ê>.�t�:�ȍ/$j*0 ��c)�E���cv5]�\�`ɕ������N$Vqn�.T0��3�w��kG�a�����Z޻�*o#���Ld�O���lC�Χْ}�-o�"M�OҠB��j<s��-_ �^�6�Z�wp�̶�3qq����H'���b�D��(lg �41:Qrx����p�EE%�)��`��]�4���E4�=`Ա�Y���,�,�����a�Q�LV�|���-T��F���&B�E��8�o��4X&�؆����L���geus^�N��@���k|� 2�	�3C1p�� /(|�;I��U�����n�1nQ�YMZ��_ߍNt��(�Ykj]�"٧)���3�i�o,�l�������l�)�w�j�ܰ�9�m:a G���k�ҳe��2�Po0�!7bI���	z����]6S�f
UM�N���A=D&<}�[訨��)�q�g�n����z����L'�15�|����i��߼ܽ,|e��	��i;b�g�*S��Dg�-ua�1�z9��U|�:O�V�#osV�k�41�D���4k>���IT���NTHOS&c�t�͎E�ŧ�J�0�^��s�÷�C�n���[�_k��c.�)�Z(6���B��j@�GQ�7�t]~O��	�n��܀C�?���['n����m�2d�P�ǂ\Fr9o�_��[��������=̙����`�\R�� �Kf:�I��0a�OR���$xӌ��M"T�"�����e��H�Jd�+ӡ)A�VF��USNh�����'s��b��*�,�p7��Iv�+�jh�t0x��yً���J�&�ѩ����گI3��ԁxF�HGPohb`HT��Jh�2Y�4U<`P�l�?��k�� ����j��&�ϤgiYj�h>���K,,C��E�
Ob�noe5w���N(��rE��Vm�[1��{�'�h���I鞗�J}��?������z2Ȏ��|�qy��l$<��R�����:�����"A]�+L��E�'�w����4I���t5���-q�u�ga�+x9jaWb��ѷ �hԌ� +_��`J�w���� �������S*�?��nƊ���&z����J�E�d�j�m[y���X"_��s�/�D�=U R���7k�n��w�s&é!�j��(3{���H����,���&\ݏ[�s0���]��l`�i��2����헂_߶�:0�W-@-r<��y����5%��֢1���mŬ��ӕN���7ex�.d�YCXι�q�B9�p���j@��.�K�'n.*�^]��e���������.��?a>�$�Z�M&�%�v��߱ʅ�1��?�6 "��i�#��Y�7=��VH�Ks7/�ϵi��"&����z$F���j��?��q&q+�(�����#,l��^�6�O;~��|C�c{%��0�~j4��jhXS���~�X״�D���8����i{�/w���m�,����b�Rmt��)8<|Z�/;��/x'm{���ZZ���C����XUV�Qa�|>�ҷ�'��Ċ�u0�9���Ⱦ߾u�H$���zd��a鐁šM�'Tm)ۥ6h�8DF(2y_T0E_T�����}�l7(R˻�~\��蔸���:���.�{��S�ŷ��=Ѥ)�t��&uO�U�2Kˮҡ2O����=�Z>Co�o-���B$��_\u�BnX���TF%�a���!�OF1�8�YH�Rf:W��]��1|�H'��Ш,*�4#�V�F�o	�d:s��gJ��!��&9�����2� �J�Ɨ�ϯm
9Ŀ��jd<�g=H��R-�e�۳�.�j̑դQЀ>?�Y�z�nm�G�{O,�ׅ��~��oX�@3��j�l$���rJ�� ��|��!�5y3Hn9{� �4�im������0Z���Z���c�����N8=��*�-��@��Jh�]�N�E��Ffza����E�Ii��P��e [�J�|�q�ʽ2QHӦ�<��6(������͡�y6�9�]��-��_�d�T�0|1�k ���LO���,F7ώ�!��jc�FE���KX�����b��� ��D�Qz�N�Q���+��4��W�#W����L���L@�����h]J���9�;]�҈*G���9:�a���6@��Đ.$�ZT07�>Wu}���;�=���	��0����e!�mrN�60X%1����������f��{s44C�2���K���Q8
$���㚠X���������[�`9^7u,{q7��jU$��X��A'u��^~��KN��\�b�w�Z{yt[CQ�jujW
W�4�[7Ύq��lo�i��`��P0���qh�X����it��xYyJ� �K6\m�Ŷ!�Pb{�����`��J���x�rqp�r-��Yف\֝Zc�ã{1(�R��YxP4m9:?g3֦$d���+����ۄ~�L�9��J��ԑJ�g���lC�'hl�W��b�Or���&��۟�)��Vj��z��b�6��f�xY�:�t�Q�}��2�E
iv�1���� J��j$7Ր�� ��v<�����8�N}��(X��)�^3Ej�7ȷ5H:���bfe�[����K�t�dFxgs�����ak�Ʉ��� ���ٌ�.?O_L�M�Tax�_���i2��/b[�%q��f��G�bt����\�x r:x���6ܛ��ft���.���W�;�ʏV��5E�%Y��O{l�pG9�$i� ~P���y|�0���^	p��򥩨y� k��o뤛�a�<%'�ᅫ7��y\g[�<�V��?v�庻��1{k����ս'���� ��5�cW��Q�T��M�4L�47z��ŋ :0�@w=s+������ti�f�`xN��_}0����+�|-?���5��񣪆����(߃�U$�%�:?��v�a�R[�P��!�����i�����ړ�j�.��)�S�N�w��rN��Hn��v��8���"��� /�(rQ1Ag�ۑދ���֫���<�K{x�v=[j13Z�%����9���%V�>beg���3M.K��n��xr����)��bZO��=ECŖ��#�.gB38;����v
QA��'��\An�/ ��{��gʔ�\�ٶ��V���&47M�5��Q�ށ�r���`��E�R��B2�ӛL�Ac��gԯ�-ZXưݽa�bKٲ�#���K0.V��LH�n\qC� ψ��:2�P'x&���H���1�\�?)�*G���;jɇH+v�ȻsO�����JM@C߃;�#�UCٲF� #)B�PC��)Mj�|��&��Q_��0E*��a�������*4Ci��1�X�q8o��o6��fQ0��FaB	Y�>:��\�ShC/���q�-LfB����t�/�l��m
�7u�mX I.7X��t�|�m������3Z4E'I;#���Tm}O��c$�.Mɼ�"�Tw�^�<�O=��1*�;��%	K���f[d`ә�D�{����l��G�Z;+�y������.T⨣���8]��E�,x�I��1:y�r�}��=nQY�Y�t��9�s�T)V􀝯��2
�3�V�_���u��(��su-fcPe�H��߸��7�x1���"_�5�%*���?G�q�����>��ۋH^Y$P�\��Z�{x����i�����Љѱ���!4>���\�|���AХtY�����`�h]U���&�_�G��;���bA�]!��|�{�@��[}�!��ώ��h�O�P:�u���t��'I�a�
_�N���3цٝ�t�!9�*M�k���>r;���t���0����L"K�
��I_��Ǫ\2����~���&���G-�]�А���>���N6��l8�&Ad�0���y�wx��\�FXs�_�C���#/�@�J�l�][���z�!���d�D�G ��o�uLp�5^��D�{٭k���o��v8�GN0��XX�O��v#8.S�|�΋��7�;$0f�H�oCYAi�ew�?��>��5��"j�c��z���I�����4�ݫV��~Q����D�J�ƂC�$k��l#D��������z���| 3jR��	��W��1T���b�t��<��9�"C�<�s%�6&���3�{dʖa�~$
R�]��H�9�)�Q�!���IWO� Pjr�����{�)x��D�2Z<�s%�ȹ�\4�����t�u��>u>��-�I��-X��{tG�6�(�KK��;[
_��VV+x!/Ղ�mI��K��^ƋqɆ3�Td�D�4�Ĝ�*��f:�.>R�dCm�R��3���SM��˶�3> hlT�����]�MQ$@љ� !�9Ze�A:�z��-��T2#��gްaH���������������Š)X��M�B���߉�)8�Q>�!�f����)pn���\��g���6�A�Mi�r�ո�������Z��P)v߉|�J��N�K���"��)�W֚�aV���B6�!�E�q��	�A@���]¡<��G��~��!��?�k�?�N0��X��*W����k�+�	��*(,8i,&��n]����S�~��:H�׳z.���+�y+݈M��i��8A5�������vVͭ���xYu.�O;e�����H��V���s�>E%;K��8xc��X1%<�������f��G�3�v�T����C�\Ì�^�/Y�r�t��^sV\���L������OQ��7��'�M9�Haj��#�Ѯ�Dm� ����J>�&�d$�b��D���y{�EA=�R�4�W�N�P_��plBt�407�iYB����Ǥ�����i�#�ymk=�����XU�T���HLҗ�++q�_��B1�W��8d�D�]��j��v8�_��^��iIK[�@�2b��U�'�=V�Hly�cd/�dQ�ĩ�NǇ��H�Y����n#�&%R�PT� 2H��
�^H͇����AW�)�r�t"��/�'@H��w�+�B�Ax�W��S� �m����Q�~�����������(T���zhc��=󶖩HSt�[= Ņ���:��"�e3�m��×�v���������8R�&���)?ѤU�so�p��*�k+/���e��P �p)֧,����tzn}�m�������v5��`~@bj�k�hggI�a��Di�s��R���P�X0rƘ�t���#�r�m��[qjoQN�>Y��5�����z*��Ei�ؕb��KL��m��!5牥�V@��S,��Z}�|�w���H��b�˅6Y��4��k�A��W�N�K_�+{���vN��ΛL?��F�mL��'뜰4Q?�.�1��*;1���^�Kj�|:��#[D��&�g��SL�u8�|em_�%XV�(w߲�"��:�ۀ���� ������cO8���5����I����b<ԖZ`7u�-ڃsT�~�I�s�xEF Q=�
��G�/i����<�f���ɰ��%e"X5p��H��"R(F"S�n�`j�;��r��4�A��3|̾e �N�>Q�z2�}��36"��ڱ�R�L�4���;R��tڬ�c99��i�L�#l��y	
҂ě��a���av����i�Rc�.;KY�q��ߎ�O|Q�Pw�=�/�UFj�b�,��w^.���L-�S[�Z=��e�u�DmԢ"�$S�8 ����y��?�S�#� ��Я�7͘_#��e��]�a�A:����Zy��I;��1�X��Q��V����E�X���<��.�%͠�V@��4�C���BKS ~(s2�u� ���ғWA-$��~��W�g�)E��̿�'{g�	���\p���z�Vː����O,���d��,fP0b�j* wڹ}��\I��Bc�غǘ�� 8���۫
�5�ht-®D���'vWx��v
e��W��1�A�
O��%n�5�;�'!?�*�փ�b��j�	:_��	�'뷮�<@��(?x#�\���I�?�Jáҷ��gΤEð�Yΐ���H��}%�
PF��\�`/��2��� ��G��XW샸�A'��0�������&x���uVw�?[� ���c�w�1-��p��?7�W�Q�Wp~O�_ ��K�\k�X�Jd3(��b��q~ڢ2�O__��si=����_�4"[[������ÃfZ��N;Y�&��ugr��bDJ�	��y�F��{�������pyH�&�Q��`�Y���:c���
��� fH�*f����`�?��8#�� &�+o�S�Xr�4WB�M�]�N����O,�͆?tN^�k����e�mb/�����K�p�Ʒt�Ѱ�Xĥ�z�.���"�i+�pXC����Dha�#w���*�;m�tP�#��y[�F�.s1��Rt��a��Ti6;�,5P�4h��J<t�GΕ_�)5��ok����?�C��Ǎ7W�IǓ�|�G&dHn���ڔ
a�֭�."04/d!4�+\/�" g�P$�4z���hO�q���]7Ĕ�/ӟ�@'fA~ͽ�A'��)���*�,�?��Z�Á�1�K�I��<�ly�������Lʓ�NT5 �tz�}҄u��&�{4�N9�&p0I�#8�Q�hg	cbڽ�Kv ֨�� H�w��
�pjQ���z�99��/�򖛺[�c��̓^pS�z*�5BZ��Ơ�C�ԇq5.�� �g�|�]��T�L<���<ꗄ����-�3�Ջ����v���+5�IJ����������*�툊86����s��yo]�]4�8�n���v�����V�L�����3n#
�9�����:uNA-�P_�l���\�AH_���|��1pE'*����ABX���	�zX��+ޙ�a&x5�������/c��M�ά�'�z�
��S O��lBb⽶̚��_����<ʜ��Ċ`��7�2{k�S���P�C�:<�u���b����"�y�xR�iH\��C/�4

"`��6�c~��dD�h	��W�W{��P3�Cs����Q����R�F�'s>Io�9Q(�VYɦܸ����M�|�5D.6��"���ǆn�A�mV�Ov���E&~{n� �p�X��Pe^_���0)���z����\i�~��%����}��כ�D���.�~�Ц�Ҡэu[8D��ԁH6|ˌ��O;w�;,��λ��DIc�".���<x�q�k�}y����߱R������$h=3G�i	�E�㫖���^��ո
$L�؂u��:5�+3�tJ���>MV>��@&�â��;�v�Q�9�e�����4���y�Іk*
̽�d<B�O���5�7����yR֣�L�$�;9 Ib��s�)�۵���#��'1EK��|�dCG%G��]>���#�*bO9��-n�W'�A>�����فɲ ]%h��z>
X��.�:'�@������i� �(�&'�0[z�R�Qʘk�m܇��3E�썺WP_�P1.�	�ɧWG�}�l�-�.b���� �?k���������L߁Kk��_5t���bP)�=�/����u�T"���p�kE/Mե����X��|�3j����uo���P�z\\��b.
o�X#qrq�T�"�@�Ю�Y�f�|��.l��!�:�ɿ-?�6�:@xׇ��pO��Q��߻ym��)R��Ҝn=Ax&;������9ȷ���u'�|+���p;�}��d�r��l֕��<���qeWp�3�Կ�Vd�F^��B���]��G�3��QD�K�l����a�-���j�W; ߺO@m��B�ٝ[���E������b\��6i�0�;�a�?�{�a߃�Y�Na��C#���F�C��0�=�
�?k�a��a\a���T���T7<��4j���fr\���/,�{����}��!9�5ßt9�����C�X����>��A�,QO��<Q��m��D"N�U�?�+c�Wt��\�	�!e?I��+�;�[����;5�m����v�S�X�1�Rb�����|�P�}�7q��Wr���H�M��+�v��$�#�ɦ��ؖW6Ap����:�a,�! JQ!;RHZf�*�7�GoV' =y0�I+�xQ���rHS\+�C�W��%�Sl���lZ��{�����3z���;��*%�>��`���I�k<Ai!�o<��}�/g�쾙_3SH	v�i�M*{��l:!rp�I9�=�X�9+�~O��1�,]�夂e��r�[��E����LN���>�cD7����!WM�(/�oI.ag�4[���@�BR���te*�NE�M6�р����p�n3ۛ,l�)��
�Z��%/L��0�b��i}���R�/6���Tu�U8���]Ri�g����0r7s�诐{��'E�X�ص�>.�5�a/���~{u�e3.�hRN[���m���(Wb�<W�p���B�Q�B�j�(�G)�闅4❝����Y�E���$�=0��8���O�S��I(AB�^��ݥo-�l1�U�L
�t<q��,tk�m5��dN��	�Ҝ�?2aN8��W��-��8�?c8���wIt��G$�1>�`m&C.�r�)��1��w��f�b^N�ַ� �ǋ@��4���9�)�M[�@����C$��v̏�}K��ed#����Еm���nY}ͥ'q#�圗Hw�J� ���0��הNa8�!��d�����혒:m�QO%����kVN7`埁�r��&��z�o���_Ӷ�0ֹ��H�,����=���-�ni��G軋��rr)�0�(����,�*q������ĥI����] �~H�U��72��9�<][�����=��*ޥ �;��v�]�"��q)�~ɪb�*�u4���BX�u�K6TH��X�r
���K�%%'މ�WTy�ڧF�-��|	��L�q��;�w�*�����m���C�BT��R�\T�x�r��R����t��Z�B��'Hi�Z	%�!*�}�����bBt����Q�Ǐ��d�z�;��Y��)7�oFKkB'[u`Lb�A6D�������^]�=Hv�V%�	M��PJp{�R���ŝ����A�,���D���fx�� �W�`�:�sf��w�1V�I.1�$��n���{���s��ӵ�/�{���q�60��9F���Fj�h�������S�})H���C�h���؆����Zi�����[�>��;/����7��B�����]�-�Lo�m�NbSO<�f�sjl%ߝ�Tt�����w�A��w�ή�01�dy���G��� e��Q�ts�4�d�L�0\$�j����%|;�Ɯr�J:�D�h��w�=J�.ɜ�;�[Dwg�jJ�&��;\y����������G�:�yo�e���y�%�a����v�2�8��
�t��w������Sn��c��~Qf&��2��Uȿ�Ȉ+n��v͐ѡ�j��l��r�WgM��9�j*����a�O��O�!�����a�dIT��h��Rr�:���&�Q4aP��tECQ��|�oR�ư�~�}ؾπKP���Q0S�# �#�[9�<�����M���%�;Ƶ#���=8XV���>��p����F6@C���X�t�Y����g�Q~��#��f��;��H�������u�[|>�<6R�^�`}+q��b%�e�["��FX��y�E�T/at��o�$�]�煾�����-������іl�;wk�)��@̢2'O�+�B�	��t��R��̆��)g���z�4�r���x��Z���v���O f��z
���YT��>F��CӀ��B��[�e�P��T�{2�9W�aB���qs=�:�GFW�>:�'��O��9�/�.� ?O�`C?���!@�Z#��A�M,�U{���:js;oe|p�#c��E�10��t�s	ŉ��J�xl�^/D��!ݿ��͹\k�@.d�Oy�q$�w�ԃz�\U�C�z�V��Y#�_`-@��k^L�a�k�Oı`sP'�f���,�$!e���M_d��k^٣!��ܹN�G��9��j�q6�J�w9٣ k�=��q�s����a�Hq[T�c5,BϸY�Q�[����'�yW�"`���x��+Aݑ��ۋ������F�G���U����J����t�� ��P��;��EP��[��=���fL+H�aAAg���Υ(�T��IؙVbW��t�H�+ηW�*zT@���:�~�����h���ö�;����QU�ڨV�W+b���� ��C!y�U��/I��֦�YC�f�#��Ы�}���X��u"?_��H�.��%cZc��x��Įs�W꺔��-9i������t#�'_3\io�2`/��7�ԁ0Pυ�o�59�f��P��	��Qlv���~��QF5�6�v�S�lgf�*N���:���.�0lp�5�k1o��Є�.����K[�T�2w��L_������#JS%g��&�w���=�U<,�̣�	ս�O�'b=Y�l�R��Y��g/�d�^�N����/��ƴ�� l�Q���څm��ݪ�É�A����-kU�Ve�h}���#{v�/Y�\섎�l��[kMiR"�@�S����W���O��(�ǅQ��G��؟���7j�0��m['�UA���Jc�ҍ���|0�!�v[Vn��cO��&�m8���QN���k�m��艜-bG;��R��8�W��}p�ߔ��]�h���'s�� ��a9}bz ���{'-��G�5ۓ_��D!����H>w��C<b�i`g4�RV����vv�!�a����W�
++UnbR���ZB���Z�P�xj���{!HK����^�"m!���$j�{|�ui.����_A0DG	^�b��7?�x	
6+\�dT2�Y¯��� ѵ|�q���]G�m&�wAb�i�_ �T���h�7�?�8S����3[9�l���R�b�T���Xz,�*k���ٿ���K�(H��-�i���p3��=B����Z-9*9�L��	��;�]���s����\���?ιhG�V�n1�S)Z�n�M,< h��
�xI0��jm��̄2��?ϸ����8hp���)�m���b�f��z�U��:�������@ �|S=Y}2_�N31���S��h�XB7�!�٤��,`ê@���k�C�;P	����!�y}8�!����2�u.㉌ �ۿ5����Նw�/�leV�F�N�l�a��9�Ñx%!\Pg�
�%F{�$�p.��ʾ�8=���*���a��{�o��,$�}����=9��|k��ݜjΈ+b
���"� �Z�h�T����v�`2�-���̍��)UgÕ��x��g���9��Z{k9'&R�#��+��ɿ�%��.�g(�F��94Rg;���������1:�C��p$��ԅG�_�O�E�jt�qt��G�S"�B^(�* ���� ���i�S�z:U�:��[ڵ�q�֏�7����Y�!�ӓ{���禺c4H�=PC���(CFe���B�6�o=)��S���	=��,1�!B��9i��C%��j��L�x5�G���(ɘ�C�d�����,k�-�e��%ɒ�V��Υ�I�@��0�SJQ�K���`f�R��q����Ο�Z�u�E����X9� �:(
l:m�]Y��Mo��ٱ�\��Jܷ�~�kYb$N�:����7�''���Z���쾴2ո�v�~q�!I�uɄoBK?`.����}�����̔e��?�#��NRq�eh
���o#�TG8�oY"�g�ާ�`��B�uU�R�qϒ�(^�M�Ci@��gn6�%)�\6Q򸆀*���}\�_�M,�o.W�? u4�������L�?ť����}�[��u�hiFG�W��5-��)t�����8����G����#���ت.B�O����sɈ���1J�⻺k�M�pA?^h|;�``�d���������خ�|nu5@��߻%{�V�����(�G�H�^��7<�<a�D������[�����5B�t(H}�Zͬ��<U�Bj�g%D��v%<~���
_��d�1C��(����=~2�e��Of��v�v��1N�Т���.HQ��r�����c��j�\��p腯�w����==�K�����Ryḓ��
s
%�/kN��(n���_��;��� ���D��'��==G�o�����vd�D%��D`��k*ϥ?>��� gE���:�=�z����gy��1+T`�M�D�Yn�e^�1�ג�6C�I�=/Dsv���ʍ�����L�u֝��`�o�-!�X�æN��J'*�����f�! <�W!hEb���YS�&s�V��sֆ�,5�/�h ^�G�\`�l3��` =�w:`;3�(���ny�h&�!*��I�!��
� ��6��[�ߦ�LGX�׋�8$l�n�����o�jD�[��~�'-�WSOy(�ɽ�"|Dc	p�2�#/z��?�'r�|zD�s$���Dyʫm�E�����-櫠��3xd��Ln��Of��>t��jf�8u��=8UR���4�֍론昩@m����o3 �A|c����1�����VC�$܎�e� \�鋛aŇ��c�"Ţ;�h��ϕ�<�����w��5��L�����g�gV�AZU��*�d��*��A�Ex��1�bW�A�61۬�W��5<BcM8v I X��0Y?D����9�(��|���Q�Ra u�,�8�N�갇�K<����	�[�c�U]��� A�� 
�E���VY��^--����-����k9���^�4�����>��wBa%��bSH�3�?�i:Y��5J?Q��_J��|�2B����/����I���y���?�S��IԝۙD�^o�P+�j�=9I_�ރ,{
�*,y8�ҩc{���\���C���0f%W>
0Z�`|�8jJ�h�sH@;]�Mu��x\K�L��+(1�G�!;�T��U�d��D1����&����v�/�P������N��-���lB�+^]��q��k�kż��
��8S��>#��JJV���/����j«<Zs�<_� >�"$���j��ֶ�h�!��\_��� d�c��T
�斏����1�Y)� �,�u��^��S~ZZ{-5x�|�!����7ϸk$<tPUrvop=�_D�C�/�ƃ�!�J='�A?�U��f�FE�nE�Y�"�X}ӂ��e����Wx1Cq�}�߷�;�}�m�½�e�^��#o�Xc"��P�6mw��ʰo�#��Aս=$`�|X�y�3��%��9�%צ�v�՘5"�o�w]>�s^�G�t�!�©x�����KU��G�}��m_x�Ty�ne�n5FO�=��~A7ˠk�}a�ʦ��c��|`9��������Wc����M���L��P@h9"U����h��}a��RS[�_a	(Z<��g�_Hق��������vP�P�fL�:�[�^6�:O���G�\�g�ճ~C��>�Nm�t0g���:/�4�#������S���S=��o�]+��4e�h�j>�I�߀F�߻��~�\��c�����a{z� ��d`fp�U�F�������p�Lфa���Jd5@��%h,*`Z���-�L��j�?�c�4|Y*fqԧ��;�r��[���1�c�	�������X��}�me$4eD�?vl�.�LKk�oT�,�����@7n��������m����[@�AB�2�/C�$��^cV���,����?��g����]i�^��YY��D�R]P/���z�s/i�wgE�rf�w�����F�P��sp����'��3
����*'l�,���t��?�|�f�=s�dr�s�Z7��l�d	| x�)��Ob&�b����ۓ���ĕ�P���N;ZȂ�#j��,,A]ʾ�]- ����>w�2�'O͵?ֲǍ�x\���l�+P|w�1X���g���|�-j�p�MCRW���&ݹ	`��S2���`W�F�[���5c��g]�8S-�	]?O2>ת� !w�aBe|o�"¤�g�"}'��7�+��՛��N���Y�g�Z����c�\�r|�)Ӿ�'gL���;�V/1��ޫ�^���7C��1�Өŗ�����:I���=6yd�|��u�G�}��ؖ�!%
fُp綥@"0�0_�cg�k�I�G�@�r��]���0e\��\)���?c��σJ<��H��r�@"�~��+��_y�ɗ�@�A�f��a3�E�Cvx�	��%_���! ��G�sE`C�%��y���#*�u^�C��Nt�(阅�k����a�7;(��f���cG� "����U�
�r�l!_X��cn�H֧�i����-)�(ʤ�H�=u`��m&7�x�����05]��*�]�m���$|(��5s�;t�C˥��4�2��!ەq� 	thfMK������i2~?!QA�X�M�|N>{����]�������R}7e�S#S$�Q�k
����/shd��hZ���a�"�� �w��@A�a0r�E�`A'|�	C%����TfvX����1�I�/�x������*�����uv1|ȒJ�r����Od��g9$%��̯[Au���ݙ�V}+5hdz��IB��M7�V��������}Ǹ×��0�V��p�z�A�j8��/T'N|�)�_����l�
�\�\���{��&|������8���w�y�Y{��S�zݫ7�V�E���?�uD�Me{������h�]�X2�W�ǻٱ�*tg�g�Ѓ����D��f��rm��"OE���L@V!�=��L嚞�ere!��s��mi�[-����+�f�kFӻ��SF��xU�\�v���>�JC_�0}���~'�=�]���[� %,��<�]�@���V�5�_,Fw�ל�̡�a���n�NN��'/�E
�,����Lm�g�hI�ʭ�㞡�~X��l�v���Ȉ�ý�Jŀ�{,�г/Ţ�� ?��o�Ó"�ϴpvn{��]~kd�6�i�#�|������k7����Bk�{l9l���z���1W��-|9��S�����?e�;yg�B�6�=�sV(~��n�,
ѽ`�ư0� �2מ�U���dIk����ᘘU�T%X��Y0'��3�i�=�M1�H�>�6�]�j^i�L��9�c֫r�WcM�@Ck�}늣�Dȝ���;65����٧�d&²�$�[��.nQ��L�rZ��~�m��i��'i��U�튒���e�=��8�|�N>Hr?�Wq�ф%$ۧ:���*�����f���si���T��D����c�-�ć� / ���B�Uw�g�p;�p��(WnR�x�An�p�]��V�f�g�j��$��!�U9���<:��,��[�_B����!�P>R9ۃXv�-��%��J�ث�� Dx��_:�θ'��i�L���~�8�F�Ʌ�x�u�M�]rg} W�?�]���j�?�~;�/� ���4lӊ��j̀�O�ApC��!5�Q��������s�Q���`���ڕ�?���y�g���B���bӖ���K6ҧx���^����Y�ߜ�F)bUHq�s�:���Zm]�8��B�!s
��i�wG5蓘D�"R�(c͑�9�ƨ|�vn�2�����+n��<����|����|���sB�%�A2!$!/.��m?0���k0�o�!�h2���O��YI�w�v��:/+WϏ�>lzu�8�vxU�����k�A����������G�k���mCB� R�E\��,�G`��Z��e�1+Yq��Gl��zk��
;:KI׸M+�Ex���ص�`�}�6���J��K�ҹ�GU��>}�Q�������ڼ{���j���"���l��2���Cd������Xs?�� �!��'�y��񞡐c $�:�Ў��<lh�) s>0���XD�q~���؟�0���ik��r֩BȺ��Z�'���Ѻl�!,"���.G����>9���u9y��ǃ�^=�:<��T�w�S-�X�l�n�O�KM���Ua�L�ӑ�����Y)�B�!yH��F�+�@P��7n���#��ZXԺ�@�kܱ��|M[����R������;�T��(Ƙ��85�a����E��)�>��y�s��6��y�wݯ�7A8Cw��]'yq��R�J�0HMlG�^*�]t�l��`�X�M�葂%F�o�A^�7�{���j2*x�ao/��S�����-gw	�3]R�>��o�jdq��y���V�$Q0�+Q���'x�Ɗ@�`L �]��.�=�:~&踍�A�W>���:�����ʈ����}�<����}S��B�o���F"a�jx�`-�.���B�Հ?�^�/�O�oUѡ��Pv؃W>0$Mf���Q��a'6�/�(6G��"S$�ݴ�f�ˑd���*�4*�	ڸ4��o=�#�
��;�9�/X�_`�^�~P�%��?������rd�o�NHߌ�*fl0�mz���:?b��dƜ�J���0m$���q�z��?�e��͙fM���$�y�3~aN��:)��qa¨�+1i����jw|V���SsDG[���3��-uZ�h��AV�vCʺC�$c��v��d�ˆ�i��b��E/�,O��6�u���=f%0aH��ZJx^��K��C��ؖd�q+#OWy�������c��3j�u$J�c�IO�:��GI0��|�
%�5�
w�撜-�F�[�� A������
ZwS���r�i�y���	���O�+K���46�I�.�5W�B��p�0&�ͮ�r�A�*xW�-+Uc*�g]���,H���p'�ya�/�-�n�76X���C	�y<�l��ӮJj`:����K�$��@����N���(DM�����1k3�Vљ��w	F㕆���yd�=��XR�=O��er۸�Br����Had�ۢ�s��)�	���1�\·4��`X���!�6Y�L��<�SRC&j?��3%���:�u$<�.��E%5�r�C��k%U-�"k�����i�X�^�G�����X�d�O���+6���0�Ť�"��h�}� �n�����&y�]����o�̀>թ3c/��n#��Mϻb�X6�kM@�ü0�ZE�(��U4/M0L�0P���!s��'b�&k\_#�L&� �JZU?��O38ި��}ݡv������%R� .3���3^�2Fe���s5��O�2yT���O	d?�Q!x����IA��>ew�����l����Dj���?�|hbmX6?�mV���Wݎb��� ��t5�?��u�C��n�B;�����e���^E{}2d:�nb#*Bs�>@���K�[�*&�i|��{ﰠ��Wp�[���v_U=�J�����6qDD�_r�a��"w8��7g�mH���߽�T1<������b������ȅ��p>�~=�B��S?:�M�A��.�����t���8Q�KV��^w��L��V!����q������b,N5���{��q��N�f<c�V���Cp����G/����S���ʲ�5���N��!u�k�D�z�2}�V¾��R��"��"�9�չɾ�|�_G�]!8a��p廧��bƌ*�/Al`,#��>ҧk��w5�|D�Ѯ;������Kiq�ǆC��v��S�\k̓�����T5z9iY��P���i�\��V>s�/�� �`�=� j�@%%x�܈y㩽�$;'��("L���w=�^e��"�\��o�|s��7�#�N=I�+o���S�&h�\᪢;D�g�R������ܨ��9,Q��R֮��ɰߦS��vR�ky��t���[��j5��u��9s2�)���F?I��kS��eG#�q����@�c=�㢥3��J>��Q���6#M�9Ƭ�g����{���"ʮ�p�4�Mk_e�X��� �М:M��Y�S�k����B���Z`/�\��83i�x��-��^� #�;Ū������Q�k�kMu/��*-��fe��n�!�C�~�i9̝�eV���^2='4��J�D��RN�b�I�\�mV��� �(Oa�6Jd�<pS}�V+�MY;:l3wd�S�R~�4Js�1�Z}t+7w�x�zH�N
Q�X(��8p���`�� qʟ��+����hV�(�������8�O�[e�8�������L�/%7�N0���h*a����V`?�j��0���NtY����HD�D�4i)=�>�\
<Z��E�Q�7W�1{?�ˣ��Zf3B��18m��x�S�ܭ`� g!\;�PDlo��G!��	��7��J`ׯ�	 �	₃!��R7ax����u�{�L���/���d�(���jٞH����@a��{-�Vu/o�9-�����>�Yڮ �Ɣ�(oe���b�����g���Y;�}@�@p�H{|O<�X��7L�(��"�0�}/�vן��w4K�������T� �9yޞ�rЯc�X����`P`�S�f�| ��0�^�����`��C�^0M��@�_ or�~�Cd�_Ї���Q���2ڶ�sv��
��@�z�9p���E��b����L�� �CL���U�j�j�|�$�ٕ[�8`�4�mf��7d�xB�S���W��g�ֈ�D�]5-�G�&����,�Cx�r�p��C��L���!/*�Y�h�7R��L���H�Z�f��T����ҁ����rֱv�����I@�1}B�vE�@����6�_���I���x�7�[�p����8~GF�)G%��(R�T��?�@?`s��O����Tv�еP���5r�?��sWse��������	�R�K���E��E�`ԇ����m��w!T���5�+ E��s�0�Vw�1����
����|�������~���G��|�>�i�@���R8x�Wri;,^�/��"w��0Cw��>��6/()���z�^m�z�U��?5��7D0C�Qo=�~l�����D(��s^�A�[g �����0���FH���-D���i%���_��_�K�x�E�j��{��v����H�h��J<{�����p����2�r5SH�'��2��U���:0[ſ$�{؆~K�[��G}�O�`��n�NS�Z�K�B����7�̍`�#��??�3V���D��m\����g� ^$5[�5�`���Tl5kݭ��0�H�F���l���;��5*�l�R�ՠY��e�iVK�K����![M��P̜H0�  jߺ�2�8W̶'M�Q�"�m,��sK�3<�E�y]�_��D]TGJH�\4�G0˛.�i���!� �~,�����C��Ʃm�,p|[(��(��ӆc��~�9�Ķ"h'��@�Q�Թ�s3���l��Tőu��{�̩��զ[����纘���w �PTR���k:rz�0=p'QҒ���������d�� V��S�@��2��>e�H���NǣD6�r�#���!ݺA酚�h8V&�y7J�����9W�Q@\F��$5��I�w��`��Xt=v���A�Bv�p�^kl|����%���x#	 6�\ծ��HX��sN�间+��4�T��\�W��"��[`K�������J�m�E���a��u9��9"�K'�{;���^�=�c����9�޺B��3m`�P˩�w�i�F���g�`��(oO�.�����Һ2¿�f����r���+�⶗���@��5�-��"�*�� �~�\|b�	[�?�u�S����C��kP��s4��#�h�/�YI�A[Fe>ξ���H����k`j��wf*5�(��G�Z���sW��՘K�[k��@��B�ϻ�!��e������%����;�ܩ@�K��}�Dki#c�'��d��=��Gv0����
����ɪ��4A�����B�D�bF�0�H3�lk�l�4Z8�(�qT~T0�<����<�zd���vj���}\2h���m�}\f5fP</!s-�Ӹ��'��_�م|S�X>����OKF�Hؖ���޲(���tBx�Q��։�yF;��t޷G`;�御�t̤+7�w_(��XQ+U��ٿ\�	�iXqj��l�&�F)A�E�]~����瘸{�Z}�x�M���� 2��\[�o��U@������)��::�v�a+AӢ��b�T��?�ŀ'֍Όr!<��I�@��{o�y��n��M�rn��ە������槣~_�l[��,�����t.�{���b�3��b�Â�qs�����35���t�2li1�`!u�a,b��ZᓨJ,�C4J3�@>�Җ�'�o������+g+�~}3�.$��R�z��Ь��IǬ�\ĎJ쥍\�3Lש�0"�"�
cWY�#}�l�1��~�X& ��`Q-!��E�wH����2O�4Y����5㔷ӟ2�T����
 ZV�D��=��
����٩IHy��5ԋ����	̍�#O�2+�Z�9X����#�bmRaV�-�Q��(R������M��ּݩ."���:��є��+`S�:M��X�)9�ϰ�r�q_�ۄ\Y(8��@�sT�Z">�W�eǄ�{)+�Q�]��l�A�-��@�>�Z%��m>O�,�P�E����I�l�����-�xSF��TI���@�\�1�o�=� H��M������q�����Q�ad�\q��j��c7�jD[
�Y�%����{�|b�㌰�~�+��	qq{�Tl��B!�6J{����h޻s���G�����'?߼*�H����J�5��e!�k���/@1O�j\/R��#썟A߃p��B��2G��z�xW.�QP�ղ��a��X��;Y�WAncY���ӋW�u�x>����ʚ{�-���7+Q2M�b�%�+��������S��+���{ф��,i�9�x�a����:s{���L8y���Ɋ�1��e�nuh>룵Z9»>g����<�z�4K
��>������q`�����su�M�U\�+'�����)�M�p��Q�?��n8��\�:��y�:��DT�uSH����-;�[���� ��y��؏�&���rx�U"����i�m���\�(��wӏ��aw��{/)����v����yW
�]J�����`�~��|�