��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|8���e5�I��d8<��c~��#�|G�R�~��䣟�"���g��k7�����b8ƻ�a�2���S����%�ۋ��3����|�rV�g��F��[�%�d�N/W�'��##pv��n��y�8B��C�|A(��N�z��?� �JG_֕pkD�&nS�����_�Y(�mWM�zx�o&�`폽V�*�{N�4�'����"Ź�YE�������iH���s��.���K�"6�͙M@if/yWZ�4�.}�(� 1ȸ󫬤G�'�S��K&��T�נ��4WM*	�-�(��f��N;p�"�ϓ��s�@���!��D��X���3�'����I;��ۍ%K	t7SIR�f|�Ŕ��C{�P�dZ6���C��#� �M�5�{�������2�],�m�x3N� G�W~م��f
�*��t��������$�ʵt�� ��D�$�c����1��+�U� r�^�9'�K�^���ژE=��r0��a`-��!���䐳N6���ƛ��0��F�{����Mʌ+w}�q��Pڼ����{a����9��7�L�W �h�oI�͝�$���d(���T���i5�|��ꊕ�Ǆ�Ĕ�lA�ݐ!�n��yz�\�5��n2�ϒM�}�Kn���|M<�s|�Fm̈Q]*
8Ӣe�@$�j��S�̉���4���2��I�S6�:�q��w+@�0@���i��5��/���'	�1��|��~�N����GzToxIB��WTU��6��~]/V[�ڎ:�B1�H8����r�`�pUb�[����$~㊩Sh�d2Q-\jh��*�:�z-���N���,�iS���k�vY�qZ�l�I�?�~��{񅘒��S�H�H��"V*;f�ua㽁Q���!,���%MZ��q@�=��h�bN\UҦ[-�P�ac���v������<n�N�=���_EF4��j���|��!h6H8I����2�LF�ZfC�dp����b�=��H�N+�z��Dl.�c%��E���CGAJ���,�ʖ~�j�uL,��Ec�=�C�mG��ٶ�@M�23���3���Ɇ�X�o[ߞ].R���/�/:[}`=��rms�Kh��C�C@=i�W��OBb��P`�0;� 8A�5�����U "m����%v�D/6����p�[�.3�+�l�����fY�Z*�q���2�i0���,��$��[�����|~Z�5~�pxk+cW��J�_��h
v e"��� c�ƕ}�?�5I�!�ŕv���j�/Q��O���
��?Q��8�$j�O�5whO�����:b׺׬	�_���V�׼#��αM���D����0�����b����j���s��w�J����V�L�@���<J�q0�ضa�F�i�R �g�t�a=��n~XE�o�� ���l`�ء�:�3�v������L�PH��B��0y�PO��KC�=m`j�Jb|0ן�82H$|,#p(�������� �|����l�-^L��������</��ۀ�۲e�YC�#�� z(�з �xG�]�%n�ڧ�oE���u	5h�T��R���H*V�l�8�_J��&�w�� ΰ�$�~���rXVTqK�����d$�"A��M_KP��RfQD�}HKGES��[��1Sa?Ss��턅�^�t�i�x*z�kнe��rC�N�^�ɻ���t�I��F��~��w�݉N��~b�+��Y�=����
�E�1�y
K_1r%M���|��X��q�'|W�G�����Wz��aBz��tD%f�V-����)$��ə����-�L�����dؾ�6~���U�$nJM��'�����e�������Fy��e8�GU?�B]L�@�h\�?R:�ެ�fE�X�s_;3oMt�ϱ������5���M�C����f���"HO�H�_9���9�������$��bkp_�W���� �wo;ޤ _|���`b����[�]!�Ͻ�xJ��uL�֥�(}�ph��Js+&�-h����=�v~x��n3��wZh�>�ܣ�K]��)�w���+3	v?�
j}ky�TM~ظ-6�B>���w��h#���W�偞���I?GS��E:Mp�/��=���3�ںME�|�N�[XJ\Y:�4�S�i���)��L��6qyq��~�f��3��N���!��x���S56���)ZVg�h�('0�r؋\�I0;�^Q�9HOx���T/�8��7�n��D��j��}C��..d8����zoݽRI�W�݊���hȮP�2,%84��S���m^�Wd��?X����N�7���6e]G�R�ZO�r��߭�������r$墨���8$
*�����H;�-x�r��@Z���0��%���*ѕV𽶕(��h=5<�57��E�|�,����P�s����;�9�x)�	���I�'������鏟~{,8;�$�\`p\�H��W��1i��y�4�zw�!u\Ƹc��Hi/F�(fil�%��,�{����B�Y�'ԓ��5Q���;MP���z*h�ZUk�0b�,����@lIT��31�!�Z�l�Ҋ��w��
2֖T٨4���j!���m����X̰�{�p��(&������k����}��I����� vpm{������	-l������)����F'
��"R��3E�D߈Y�;|�`���s=�j�h��?�hA��	�u]��)MfZ*僓5�W-�B�}u_��rd�5a�0�4&�Ո�5�pf2��̩h��W�r��PK�ɠ�����ǌs��Sj�{�9���.n�Z���C�%��< ��B�����S�PX���8˗DU������~4�����d�{���9����r��t='G�����*;��u-9���M|n>�qlݠ=��"ɞ5X�{��@O����I�8VF/.S��\�!�?6�q#j������t>h+-��9�O+SE�a!�{9x
VG%�L�~3�9.� �[o���>�l v����ev �	��頸���.3���FG���[п��3O��m�F�O�B]�r~]ݷ:��RU
����%���J	�o�����7�^���z�x��zl$�*���#���{�C\�C'8�ݭߊ�k��a�K�F�,�N���r7_��T~�C{]�*�WoyaG�ߪN՗d�1�����M��)�8�s�b��?Q�f8�[���1������/����x��o�'ܵ*�L�~�F��)L���޲�_�+�žg�m|�6���� =Ф�N����1��KPc��?�)��:�Uěp�z�q9�&���3�})����r�ի)]4��~�=��%��یfm�e��?� �6����R�����>��%ۄ.j޳E;yx+��  �
B|;�|�'d�֒�/��'�%U��|	��٬wآf�۟�P`O �s����b�< y��&-%�g���!;���j�皭���g !�w	��7�=�7��8�G0��#��}O��)>0J=]�c����Ъ(C��t�$(���
����*�m���'{H�]��=-���rT����t�զ��!["V��_n��$dG**bӂ.W�}�w�&��)Y�٘d�����9L�Om`������&�p@��H��#�Nm4dO(C)��Ꝟ���`;�0I���v*��t�_v΃��_�K��*F�$񒻣p)�vR��5�s[V�@u,��~�%�ʮvZ��n�nK`�ߨ�lGk���Ӌn�����i@u��������T#t�5 �Wrm)w	�*�����3� 
�b���	�1��Z_�es&��F7I&ݧ�:�)!σ#^D`�&&�	��BU��?�q)z�zJ�9m�F��x����.�s���y�����B�V}�}��/����d�6��ȅ<��<6oX��߇��p�UU�w�Q)sN����Ŋ��Ͷ�LL;���bq�W�E�#� �4_�ǽ^}�E��=��nmq�o��wX-���`~��:�J�i�����)�,EٳW x"�ÿ��Ȥ
{9���0$p:��@���$��K-��Hl�u�JS�\ ��(�x�J�x�l���:��H|�4�aK����������b��RF����D̑���zw�Y$z�]�!���^��"��	%H�����8�Pĳ�������?p|�vBU������֚)$�V��]]�W���6Y�l~�%߅Nn��S̨*��n::�1׏r��FрB�lJf��Q�X�jd���B�I�Ԭ��&��`Ɲ;��u퇍~��L5��_�K��[+���r�IL踷�+�LЖ�*K����z��uvxR����C\�ii�l�8���LT]K�Kű1t8�us����@�}s���cyрvR��ů���?£z[��\LK�_���]wK���0��A��ʯ�wwz�.�������K	��1=9�+�&tM؋oi��/U/Ł%?�C�2�����1-p�!>������'�*�[ze�Z��t��ia��z{�6 �oe�"����P,�m;޽`u!�Ň���9s��s�y�*?��t��t��ܭ�v�a���1�g�t�j2�2�Y��w�|!�P!F�I������Y�zSPh��RFPa2>C�ez�T�\?�C7{/��˖��Yۇ�@R�b�+b21�-
g��+P���H�@��&�P/RNv��	�v�*���H{���ER�+A��GZ�J��G���qʸ���С���Ӎa�Š�����5��͜�ѝ�;r�Gw�!�f.��c��3��ۥ!�[H�֟�s���_�ک��6���KG��"kZ���;G�+i�kwK����~E���z�����:����1��*��y�c��rnC��E��YmȊjqh8=Sַ#�G��,I���p�mΐ
@59�=�&-�8��=�.|Rn�B�,�2�,k
��G��b��<MN���N{'�?1�5���P,v'��b�WM�A/Yw|t��S#6*�t�m����,͓�>
��F{^��7�T�_��=oA蔇ɡ�)(�"��b~&�z�E��q��Q� >j��m�@f
����>x�����Z����e6�U�ZRu�.8�_��?"�/�<@��%����^ ��F��H-߂6}T�4��FH������8^1�@vn�ǳ��j�m�[��a����=����v�#��J�>����0�DL��ĪA0��2����gUrC���)���Ys�^Ӂ7�3�Jl�/���./�놝���M&���R���.�W���)0s�����7�yB��v"�j��� �~�˰�凘Yk�O�������_���K{K��3�.�‭�V�Hc/[���MM@���"�re䳱t��R ���������J�x����4��L��OD.~D��t��|�ߣ)/+�wfn��]H,���PN'�Y��́^�Ènl��}·�^��ۂ���L�߻��K?���k�Z�)ߺF�Z���-�]�����{�Z�F� �b�7��!_�<��@��L$:Y<���5�Y�7�>1���9?*`�V�"唱
L�JϺ��[@�	��^uZl����=�e�w-�����5�p��#�v��@e�s��6�~��}ñ���w���a���B1��>�j��[�ٙ8���gDXҮF^tY`�8��b�޸R~��q"r-P�IN)e-�꺅	�ܙ�ib�d���mt�'���l�7$|of-��ȇ�����9�3�wz�%@��P�4'k���>�	�g�J������]Y���C�7]J��N�k��$����Dʫ[#*����6��-|�m�m���Dє{���T�y�Y�곐��Z;v"\�M�&{O9/[YA!�u!2G����	2IY)~��Fk��6�׈�N��I?;g�ӆ�D�H��Z��/�+��}��#*~����rb�����C���s]�B�*�0й����܈�[�}**%5���߀s�!��?���gk_E�c��V7���Z��8�5@R�=w �].��b�3C%ؚ�1o��TI\�{�0���5�j����$J-O�mII �����,�y5�Ӟ�6��`![�uBU�̏(��Yrm��v�n�!Hy�U���P��-d4D���
��DQ�֨���0��������0��Òs�� �ݒ{�R_ڏ-MI��t!Wj�ﴼ�j,!([ڢ�P"�/�.�mR���^vD}��<�`fS��c�lwP��~>E���8�P2S��`Dw�a&���O""*���s��;O<e��W����A0�{FgR�?���o�b��S��E�C�]�1&H	m��^]�tZ,>;�4��.��?O'ry�����
;�o_����|qj�O����.kԝL�c�2��Y�q~N��Ӷ��W��j���fb����"�6�=�g��ע�Wl��O�o���o��Q��ZŊ����5l��'�z������%-F�l^�>�轀����dN:�^��"
yY�D�,��c
�D�UR^��kw��_��:D�e�������\�pl�Ͻ��Z�3�O��M���)�tǖFXW�����#� aU֘9��{3�"�����2��x�>چeD$Wr��{}��:����H���,$��m��jVt��A�9(o@�& �{�����p��2�Ŕ�{ͭD�G&�S�dh-��}�ީ&�`-������)q���� �\G	W�6.kǕ�s��z�#�E��X�̾��y�I��1��S��k�1���ɹp����B4����;�����O�Y�|bq��S�*�펞��t�@��a�)#¯;!wHe"��|���wT��� >F0����*t�=�g�jE�d�Ս"�=(�J��z�'��Ө�$��SOgc5O|/�����E{�NX�%x��ὲ���A^1	�@�$؁���I��o>�''8�c�3��R5Ӥܴ�v@e��/�ŧ�\7C`=���"�.i���L�/��1�����08[��<�k����P4���j/q@,ʳ��{;���j��zC3�U�1k=��)�Q�ѳ�h/��e��tb B��2��b�G�@��'-�� ��� v�e�;���B�*��e�&��|zϾ�N�����E���)��ө�!,���[�f�Ϟ�����ɟ7�(Lv����Z�kP���l�"���CuP`�z�9��4e(��<�&ú���4���R���(���s�o�����*��u9v�S�"Cj��|Ğ����/��v9�z�>��V��3����,��ܥ��������jdN��3fW����O>d�4���8_$$G ��oh�"&����)����.&3�Ø�H�c��yĈ�"2�cV�*+����>;���|H*DJ�˗q�38]wU:�|~g�4*�goB�
O�e��V�G(�o,.!p�9?��\Ѭ�.kK r���|��odz�ކ��R ��T=��f򍅣��J�:3�a\u�Tn�
� Q�o��S���d��6�;R=1�4�*����REq�K�&H4�?��$*Jd/�N������2A�0���lL��N��2A2��q�>�7���*�.��9�c�Do�p�������?#�2{hw�
r7k��3=h�#��'M~�/v�{f�u�F�m; ��t�9�듺��m�q��i�X~^w4�;�M�Xs_�e�ۑxK?n�r�}��6�9��NK��o���U��>IF�m�E�+��jZ������8F(l)T�zR��l��@p+p���Z1m�`��z�}'����0ZJ9�����J5���A~�+�Rƻ�L�8�w��\�`o�9<WDM��]^)�^�Y�6�C ���9�6��I��v���n��Y먆D���93��-�ح��=�@I�7�����m��|J����PZ"^�VN�Б�Pnra����	�KK�g�.p���"}d�chP�ɭ��g��.!��-D5�!5vs��0W�Te\Oq��~u���tN#���bo��{���pK��^�	J֧')��rsE����B}�N���^1 �`�I ��<�re�h�lui�sB�z���π�ۤO&�ָ�Ό;�beه���=���3��b�;L��R|�4�,��ʸͽc�
��{���ܫ\Շ�&�O94a��>Y���Ɓ�D
u�e[xE���ѷ_g���w?c�W�	j�ҧ�X�ւ���4B�Z"��2�����j/B3"̘şg�k�o	�E��GaP|�:���A�W�t7����4�Tg $�C�W��yT^�ߟalG�_��cd�̅���hl�
����#�	��SL(�,�YC���,���>�@S�[\	�ׂOU�ϛѸ�XCgȔ�p+�ߢ����3���b=���~]�u�P�� ͛�T�m��٭�J\���~���Qo�����I�z����,�O��<Θ{H������1nil�tw/,M�Bg�~�HB��T��5��s�l���k(8�tK~J�_G
*��u�%5�A������/8vqP��l�@���/6ʨ�������مvҚ���ay@̻����s�$;,Wަ;��\>3�s�<x��ԕ�J��"l���!Ubā��`����U1��0 �� -�Y�D��m�P�Ê=�� s<A ���
=h*o���f�2!�=�BO���=}a��{�Âv�Cg��;�a�.����]4G(����R�Z���E�%�[�U���������M�n�'�zB4�T{�Q�h
�y6;d�躇�������쐲*��1�O����p�Nr��ץ��}i2*!7
�h'1 g�'h	+�%P����9��X���Àc���s�D�EAc`rMGj�	��%�5u~���e�����wq]��
3{c��CGAo�ë?#�G����w�u�}-ۆeS;�AH���Ɓ�5ńP�}��*������	&	-�oX"Y�� �����2�[w�,��ŴZ(�=����`�7�Q��q�@v�L�m3>�ȩ����d�B�r9�8v��޿A�p}[�K/mR�*-z���?oP�DQ��@qh���)E�`�Y�撞�p\�	���t9�����M�hO�bV����Aǜ&���!
��Q���١��Ъ߅X9�_;���}��4&(ŕ�O��k�y;�]�v�7l�r8���-U��om��9
����@Gm�Z���M��/��AP��wVk v���1q�󥗣���ƅ��p)��\e4����K�R'GV�ư<�G[Ѥ�M��,pR�Ӥ�%�wT��'��6ڌ?2�%���Q�Q�x��շ~�`I�aj�����`çZ��'T4�o�2�  1�"�}��i�Ҡ&4���jE�>���Ɏ�<����W�@I�����G!�t��<�Ky2�n6{ �{��G�{�]u޲���*,;.�1/���1�<~�Z�[;�/� ZK��=h!5حV���J��[qJb�O���2�å�������Lm͑���O���)���>�^4��rW��mn��f>ż�#]��cΝ>�鱵lZ���v��8h�����Ћq��r�lL��'��`Y ��Cf\{xp1�!���l��8|�v�lc��[�ǁ��a����L�z��-�#u��-m($�#���Q����fμ�6�3f����z̮��l��9S
��&�6M��p
Pȼ�qTR��]�Ļ�	
�M��'���9�U\q�y�u���Mj8���r|ua��V��w��UlU���C�g��U��,���ٔ!%�\K��}�&U����1��S�@?>��-ja�5��ݰ.�ק(�09(�Ϟ����D�ί����u��
������>1��uܨ�ޠ(����!�
	؆bU���I1��}�N �f��oaU����?��:^��%���VA�l��A_��Вxݬ�h�q���#>\^Ξ�Mu`맖�x��1���wF	V���ct��o0�Aw'��e�X��(�	����KE`��+�qNcҺ6)�D�p?r�:]��J=�Ø�^7'[@K��T��zb�p:P(g	;Y������ʁ+��)��c;)�R�ٶ�6�����lH�j�MJ`�Ӂ}#��@���|�����$�^��P��<R7���38t&;vN�G�W�ڙy�%fL:Œri��?�Q�W�;�Xz�����zM�
B��Ij���䬱g%� gr�y8��lbM�=H�4&�@��܍�� x�52�tI��-:�O>�hs�܆5��
J�5xެ���&P$�^�~|�JD�}��Uͮ���3�;���!��ڢ;Hde�����|�aj�ۭ5pr3{�#�'n���\�,`����B$M��a�Iխ�!�I���Z���a�J��B��-����j����я�2���
��.oźw���(tކ^^������i8�{�:ps7�pl�f�+�5��K��|K����~�(�X������7��"Н�텀�!:�R|�$g��4�+7V<�;1?�A�r��ȥ_K��L����sK}��_�0p~�N��	wӚ��G�ݵ��ÀҦE�s.�������`<��b�5��L`�u)ai���t��e���`8��v��
���{�4�$9�/�Ӿa�s�������-�i�����#����n�Z�D�ܵK�U�rlBH}M}�S��N>BT�������ŗ	�dp��0.OPV���:Ͼ�@��-�ۋĉ��5T��|��Nn�)�D <����W�X�/y��y���Cb�%��9�wCݓ.	�A¨�����`@	�SG��3À��z!�a�g�߱�L�e���st��w�������<Q�w8س�K׹�����q�F�@���c�Z�?�͒���q5b�T�OvMF��E����s�~��x�x�AchC�<�R�rV��W4����~�?���e��	*����P��Њ�c��,Cĥ	����8����<���8푮���F�9�1��ަ�_���k�BO�Y�ZB��f]K�)�����>�)X�D�H��)�W�㲨;sB��������������G�gb�Ք!I׹�Q"U�����o����Q��NT�ak	��D=��cT���}�'d�Ob���T�<��C͜-T�^?R�P������4�l">��h�%3N�;Q	o�g��oz���\��ƕ����&3;�%�*v�� �8E�?�E�0�Gk�W�7��lSe�*��yki5�����!���b������QfH{�BԳ�><w�{as�����v a������&�H}ރ�B�+���xx��
�C���x^��&3�gM�~�M,aD���(+�۴Ĺ���eʍB�`0^֒��K�!��G��?�wȻ����l��A�h6�/�/�O���U!��l|�X��}5���Z.uD�����Yr��XU� �2�վJ�P��L¡��"cD��F�}�n"��?���(;�z�jTT醥¶�Su��
�R͚U�=�h�l�HB��:��k�j����f���WqUsqc��;df�楂*���2|��[Ww��=b�s '�%ړ�z�WxZƿ�5>��|f����-�(N�C%	V1	��$2/����Ź\w��T}F5�]|���R�I��cj����]�UV����<�ɤ����&�S���)�IHk��ca��.?&oJ�X���`�F]�[�N�Jͫs�0���I1k2�.��͇9^�9���Ki!��R}��9Q�L��f��F�ȧ�IH{\2Y�"�6e�Rt��E��b�V�7���>�kŹ��ʕF��4aJ(oȴܶ1gZb7�ӏ��P11M\����̵}�٦�[�5��M�H�囗�?�Y����GMmR,K��/��V�u�YM����y&gr�}ĕbo�%�J%�r;�V+�s��H!�=��-jwt9P`�_He�B��t�j6�f�I"r ��Ftev�w4��y�7���W@1��U��L����9nE����P�Z����^��8��f�q�ċ��v2��i<*�#��?+�1!���9���u��1�k�?�Q������ ���7P�y�� �Z��;y�u��U�外�v%>s�����Ns��go'α����@��>ۥW9l	<���b���:cc�a}�{*s:��z�b~u�X -��e(V�T�4�Dy���b��,I�����a�8�R�vn�ؚ���M���ѹ��iHi#q�#�Q��[� �)��Ŷ9�+�D�d�5��fi˷�i&L���^<���k��sn4�2��u^�oge.+U���C��Kf�z~�BV�ӿ}��gT�K�b��UUJ��͉2��'��:���J�<�Q�s�g��L/-vʟ%�+���S��oJI��}4�{���d���0���
��S�C��{G�ܝ�d]�n�7��<�U��<�Ȥ�k,j��$q]_�J�/��b�� GD�#�0�]��LY�t��o��l��rP냦�a���/L1�~V?�e��V6���Q:sX�JwXO=�x�E]ؿ�9E 6�QN��\c�k$��jR��2���&$^b�ID#'|Iy���E��n���8m�
��ؤ�Օ�c�>T �m	q����cs�d_��5U�n���Ӣ/o7��M/@�:'�!^p��mH����4j����?���r�c�	J�"k���\B�0��t����������C��}D5\�Hx8��	�:�Qw��'������d�M�eΟ��(Y���h�(�$WF��� �hڊsI�q�]g��z��%��c�T� #�3�'��<R�ȝo��M�/�Ge�s�Y�h��"ikbI<z�z�宋8�L�<6��2u��;Ҵ���诸G+N����G��O|�����.�j�A��l0���:����R� 5��JA��,���{���U��������(�P)��7D��<%]}���4�P�,gO57L�,��w� �IA�>0��0�
`�I^Of���m(�ԃ ��DTy$�Fzg��St�EI|i��r�~��Q���C�8E����t�]�]�-w1MݕN��������>cٗ��}= m��"��ˀ�=J���� ��q��ݔ�8���1���BX�>��vZ�h�)��`���%�����e�M@5���TX���AN~�G�'��Ǿ^qV�崰W�:Z�#f�jt�m����GŤ%�OC���EW*N���E�2R^A�.�k�>��~�]���a�����|v-���^��VY9h�v������!຾�Ix�ڱ���"#(;yQvGz�
N1����11f���Û��(���a�f&�{��ǈ�p�����ë��%2����yjQ�<�PWc��{a�f�3�3���2塃=��D4�i{�R�����*�!���0ꪚV�z����=6���a�B;��t����Ju4�8��dX���@n����O���`�I�SFA��љxp�	�s�[q�·�,������C qԪ�L��*Yh����E��vwU�}=4�h�矼"P,���mˬ��� ֘b|`����>?7HI�
m�c���(��Y|5ޞ�������\�fh�)# ިQJ��� � �h!Ũ*K���$H~�{l������D~Q��(����Ū����(S��k� �XG��z����;@�WG��&�[�`�1��Y�*t@�-�Ϡ|ތ���숻 @��q����NN7��A�\F:2�(Mӆ�S�Y WW��ę�@X1�����I��T}"m4Հ+Ҋ��k�ac��E�.��IE�� ��T�%$���g��w;bm��C�gV��p"A�<��M�U@T�rq!�S��5L1"�������b�JZD|���+]�nơ��\1�7�#�R��e�̻�(G^~����5P�`���,�;����$��	���)��(�4�b���[=�n[,&�.�:UJ/L� G�E�U�+SS�;�H6r�.j�:���S|u�ǿ9�8����+����k{��>��:��-O�%�O>����&>�Ш�ch�xxA�R�>	,����&�,��+�EN��,�ִ��
؉��#��a�ޜi���ͧ0G�*m���#YA|Rw�i�&"74s�����1/YѼ����;���x�����-�:��]{�D��J��˾�;w54��2ޒ��n3 �v&lv��^�^��� �T^tH�	��Lק�A� к���u�_����bUІ@t�|��ڰ�ZWF��,��`FʭZ�P�tKC�B����kv.	��)|�_����2�DA�x�^T�ݳU��St��.���	k��"�o�{��R;)�����B��:�����=����ȑe�!�N�s]���BA��uh�yI:�����}
�ߴ��4���1U�lt]w��ZBY���Ńw��SkO7=J�Lf��Ϸ�7=\� ��S�j9ڢ���Į[@�0D5����T��U���4sqS���-�9e2�g&v��td�s��-�ٿ����~��+����UeX�*,�����3�6$�B��3C���G/O��1��@�h�߅������Bִ>4}b~�3޻xG��i46?���;�W^���Ӛ�D}�|V3^�~���5�����������ַ>~��$���nu�i��<��`?E�� B�C
o{��ݐ�a�)?�H�B�?Ɩ��.
SF��#3ͤFRZ��\�������u�N۔����£���o��;<��a���>�5�\|�^<���T��1C�l���MP� )���������*��! A��z���ղ`@���
��r��j��Y����5�K��Pƨ���OG�8�h�wA��+��nF�R��Y�� ��$li�So���7�f䷘�ړ|S+�S���9;�pRU�o�LTV.28��]��0�)Q�߄�*R602FNYm�<<vI&b��P^�@�@ʬ���>h5U���4P�..�t��jn�$ﮰ�<_g������V�y�u�3�����U��o/(6�,H���op��8�4�%���9�ʥ*�	��<��:'p(x�F��!�.����O"�mv�sV����voT~͞|�a�H��i:dT%旕�����M�5\c����^T.��lm9��]�VN;�8��y Д��,�G�$6✺��	hSu/$�K��>~��_����߿��x)�/Tn�ޅ�~�
vs� \6$��R�����W����f��Q6Ix�w��!���C�J� :��c��#H)g>� �0�v��9��	'+q筡@
�ƈ��R�M���(��:���[-wt������B�L��C�n�U�'���A�������+7�U�`����i;	0��zC�@�Ř&�x�OE��oA��3����Y��~d�qn���`{���i�;��Τ�q,�v�핔��ga�N1~4�cK��[@�c���O޵���+�5Hf��\���"i��/�q;��6�K9l3ܠ���p�jt4k�-#�St�XFA�9U7e�c���M\��A���T��I9g����ο�4^w�M�	N��`�;��jR`��k�ߌ��|�P�~�*��g�Ax��l�;�bL0cx�ya�u�2��k��2/b�~!
`>����G�T]���������&�6�#���R��bur��U��i�y��������k&e��!�~�L���2L��pt�� lGrg��-�����fjי�ƒ� ��"^x�,7HA9%�ޗ��ddUWUdl�{��?}Z�c�'��v�±h�oo��"���A�
����<)
i;c�'j�pwV)�x~tkd�n~�V��k�f�i�9_e��>|!��U!�V|ᔾ8�/��6mO�G�y���"%��c
�Iΐ֟�M�B%/OتO��U�ŹlW�ʭ�9a�r��@v��w"�� ܵ�����8��� n�e��Fvur��⽡Q��e�*�9��v��1G1z%��?��H���.�g��D���3�����_W�3kE�b��W�q+��͍��;2�5y�4�J�O�:�U
j@��o�4�P��ٺ�{HaΈ �Q��dN��o�\*S|�I����x�	��9�%����:��L�W�Ӌ�Z�x���o�)���ujIjԨ�c-��@���>��0���K= ���� X������G�]t���6����o�K����S����Za�^Cs/�g�k�|�Д!	�P�H�N͠�H@sT�,���\`{E��y��)���e#�N}7O�Bwx���'%��C$��)�L�>�,C��z�+:5DB��e�Z~�9u��������ŷ^��,����I`	����y�Lc�q�Sz=��W��?a.����;�ǵm�q��h�)�Ik%G�����}��D��d�ӈ���o(���Hs�mZ7K���Fr�ق���`���Q���`��d�7����1Dq=�K#辘�">-���b.|.���&���`�ɱ�j���U������	���{dZ5A�Fs��N�������,1]��U���`)~����'�B��B��k�{8.�����/K���e�	�p��m���(��Os����I�^*�3�p2C��I���c����ub��ߟf/��C�q�N4��*�9"�qvp+1�7E��f�C�hVX���L�"��9\����R�����2N�P��((�y����&�nC����mr����%�Zۜ�}�8%0A�8���N��0��*��N0\uZWN��E'h�Z=��@�-$���|��Vj�p���-��*��j!��VS;��d��K�b�88�Ӕ�!*p����1U�g����!� ����ͬ�y+���S#�P!�yz�R��"ՙ˾V���B��Vb�x�b�$3�����3�Ke��Pb����&��I��J[ȼ}�J����*�7X?_����i�7�h����|�=[q4�M��I��\̗���|���^���dv3'
ef;�	꼨,��0�:\�k9C��b�� ��Cž!��A�J�X�Š.5���a_��y빓S�M ��� t���3�,OC;��SR���N��|'��a�3%�e�~��J��*�=4Խ���JeM���Kt/�"�� [d�n�B��2��ѻD��Z���*���<�N6���Ĵ��Ф�kW��.3>E��L�����sq ��'g>SԠ�r@�<�xn���KR�a*�{��ѴG�S">��� /�%�t5j�� ������@5���#}0�a�9h.�w�&�]��,�$���^�S��+�@&���j;��� �ǡ���pd���v ����45{}��z�7�
��x$�գ���nÕ��V��x�!��!� ����hr�[��a?%�sx���N
���՗=%~=>QA�Վ��`�9,�I�И�^�Ղ�afMF�W���Y$|�6.p�y��Q0K�٩�.IB�Y�/�����"�zL�sx�Z�)g�eڳa>���(�J[�� h�%s�	2���I����B��8C��DoH��e5/{)	�}����|�s��V�^ʰbv���S�aj"x$s��sɡ����f��PZ�D�Ay� C�x)q.!��Zݟ� p�;��t�ӸB�[�=�X�N+�*5����:\����6zi�~���,v�<��Wrخ��u���&���J-����?����M��O�w�Ȍf�5�BO���2��I�Fn��;�8,�)��GY�Ǌ���1j�f��YZ���9�zv�TS8��8���D6XK����o�FM�t؂*��:�������fo�]DZ8� ;��a-:��%�����=�bo���}�ZL^�4���,��D��PZؖ��3�־�l���?�5 ���2�P�j��q[�q�n�Y7	�,�3�|�{p���:ؓ腷���T��*,���L�R;�6ò�,+;�%�k}���Y���yrZ�NeA�!fWW����D�5�קT�j]-!"��M�mcEB~�`���G;��_������_�.6/p}AH>Bb��I6���-�?��<n�Ml)����[�H�ŬF%%��B��m1���H�:S|�3ރ��<N�Z�u�!�ßj9�L>��'lu���r�9'��撥�� �Ln�dJk�_����g��=˕'?~���/�X\������ Gfz��=W�	ß�k2�����(y��)���Bۍ*���J��� z�DPc^q��'OƤ��v��he�>�Ɗ��; 4��1ۡ������w�DS{C�o��/��E�ǘ���������F�L�҈	�$�-�������N��9��^�������;UwDqQV�kQ!��GUQg���K��S�n6M�s�	�bn(�%=�NLt�<��8���6����G{ZjP�R�@R����ڹ+hy�;���$G�x��:�z�	�hq��k��Se�����bGl7�g��Y`�U�`@w�
���Q�dw�4;Y�	��%���j���5N5��)�E�ns�_��m5���b|�l8��H:�xk�13ҧ�Y`6�X�\��NUX��dG�>&*1�i���^/M>g�V7��y����Θ:L��5(Mfn�G��u�W����WX��8~���;C����Ty��;j|�rUcZf������J��j��R�,���\'l&�0�=�u�?PS_hw�� ����R7�
�����P��������X�+����x�}c21Ő�7�&Ai�;��)�1o��kE'��t%�9~����n�I������5#d+!���<���F���4��_�c;~tC���)h����b'��{?x���0�l5��I���l��������k�n��Q����>�E\��)J��v�[F���u� <?ZD/�QTO�u�"`����?��x��]���pz���9o�QUa��N���tLߎ���<�b(� ����D�w��\s�w��d�/r1	K�V3��|~���&񇣖l6��@��y �$��ǽ�g*&aT����U��Ź-����|w���p�QJ�"Q�> i�z��C���ʃe��nxk�u0�B`=������h��{Nä&�	V��o9P��d��d/��E�4��y_�v�8?����w�U~m^�R��������W�D�$�P�_Ң􀋹�!�F�^�iWx)�տ7��g�x=��B�>Ʌ��T+o�������V�;���N�j�w�����E��z0jyd]�W'����;}ϩ�5I�I���,�Ѷ,�(w(��_���
WA�[M��'��T{����KǷ� LVaerDy�D�a3Am~]tn�`=�L��B���5�5Pos?��t��<���~��]6M�e��7�d�V�1����歉�ob�[�&��t���kOE���G2�����%4Ǯ-�b=����H���t4 �ߤ��D?C ��S��_��p����]��ݚ3M���s�ş��4&�a�����rB���?���9�U��%�_M~�&?��n�傰�T�B�e�'8����BN@�����<�g�i��Y����Oz���|�����?Ϧ�|ս~���aWg}c��wHn8�&��!� �\	�[ߎg�&�uR�	�azx<bLD�u!x�|ڴAz�hhQK�=���&p��)���3��x�"\�
�~Tӟ��7#m𠚔v�=�x"/�џ��|�8�2�-o��:]f_�3�l���k�����=��MF�Jq���F�L$�jG���ݰ���ȳ�A�n�>y�@{���|TJ0KDr�VN�6[��;�u�7�ҴWOv%LL��+y�t�^X[J7��֤�|�۞�*�ژ��2M�<7���k}s�!,��a@M^��O̐�BH9����NÁK���f�qq�-���T.��C�Q��Z{`���^�,�Az���K�i}�7��L�L��#;�Di����w��U��I1L��j��{�����v�����߃�or�y�K����;�7�ŋ�%nDCHض�����W�5[k`��YH��s���)�"u�ڃ������ݘ>8�r���5�_��Bꭍ��*zb��(~;�ZǱ����`XB��3:tM] �����Y���^s�F�x� 'Hץ��ޜ��i����Tf��>g ���h��c�[K�9e��L�ҍ����j�e�v!CԮ�ǔ�:�;~�S���-8,���1�ԙ��'ϝSՠ堛7�:�~�h�5�gь@T$����H��Y9t��?�.l"F��{ޏA�:8n�����]�z�Z��@쥁K���u�����߃�5b(K�2�<�*�>4���龖�|�t9=�J�U��SV?7:m���J2�m��z-�M#�3���I�	 ��Jm� ��B��i��n&�M�DE��7Ǣw/eB'~_u��\�i]�6�t��w�>̞}� ��!ۀ��|t�G��
�n$���J��7(s��I�<��>I�r$��:��':�>�A�qX��'p���	u31ww�V��i�JD�/�m'8�K_
"���ZW��~@S�`/�]{6x;���0�Ox �
&I���?"�ۓ9 ؀F7냔�^s]t��`nh�Z�W��zg�ߜ��I5�/ ��$I��O�.���Wy8Ik,���A��;���Z�z#<x)(��6(�w�#����,�VݏY�Z�p#��������/�61��=�O�T:�6�Oɂ�ןd�ϕx�R1�k�4O�$��	]ĭ�Y���GR��s"�_��JV�pi�{�X��2[��8����4>$.0)� v��%	o��g4���zS=U�����`�4VĀ*z.	]=��˧�o�ibbwyp�q�X]&>���Xת˶�֎�;�ehV��%!�.�P�LN�T����JY����.��勤�X_}�ҧ�	&h�e��u�_q���t�£�y�}�[R+�!��u:T�i�Ft�5v���acO
J���r~���9�����z3Hn|n:�Ϛ�Y���Y5&��	�Q��3�d�$�[�j���wg��]��%#��k�O��&ɞ`��ؕ���,-�;}���90�W���&%L�-̞����J�Y�\a��:��&ݣB3�)��}����@a��p�I�%e�;Ί�����I�S$_ձ��+�g��y���q�w�!�����A~��S ,�:

+**0�"�?P �d{ԯٙQ�G�2�����0�납YnR���%��c�SsHi�	f�lZc��ެ���7�J���`
�G�c�SY9��r��������S���
}�p�M�tHkC�m��Y�%>���,ȉ�sy'Z{5Z��&NT��$�v�g�˄�&<��FD����Ī��[�QC���X�9�1Q�:�1Q�۱���IϢ&����.�K�]Q�l���������VJ�t�f���s>����D:�T�p3,�C+7��!���Dv��=4�����]/��p���\*���R�ˤ��C�߿�r3�ԙ��>N͍B��\_ulɩ	z�Κo�P�@S�CKr�^�6�o�U�r��20��x�'ȸ�H������*k5�x�S�b��X����Yl���<)�5Z��3�/: 3��#����-b M��
��a���@�:&��f
��Q���/�ò�W�AT�<�n�7JV��[�v����BMf_���u���O�|�Kn�j�"��t�,�v�t`j��y2� B$=2�Δ 뗵p�@��� �)E �w���ܲ���G�%�LO ����8>�G6?ɱ堎U{d!Cn�����������{|���#&���|� ��[��&��&Y�GΟϼ���\T`�v˖��(���sw֧�p�i[�ܣ�J��b��ʝ�Ae�|Dsy͠n8N��j��^���R��l�:�@l+�jAŸ��YY�H���'`��pZ���+8üڌZ�Jh���������t	���g����"{�l^?_������ �O̳����ԮKCg����*�0�]/WmL<��*����K2��Ct�'%i1�/B��ϖp�B$��j�4��g���D\\�<�q��<;{���T�������I����:=�<A�)�忢^0���s��(́�R�����S6P�����9���Qr�2��R<��I�>:q,���xyc/?r|�C��*��`.$��W��NN��.&g��K��I�	6B�Wu��V��a�TD�^GE��<�:�'����mg�)!4�p�J�sM��+�~!�<�:d�&��/��ӂY����wV�@�F�G@Bb=m %[P8�PO+t��kK��Z Q�	|�/��?���^�c�� ��,S��l��^!R�9���R1��D@�ݨ ���!4�غ��N�I����#ш���H���L�_��4;\u����؞�]M-lG�⩬y�~yM~a��HAE���M �����5���Y)�u�'s�c�?D�t��̢<�����y��L��%�3�'�c�=�%	8��߷�:�����C����� �Sis1Z��8�ʡB�w� ���'`˞���W*i��kV#��6��>�5]�d�zL�� v�/����On_���0�>�S�&1q��8�^k�q,�XC؇,�l�"�+�n��ڸ����1�G���F���b�~��e�I�!�X��(���[p"rݦSO���y��I��A�% ��z-�@�{Pm��������o2Qh�s�~���2�r1�^x����))h�H伱��o�O�#p�U��ꬠtoc�����/�$3>����Ba��ov
*\f��x�=����5et)��w��1�I��̽�c<L�C�љ�o2���`缘��fď��V�場2:r���r��]?�^4�H|j~���J�2��HF�:�D��ׇ{�h^Ȟl����qkd�H�p��f��/=7z�К��/�����]��+H���S$����P��y5>�H� ����aQ+g啼��	��9b�R ��@�U����r@�wLY�e8�!��ح�S/7�� d��gg!�w$Z����H����%�A���yR�QJ@�Ԉ�_�W���U��|�%���!��!M��(ڹ���R�"�a�*��r�|����HryHg�l���fapT��|��<���:�����I�|�StHy�?�ҙ	�M&�M���Omd.�nm��&�Xf}&��M ���e|�m�L��*��^B�V'4?�3�i��[�?�S����t��)��Wq�?�,��/o�u�^�/�Lͭ$�Z��\��t�=$/-��)P̹��H=-�S�%Ȓ� R���*�Ef�җ�3>�����XnI[p3� s?�l$��˳Wca��F�!/^닏��_��X����]�����+�����[�$��v�m(�/ڶ2
v����0�0���'>G�F��=���.\�P�ɦ�P��l�*R�5�[A-��;����؃2U�y蕖��n�'�D��9��K�hnr�����◆�/��~�0AN�3��%���[����yR�خ֊�D�f���?*�	*��Hӏ_��MU� tA�Rv1� ��h��ׯ�s��~|��!��4�؋,��%:	��,��!5��g��_t�_>1&~�,.�;�Pv��j�5Ո'�Zk��6������6�줞\ɫ��=��'��?��9�+3KNصC|~n��Ժt���H1�{"����~�9؈�l0	@�9��^��a�Tx��$� ���O7����,����V`0~���c�|��,��%���CP�֬��:C��Y�a����Lv٦"#7�v����_��f�*�q��hZ����V�CZ*�6ry��p���;?�/�pJ�嬨VZ�|��Ǻ]�������䦹�`КW�k(�z�<�pcR�O)dCOh�p�X4��e�B�	$�ۄ��	wtL�6龍�{�v�)_83���2ߊ���99�Z7!�ʄEIF�u�rb%���m(V�]�zvZy��/�;�"%�%j�Q�<�ھ?��DL�����Ԍ�ؙ������J�<����]M!e�V���7���LL��3�ɉ�+	�����@���'�Z]�-D.���Yۂ-����e�G�n������^v+w��^��U��^jb���a�z���2�?�f��L�xگ�i5�a�no�!�SU�[3O�į���A��f�]��2��GJ6���|�x���s,�oT���׎/|#�x�;��R�Y�#��!�ߣkzQ��16��!�������'���p ��yc#�PJ��}I��v�GJ2�A�a�0�����՘�-
��~{�+J����.��ŨB#����c���֘[FR���m��9өM���TG���{A�º���`�?�`��1S&>����t���l�F�X�j��'Z���R�P>��w?�қj?;ɵ	�Pv������4A���ʞ~��쒕�`~�2`��r*{�1Ue�\��T�����d�H�����i[���RDTH���n��}�(F�V�фMU��>(�]`j�2���b�"�Tv��>���Czoq���z?�o̦ݟ������^�"nh�<�J�i���l�&Û�D%~�@EO)�c@
}F�_7گ��᫨�bY�N�Ń�ƕ	���Cl��'���L欮�B+b�F:��7U��z�x���G���e!B�m8H�oͬ���-�B�¢���aV_����'�Է�a��P�Ɏ��sԌ��O����� ģ&V��bJIkU�����
�r����){�8JuM�<i�kN.����h���ۮ����Ng~���iY5��G�U�Җ��_#�bX�WR4$v���M��Q����;E�x-���K�+���i�ǒ��LZ�[`��֬'�8��<���es1?�Ÿ��Z@�h�=b�g��w�����l�ʐ���I/Q�1���T�2�p�Pˇ?�9!��B�Iԗ�S�&/�ǂ��K;3����ln���g\���i�0eG��ڹ��323�[?Z3x8Z�\�|�g��[�3�{�TUbZ�T�{G 8�د�S�6�}z1�7ڗ�9����qA<D4�KNH����<)yic Eݗ*��^G�tI�0�@���z�m��/#�~k�6��F�G�V13�|���Z���~�6v7�h��%zGD�v^�k9��i�ޜr���5I�<_�/�*U2Aյ]J.oS���<>����bI$��@�I	=����S)�2���+�@���:ݭ�����+����v 
��M�meF��;.��ܦ(F!N�"���2^�ZU%I:DBd�]�(�i�K�����՚J�m6����,"�\����MQ�ԋS_�t�#�RSFY�C��u��y�Z��n�(����
��^Ƿv��=�k��|����c�T����f���}{{��q��o5��h.��t4�eVڀ��ж ��u0D�ϣg�R�yi�5�%����Ȼ=���jy��3A3x�VhXA1���|��U�gJ����'�}�J�H��ҟF��H3o�Nݛ56���>I!��'��$Nv����j��k+u��S=�M�=�V{�Z_��Q-��LV�rF�K�q��ȾD�2\=M\&��b8��=��*eʠ�b��I��P�ڝ]�â���p��Ep��œ-�[��`��B��}�_�&v5N��N�3�֑Xl�M�i֪�r@��s�V��p-�5nɱ�t�=S��>�������1Tt/ٯ<�d�ݑ�&}��������T�}�/���\S�>
G@Xn�Ǡ����i���g��){ٛ�qej�#���}mTOl=���~b_"�n�/��>�X/Z+�w�2�x�3z�y	�(�@^���H«5lϟ����f;�؂?d.*��=�Z`�Ht�����:F C�a��V�єZs;(���a���Uo2�-�4�MQ��n�s�A��
)�AlW�d��@��#W!�
�<D�`{<�3��T����o�E|���՗��Ҁ�� 9=��W��=��Vg�����C��qT�%�����t���1kG7��R;'h-?��8��8fuqI ������=!��.8����0��W��̗�8�b|%���tcv�v�hl�_Q#C�~1�C����5�%@��mf�X��B$�G�_yR�+F@H��|�I� se���p�`D�'
��[��Xlf�:�BbbNc�4�A����5�M	�ZQ��"����3vt���"+�YN��GW�g����.����YNǢ9Yz0X/�\ӵ�z�R��;ܻ��2&`�����.��<��(��Y�rhv��G���Ho��7�Y�=e�F�q���*����ҪR2��2q�e�zAm���s)�-p�w]�E�Lb��p�
�;���	���\Z��+�.���i�{��,'��y͓:Aŷi�(��s��Ab�kv�'>�����&S8��2"��Zc��^��
B0��A�S�\I���2����z=��J2)�f�uG��)v��XkP,��FrO +������?�qZM�eQV�(k�J@a�S��J��3xCJ�Y���"0��F��ҁ���a�Rkmx�>��n�_�M&��z�k��P�����D�E�����Y7�u����.��W�v�y'�#��ic�:cݝ�bR�n���W�+�M���P~����2M(�w�]~�sF��M��1���);���M�����W04�Z��q��i�E"C!�:�Y�(�