��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQ�k��s�#��ݎ�4Jh�}������!2����s���kW�YCu��ߥ� q��j3��:��ʥ�C0�S�m�lf@q����.{�.��Wgۋ���ʓ2v��K�U�@����vF63q�^�6��\��-l��P|<��K��S���]VL������h7����_���Z-�:K�ó/�-M�fX���I�S@�F�R��b��F�\��Ǜ��`��dS�L½Wǳ�/y�nV��A�Z>y��k(�<�W��^8���W��;�u)u]'��̱&�6��*XV�����2VB�98%'|��(H�%�	��9N�T�1Z��QHJ�T�a/���,,IǼw��l����=��B�&S����I�<4�@#U	8n�j�n}l��޼��櫐h�G��R?�x��i�ҕ�$Gc* F��%<	#c�b��M������_��{nГ۲�� �C�۠~��$���Tp'2�՝��Z�Ō��9������U�_����H�
�ȂQ����}���A��~%�*r�/T�"����4��}N(�t	���r�X��y�#�<�`�I�k��Y@�
rA����Z`s_� lc�O7��WcY��ö`ă���|�1�b؎�Z�	����km����3×Wh{��l��o���C(hEII ��-:�2v1�}�$�4��VY=*8����G3�&���������K|��ngG�S�)�|�t�zn�ɓ?n�L���99��w��?���䇏~��=�r�&'s����}<}k�	�e��*��<s�l,�J��3�8��0�o�v�m���:w��Wt�~�	]�*16���V�0!�<�=@v�����s�3yx��T�X�a�S�{��Z�HL)�JeT�D�sr��n��k��@�Ꞗ�I��]�IpC}[df����������OkY�O{ɛ���H���4���%�:0�c��^9�}���^)��&�qo��D
�hVlkl�X+Q���� �T�>�q΁�Z%%�&�a9;"�V�0�����c	60 ��Iɯ���-[��7С6�Q�R��j�r� ���'�)3T�y�̘���5`���x(f l�P	"S�Z %�`� ��z�>�:d��~�����*��c��y�u!U����!���0�HC{�ķԬ�`Fڲ�(F%mh�>�(�o9�8�tì���U�����ql?��gXP���� 1�[ګO����i���c��Z����تIU��e��Vo��"a�%F۰9ȗK�a1�*t�p���{㚫@)�Կ�Cx�mY5Ts�̻��P�����oQ��C���)���S��PBC� O(�R�T�di�B{��9�Q� ��G��7���cw����yɧ+�8A��lc(B�Y?5[6�l`�ÿ�V�WW;�84�k��#X�Fؒ��7�u�.A9R��{��6�S�K)��cU
#b�āL�aOt��.eL�b�PBA�]L���I�.��Y�|m-~AњSmdĕ[���=|���dYM����������n��o8o�Oڡ������k���'$i ���\��>9�+7D0�7�W�%;�~��d=�ߙ���=��������b�k�G~r"���f{���/����V����ez���i\ߝZ�C�$��VLg�?��e�����9�P�P�@u;�d�aU� �s8�l&=�����==ա��6���覽�־y'j�e��^qe��,��O�Rdd�j�� q��-(G�Y���P#-�_���X�T��d��:X\;�D��6w���	4N�#��q���L���}��]� �P�T�9L�ʿG=Y�v�r�:���p�#$���%�� 
�|���7��C����DV:�|-�z�߆2'*>��:l&J��(�&-���s���$G/_�� �ڸ%�C!����ޛm������2����(���ĨXiҡ�}��Ǆ�Ӈ3���#gTN���`AU�ɗ��%
�����b8ϯ�'2J~nxc��FܮAֹ@�0�<���$�P��e�=���*�I]�RL�BWT�?���jMt3YH���7\W�5ep��$���A�W�؁]F]���"p����1���Uzl�u����#�X��l��,��M��痽�9����,7�,�WQ%��� �j~��`���j���N�K���H�n�i�\��s,q;�-�W��o�	I���銕K�I��/'c��܌�y~}>��!��I��X=�����!�eQ?�0�Qu�Mm.������m��tF?*�&i�}/�(�-dr0=�e�_�ٸ����'�����$p��ʟ̺�-%���()d�rR�FE8��lr��͠��[���S�M�iˬ}�J��J[��e��:r��O:h�ǌ4o��M�bM�i��T�biq�a�O�3�
H���!��Ѧ�m�55�0�Q�0���~;&mV[(M5���k���0���Fɳ=%<�@dh[݅+�dp|'����U��}��J��z.b�ѳ�40"�r_;�e�Y����×�n%�-�q*a��� �M�n�/��6���㭬�۞I�
�l�]ҫ����-��|V�HCF�.�d�'Q'�d���i�h�ڕKB�q=2��Âr��*g�=9�*���r,�u�5uAB��{o��y������B��`һi�1 ������O	.\����Ds�j�\�98�<�����_�#��x����@zU�꧁IL��xL�E�?A��Ff�k�8t!�Wj����1(�.�:�p?h��9_ܓv��Q,
m������<�x�,;Б=0��
Vy��.ʝ����s��D�U>�XVu�0���n=�&&,�\��o��r�e=����H���UE౞IKƭ'JwO���N�G[���w+s�=���_��P�8�V���F���
g�ym{���;6�US������eV��d��ҢfL]�#u"!̶"ԗB�Ẍ��PAW�<ߓԩ���L��e�:��ʯF�Z%��5�0M�3?QRν:?q0��������MkBٸ:e6Ր-��f"I�mB����J��6zx`���r�(A3f,-m� હ���O����q���!n,�}+GQ�m^�)I>��_�ۊ�io���"ri��N�R���)�w�x��c��d��J{�B���B?��B�j��ǁH=�a�v�bi��bX_Amu��؀>���5�O���v.���^'���]Գen�A����Qֈ���t��3P�M�ݰ)�-�>�j�s�m���i������[���0��~��"�!��h�4��d'������U���~������$:&�vC�X?&4c�sj���FF� B�C��:N[�����mˬ=�i>�எ2W�d<����x��ߓAvV��q#����5e��C�ʎ{RY�z�m�~�?2�j%ʕ�/�?�o:zU�$0��%c �$�Gز�tK�4�|���f��Ge�ݪ�x�1�(D_�ߔ��yHX�خ/A=�z�6����y�I_��ǣb{}
n�6��ȳ�r�>-�D�%&Y���+O8���b��}�(e^y>%M��ۤ���B�G�}�+��!-�?s���)��K�Wo?�Ve�H�:��Ca�aEצ�����ES ��u���v��u� �#��T�E�!�^�Xi��5)�3��ϛ�0\M������n����tIO�0;\{������|��j]P�s�rm,�(2��y0��h�j�"�v��}�+&,�ʨ�kԎ^]����q���\��Z�e��ut���7?��&1������u7�	�wB���RJf�r����e��;�I� fN��Cv����Jo>J��w����@g��`�E;��rWh�;:����bEiGW�\*+��*����;R�S}��Ó��Ϗ��l�w|��d���R�)_�0HeM2d��uӏ�X�A�G����y}Ù��hh�ҙ�����*�,/.XN����T��-2�0B:0�v�y��Y���j�a��!�����M�Z�;�O,c���h|n*,��	];ԏ�buV�5���e ֒*�L�KK��_s
��y��e�|� ʷ�~�sUc��8Ix�\s'G�nQ�S�QA���0{W�s��nQۤa��\�Zm�n |_cMđ�a�M�m�jҝ1~�3��]Ph�[O8�p��%�g��-�(!{N�����?�ƻ`!V)K��>�_��Pw�9��E�c6k{��6�`ja���[�l�e��8�f	��coS
ӌ@��uQKR�3w�
r�]I[i O����0Z�b!�.��3�p���>X]���
y�y����az�U8�M7�A9/�B
E��1�Z� ڕy0��?��ݍ�����Nc�������g��˃~�=+��y�u����T�
о��G��@;���3����l\�O�XβT���i�՚�𹮴��.��	�"O��mV.W����c0h� ��!SxD�
!"�7���݊��;j-����Ϲ�2:Zx,(%����%�6�!�>nf���+���w �|�D�������*r� {B�����&+��3x�j�Q����k��PI��
 �������,h���UK?E�96X�kϋ�6� d��V���7݅��:?�3�̇�X���(&vO;�������m.r�c���@���Y�@W���T�L����~����,�zo���� j&���1c5+���w����E�z��������9.���.�T;?ÿo�I�ˈ������
 p(�,�gѪ)�^����!n}���37�T2������YܖQ�(VG��.��P`d�TL�:�^t�����x:���b6�"�Lk���|x�(�Aq��yÖ[�=���%����� LΖPh��T;:Û6<�qů�t�UO 
� �C���"p-����.s~�od�ʯn:�ad)7��+�ݕ	��J�@FP�q�˩4����;N��5w�x��i�.N?�l0t?�U5R'��G��4���$AS�	����ۦ��t�����tնڳ4B8���V�naI�[z �����ƏJ�3M�.���^s��YE���~���W���k+j��� ��i�1�bL���]|8��F(Y�o�@��8�����[�)6��<��b<^S Vϻ U��+��7i\��r^��گP���W��l`$�����z���Ҹ�Y�*Q�i4��5����;A�Wp܇h��ہ��R��I���`��sR���m�aD�$5�q�{ �g(<��9����{�����no�'���1'śyb=	ڱ��������������R�R�ݢ@��Z��X6�H)���0��_�� *=���N��6T�n�Qm#<o�� �+zl�/���Je-7ai��G�5[0ۑF	<^ZT9�ch�����&���>�1�Ӷ�bǛ�VDc�fw	�ݶ	H��X9G���ʔ۔�+�{A'cNp�gf"�'%�(������2Ʉ�	��~��]F�d��2�x7[Γ ������(tWfBV���A��'$-��'���ѱ�|Ɂ6-ȃ���o�n�N�&Ϝ����ȿ�*��P3-�X�<� �
dE'�z��q���DSwJ�tu)l�A��7EٿN�|�'�
I�.xPA�rZ�e�D��W_����LLUp���/\f���zѿ&��֪>�[e.CkmYq�
���4��#����@gb�D��9>�%�K�M?�SUZ�{ OS����,e�R��r�2l]J�!�l���.N��{y�3l����aY*�����U��#sd��s!?�7��:�vķ�2S�G�u�52����:C4����ЧX�R�ކ逻�p*Q;�ŚQ�G��P}�m{ir~n�#�BI�U2�ס}��f9�~��̇g`h�vɑ U��p����9tJI��U�\�ߧ����)b���MT�<;��yu�Y�@�ز8�ȿ��PLؿ���>z:|R���sRC����}��m�}��3���޻�{%������2,�-���G��6უ�Q�eH�5��?�AV�������%�d��-��kϞWJ����7\i�׭���/����:�>���ӿM��&�s���L�ruԺT:�Li�<.<t�
�לv5tD�X��OxK5�E��Btc1��s[�������R,7r3�|�,�-��wS���0���y����~�1���~�=%�_׵8uA�]M8��-�d��FU���%�Dw14-~i�3�H��]�cnL|$r�D��OKP���V��`���Y���lZtDd��kК>9A��W\�`��)9��5���\o�`��-�{3�ֳ,i8\�haJۜ�cqJ{Z��{��i%�i�\�4�����V�ep��G@]=�&[E�#6j�+�S?Y�~ח�����%$�d��a%V�W��_�|�-�I'�����Dn��AE���ъ���*��u8�gW�$?�̦L�*�ς�|�1���gA񚋢�j(�mc�!Îh�,�P!S�&g�^�M����(zD�PY�#�������ߔԏ�9�t��d'��ӿ�W�Z������v�8�h��nٚ�n|��$Q�G2�оz�����-��ō�f9Wi�-.W�v�Ę��	��J� K��덓���'�$�F��u��s�d*�pW�r�ܝ��#'7;��K��D�`;S;��H)���5;�g&�,E�f��46p�����ƭ�P5�K�C�a�c�f�5�$HW�Gy�>�V��dz'o7c�C���5�"�<���el���7�|�~���-(���$@}̔G�)��^��(-��uT0��9��uz̿���s����5��8ж=X�Yj�*]�����yh��#����W��q��5����X��t���?k#sT��������_M��$ȁנ�t���.*-�����U�Og^��~d�$;���ں�o��8�0��%�>���B����Ú�l�G��6��"��&����������ѲoB	�QG	�1@(}�w �$/�e߆+�u�4���k�?���V�e����0���f�ti��,�Ȥ�c�x~�U�q������*Z��?�P%�OT���E�9���9뿽���y�s ��h��0�祿�u��c/�vdY@�'�:5x�G�o�Rx�X��1v����w��:�{�l|��sK�DC��!��#�uK�f����p�!�y�/K݉�	��y:�c���D-��} /'+�M�"�`9�N���M�ue^lvu!Y4¿�L�6�}��PT�W;׸U|8�� ��	b��/Ll�
�2���K���@э�vB]0\�M7.|تP9:����0�R�%-����Wȋ_^�MV
�f��5�Vկn�.���:<�ڑƠ�#�|��L��"�r��M����ۣ"���KN�MIt]��[���?ߙ��Z���gg/�ǚ@���k�	�v���3 -����D���G�"�Gܤ�-�َ�E��Z�!��|�V�9C�+��g����jMAK�0?�ϣ�8L)��`u� �~��Ψ��Lq��tB�A�PS�X��-Q87�ԝ~))�O=EMN�� ��o�\償�{6a�W)�W~Q��Ѿ8b���O����~�fts��vi���a�Pb�XO��4��'�762qAϫ��.=n}���|�wqXu^�V�J���2��1Ǆ&8v{�<��.�mC�0���� �3;��c�B�,=��o�	�/�����&p\T~�e���p��s��n�|�fKT��Mgmq����ⅳx��E�/0�a�o�d�x�)�����ژ�
�V�:�����Z�~���69̂����=A��-S���r���>nrm��f�����c��<�j.lc�(R��~��+�����fе�6
��53V���T2���9X̝-���~�o��F��!A���:ԕ���o���<fs�g��4��Md����_e�hs\�nN�-�L2X��B�*�RR��Lު���3�A>{�9H�S[���50����p+Ǳ���.��)���|j&�7A����ہ?���J!Y�lk�;�D&���=[�RHz��Q�:�5V��}܅Ҿ��I�,�k|������!TO�o������6_jv���g�"�)���j��o�"���{t"��@��� ,}�*ְ��ʉJ�F�S1���n�yH��vH.]4j�P�������y�X�q��˰�YV�v�u����|��'%�>D�k����yk-�d*)$���.4�N����E!;�%f\�₈���!�zl #��}��̄�y�j�)س��/�^mHwR�?$e�H��)	)��L�׋7D�j*k�k@�*F�6{��y(
��p\m�s�0͔.m/� n��"�����FKH$��ۆ���������ߗp��
�U����Hg�ãK� Ys���ڇ*������������"�A���a���e���ɘ6
<���\藺rRH�n�L�j��-�!�c���G��q� �nw�Q��b��#	>ʕ�V���Rݱi��}Р�E��2̕J	����(��hdq����LH#%����p�5���R���M�+s۶�g�r[�>ܗ�]B�J �6�}��dn�r~������/3�_�T�G]��r���3��*Ζ���x�Rc�%<Y&� �Q��W�h1E��_����]�\�_M}F.fMn�8 �>�׫�G1R�w��̪a������g$�pa���h�/��~v/����	{_�-�]�3�bZ�ڵ�n%� �0�Yh5��7��9ms<$9��K����#vR}Hr�7"�<c�{�ē�Dd���߽ �U �bP�|��������hs�"Ƹt?;��R_&�����ÿ('�Ε��P�W* �J5��Ytc{��X�I�f�t��ROv��������K58�>��D�^(0�q �O�L�{�?�>�r%aX���]֠���w�m��h�f�����e�a(��� Qj�
)kmW; a9��o��/�g�8�t�
���(�};���I@���p��w�'��������r�����fޚ7+5��T������<FE�	�_jf���$�W���-1��G�Ѫ�N��8�H��+�u�u�K�K�6!2�� A(CYG�� �=�k$�+a���_����e�>��v�)��6���i�X�(���7a������6̽�H9�ƚ��|&�rA��;[���o�)M:�!ܪ��]�҄Y���3�$j��q��%�<r�jvց�W�3�2��i��C�P2b��)q|�oG��͛��/��C;�-��	��)� �8�J~%�V+-��Pq�������ʲ5�[DFD�!�SFA��G���� �<�����7	a���t_���(j�g�nR����9%�[��&g�z��@�&T��d��l�T�dj3Jqpp��*��
��?�{RV���C2��R V��f��j~�L1d�rVϮ-9�P�ϫ[P��'��0��%,`�?�7K����b^��f"(�9w,�٩����~-�y���B$�̘���<&¦�<iw�^xߟF���= ���[EF�Hzh)����Q�͆��x�����'����A����~ܨ�%��~� �k~����>�z�4�iZ`T2|�x؅q�b���6�3������A&	z�9��p�.��c0����+b�����s���<�	D���e8�ýD��;���\���]� ��a�.l.�M�$K����ۧp4ŔNx�|�}*Z��N2L�����_h07n���d�)�@�f~����BU�e�3��(� ���븽|�Ž�PTއ]��>܊%;�^F�	rM3�47M�ƶP�?�D��c��l������)航�]�1��rVhz��;n�|�S��U8��TH�%lw"�3��xn`�:�@7v�ɰ����jt��Ơ`��Ֆ͉�Q/�FR��#�8��9Uۙ[���M�}�_W�`,�FȂ�~7ߴq�%�ȁ
�[G�zg	Yu���'o�����n	L��6(�ԃfQ���K�:����}�xmNq�e:}1�v�n���)"�����%[�!�O��SD��j��0Pm+��8�18&UX]��q
�e$$���u��.G�m��8UR/�XK}�	J��LEA��U��&��_,��X�������g��o�*{sT�xAA˕�����Y�O��oTp�&���u��\��pף�v����-�̪W�,�? [�u��
��%��Zm<�o�r���W���EY�EH� @�+�q<rـ�����mC;��$�2>�@���Y�gr1$��)#��׹a�=��X�W��E�ҞY��Vͬ������S���s=��:T��x�<r�Z��L|��\'v�6�Wz�X4�v�_\����&�p��o��A��c����k}����+�>Ĳ{������<+���7T��*��Lb��%�!��=I�h����K2cj��1H���~�OT��>�ˏ�L���%���U�Y3P�2��W��Ҩ�+��"l���a2����]0�0��Uz$Ō���A�(MY�����T�+��U���6s._T�Z����O�m�rT{uq��Jb����0tX�1�s�{X M�?2������B��W�LO��Fhr��o&tBn�\�=_rԊ>��5�G����_1�P����o-�\;RQQ�c�� 1�9n8�4]��L��-��RHX�I��g}�D�)5bPY�!:'���B�3��,z@M�W(��7��4]��3��lE�����o�n}=�$��3ѵ,����B�0#2�3��K���2��&<�.��|���V���Z�[e��~�r�>AR�%e�W�y؁��#Q�?�U�n��u�v�8�Ƅ���ȍw�/��e��HI�d�o15Ms�!�S9���<bиM��Ġ��:��)����ӫ<��������\TPX�#��͝9Z��׋��A�xO2e��M��x�m�r�I>J�&�-����Ƚ�B�ԋ�o��"3H��!��ϰ�w0��n��ɽ�����S�S�?Ȝ��V���j���[��kdz�-���WG޲��B�&LU��"�RT�ЛɎ�o>����2�zɎx/�~n?�^����Y~����@g^�N0Y$�t%��O�E�`p��<��(Q��hs��[qw\����J4o&~\V�o�̂�|9�G	�"�/n$q��u��D�7<}lEĴ!��W��ڗ��RF��^[�Ds�n[ׯ�5Q-�.b�e��;���(�O�a�d4܊��j�j�<�#�e	!3���ņ%+Yb��v|>cYF�䔫�@�	WZY'B�D_ⲷ�$�����d��F��r�����l���-M�����~\�ag� ؇I���#�*���wl �X���H�J��^�3+�0D���̞u�s������yfFcp�Tf
����ϡA�V�$��6;�g$������޵e��R~�����HI(>ڜ��t���8-�l�	Z�R�p�hϹ]bX��w6�?�?i�h\Vq�7�f*�B�+1u^������ė�XG�> Wg�]��>���}s��r7�7zdѰ����|�݉mc��CW�}����o�~6��%dzC���UgT���l�r���h,O������ӧ�:.@�n��u:�6V��e��.��$���F�£�JX>�'7p�*�|�\�T���$�Nt����������^W��8E������%�u%�a��F(����$� BM��?�� ��M�Q��P���׍WN�<3�~���kṠi��#�:�=���	.��١�� ��6��#�3�u�+��v��\UJf�kW�_�cBl�1R�K1�PA4p��H�����@�V��c��[���� T�U�>�mm-�4�����fa���~U����V�1q�onc�8������#�[c:�?�0L kn�3ҸY�#�o��W��Nqq\�鯎����[�F�sŎ�j#d`/������E�W*� c2��/�-K�UG(d!��9�-K�_��l!���(꜄�|��b{�� ������瘩%y۷�wª�>/f%K�[�8�K�!�7�4��"�p�Qָ7��].�#H�8��^??�,���G�����m�_���q������Ԥ�k� ���ܱ�L�}m��L*�{X�[�ʨg*}��!и;��6x]y�B�}�{�fx�f�~9�Q^�O�A�<8s�2��Y���p����N_Z��+o���`agOP27C �6�ý	og�S-ul�^�wr����ÏJ���;
E�i����t���0=U�D�̔x@��R��S65ź�%l�i�b�)U	ƹ\tj������!�~�ʤS�	]��/���% D�X����¤5R裌'��`���$� +:q����?O���)���!�҂�ƃ������.,�M(a�ib��4���8q�o���k�c��b����bb��/t�.C\l%�.GIL�6������&��W/���-�А��Mm�_��hݽ�


,W�¥BdS��	Ŀ�LǬu9[��u^%��"4o����`����YE��r������������B� ���VRU�L���0���+�{b�0��0����G��|:¬#��O���W���>,��"���˳#M���(��-��:�v�4C��$L�=�+S}�M�xŔ�ٮ�ߍ
�5���H����-��\)N�e�{�����&Z{�>v����~Z��5Z��+��C��DZMV��Qh����2�	�|&���������\2o/�,q��9`�i�­feb�"{W||�p�ʡ�~�m�h�Z����]#B��)%3���	wt8ĺ�K��i��oCC�dPz|h��/=>3�A@��%3���]୶h�J��9ۿB5S���!ϛ���Pt~�2��)����0�S pb�d�-�RSґ���#����?�Dr�Aڑ[
�c��^�_,K����/W�>t�"u�M����æ��{��Gp/~��t�Q�^�� 2�#mB���"����L�G��8؟d��������.�;�u��1�қ����y����x���=��8V�M�'>Y�L�d'QK��bG�ۧ���O4h��� ��0��"(��w{Yp}��4Ċ�q�Q�*����!�л�`���z�B���SLBnZ�Zˎ�^d3�};:8�0��[M�P�H�4�b������Y!r�1����NE����&[x�ߞ"�+�����-��i	3P;a��k�c��^��Qq���)[:Kg�n��[>[��X���?&�u�g.}��Bc��

 X'��ah�E=:�qe>Mt����ZؔF+!������l�wfC�Wg�U�M�Z���zM���+�z����g��G,��pp�*;v
ܕB4U�)��,HC;���
�¤�=�٠�	�Q��_&�y��ҹ;v� �.�+���!�5]�*ϗ�������[K�ӏpC\�%����>C]�Q�� ��i _���{8/@�Ԏ���T�>��&�b>������-M�N���<ll��|~�0>s����?���$O0��YQ�0y��������	�8�\�d���씜����z�C}X��9,�\ak��7u;ׄ8��Q��k��	rR��d�RěWa�����8zfߤG?��5�zq�P�t,G��x[� �N+���3U��0U٤�RD�yG����6�?9��f �1T�?i�ߧ�ǜbў�u�A�<	�q�7�8�Sٰ_�e�dBK.-.�enIU��9���%�0��s��x���%"����,�����s�{��>�{,i3�c"fd	_�x��������p� �ҏ��
�$�%ް��D�D}��?��%�yLt;��$����0�c腹���+$�i��h���Ϩ���g9\���l�ҷ�o����{#��h;H�S�0K���\ >��Wѭ8L�x�U_ݚD���D�,ci�x+�|.�Vz�?���C����Q7
wR9������x�Nt�b�	^Lh�fHl� �݇�`A����=�N3���ֈ�!�ǥ9��6����6�Ƞ�7�_ڭ���'_�]��+�7���x�}`�48ҷ7d�.�c'X7�sˁ�f��`����k{��B�,,dF�Qy!�Ch������xZ��BI���\��f���u"݁�����n!�ꑒ
Iq�<4��c�������8�è������4��q�|�]I���8&��%s���^a=�8���m!X־� &�u��1���lN\t���o'-����>S.�.�o�e�J4�_5�x���C��Sf��#�hY��[m���;�����ІLŻjM\Օ��٢i��S�Xf�T#ͦ��1�2UqW@�����FB=�D� �A�*��ׇ7�{�R�6Ǡ������	ÁX����h����"�(�9;��.��}�&�������(t�ܦG��2���Z�z���R��roD�wmEm��J��IN2A�lw�n��\�~��f�r��q���8/��O����h(�VOx��dH������B-9����X$�t66�-R��X��5�:.�IW���|�ا3vH����jј�A�i�6��N���T���M�}S��N���<e�5gl�[4��,`<����#6��|� :�W�~p��b��
��t����E��;X���ڌ��}�?�^��hN���G���Mw�bBW6�0�U�U7�����ɾ���@�Y� ������X���Ǫ�+RDg��G'	#A�hv� �Ŷ)(OT���Ҩ�z��/�����{�,$��i{�%��(}E.ð*y��� �.�U��]DMs�yː1B:|�c$�ż���JJYŁx���45�%�z`��K
�'��9 �ױ5�A�=�h�����5�#,N,Q��z�KyUë�L�S����|���N�{(�Ru��1� ���y�����s�j�!�W��ʉ���+���c�ʔ�h���4V��\Fx��O���
�4����/�M��{g,+hй3`P{�9�Z�,ʭ��sS��Il	C�[���Y/���sw��ga�A����s٣�c�u���<��A��s�ݶN������.�i_� k����'<�W :�
�2>��j�iC6"#�<�d��%3�0����H�ܑ1�<�J�8�������b���ƃ!;j����R&]�3zD5��݀������0uw!��%{�Y]<��*7�)��Ӳ���&q]�#s�	!�B������&�I��.��g؞�0�V�
.�]/Q0�Z��m��8��v�-��P�,��S;�m�JKh�"����I��I�vQ��z��Ox�?w1}@�:�?�;N��}<R[��(�]Lax8Rz��)��A�㬖�AD�+T�Gz�ɚ/����v[����@=���<;9UXG'9։4/Z�SP��}z��k:�-]aX�A��[�_��zF����G��J���a�Hmm|��t_6��|]@
���//�o ��jB�+s���.��k!�C����_�;)cA�Cu+S|�ّ!��C_��6�Dz5:��2��d�ui3;M���<�m3]��P2h���8��3��l�~S _��\�7����|
�
��(ln;˰C��
�%{etz�M��؆�/��3v�b�	��+�
�^쥲���8�ƾ�ZH,~�x,��Lڮ�U��:&=�����#��ԗm�Օ�q��Q�d�>J���G61���7�;���ӥ];AE�|�����lٍ"��8�f��UƷH��CL�D�U�E�x�1�"P�.��b��}�tE�m(�aIk�ԕ�Ļ�C����c���b*�؁Tg���]����J�#�� ��-�G$\��ot�<y[�F���/� ���8�S�s���o8��;#���W2;w�l��Tx&Z�`*g�z(��a�����1r|!^gҁS�C���v�����LD��w��`�2Տ���g���eAlA�@����s�њfdp������w�����;9���~������:��䊆��BS�����/D��'Y-&_E9�Ę]�U����]8|�]�jsz�?�`R��w�������z�W_��<B����l�H�l�+G�t�[�KΩ8>р��@�00F�3��w~M��[8�8�����J\����J���e\��i8���#T`L��+���a��	����:)P���� �Q�q���.�r����g���+��&
R��l�j�ǩ��b.>�*�Csl:�[�� Z�ۻ������_��J�CI#�T���8\r��b���97R9�
��Dx �猉�Ty��O/�4��T���7bH�-�03cп�4"	�F$�D�{	>6\��A��m0�i5@��&��,�F����D��e� 8a ~u�b�c�ڶ�HX�t�@����ī�V�3=1�6��l��Tp�H��A,6?���.i9�ߨ"f��;VN;'���U?�&^�Û	�\}��%�0��P��%�	��&<ؚKW˵�o4�-J�!ZJ+DN¶y�f�GEE��[��]a��\D���-��8z��W����3ݤ��g����˥2P���B]J��i�),%�c�{��D�!^ُE���<tU.�:MY�YyH] o�ʹ)�2�R@����_�A�j�0��_��d�7h,�3-��2l��Kּ�ǡ�)��d7`o�|�j�Y��L~�S=F�-����4\�SC�kb�M�Z삓>��6V��yXL�*��Z���F>{�!E�
ߑ4f�X���1��Y�}!tV
2_�;��������x��T���a�6o���j����<B��֊��l��Ow�*Uf�;����!�iWyM=I� �����b����2�5��޾��M(k-��2�rt_�� y�j����{j*����%]a�*�F�e�uAei�����G���=g�E�ve��"�����Q�zV�q�}V�:�xFR#𖞣0`}\v ��oĪ�L=� �s�X1���QDʤPx��F�z�}�H�Z�]ԍ���a!l��=�������	��*ΙʌC���Jʇ]�IeDU�As�j��e�s6 H�SS��y���M���1@�e�x�꿐Zd5o�qOg�^cxWP��b��%d�Z&�.E<U�:{+�&�J��1�]!�?Ϊ��<�B����t�(%%|��|�;�� p���$���lNt�ϖyQ¦)���H)C�L����^�P��u$!��ĉcV| �H��{��$�d�I�|:���O�V���Q��1|�UM�xG���!k��(��S.�r�k*�7Wc�>���1ܤ@z�$r'X�����;�0���h}�?���IK�`
_�6�eM� hru?�S�M��G�����@i��9�a2 HB!�d��l �3&���\��b�Y��;���'2�]DA��p��qv2_7Lf���X��U8#���	�{�����`q�Q"3w�oi
�ڧ���8B��\����y�-�e�3�,�����'�۴ �^#�\?a :A�o�D����L�?�CG���g<&(���K�rZcu��^ �7W��ylv`��px��`To(�d�_*��'ɧsL{�A�EYW�Q=@y�0��y`
;�o_
�Cˋ���Y��h�#���3��%���ya[���>���G{��=�9�P����E�Ճ���v�
:�Q��i���W�e���}Sl�'�n8'�P����Q�sNX�"�I�	���j[h���J{K��!�V�Ŝ������[s@F����?�?�����2�ӂl�B�q=R�\8�c�:�Ԫ�;Q'�����?�~"��c�'�򑌝/�s1�GW��qB*�~M�����F��0xM:�]t���c���[P`�6jY¶��?�y��B�Vv�r�b촫�� �x��N���|�Ӌ��}�R�]��~��a�x�.Z��㉴z}f�r�= �ލ��ӌ$�BT�'"չ%"�Ġ�K��|�dH������sA��)���ܮ�PX"��=��}pIZ�J�MʪYAv]0�/���P�׿Tb,Q��&�m>V������m̚�*������c5�n9n�6\�i]��pM�T�|4ϻ)�1�F��8 c�����cy��0I����1��X��KT�0�����:�ѱ �['���r ��>��Q0���2���o�"~Oư�s�e����A1�>��m ����X{��yVO�������e�@��ž�<����١��&	�XMx-������n�[Q���p�����l�T�� FƱ-BV��$tC��э�P͗�M�<�?�S9���u��y �Q��H���X�	e���P���d��/�I2�E1��y
/o=�?���w͝�;i"~&�8v6!�I�#RC���q4/��%~Z���.�Y��Gs���2�CLi2b�%~j�?($ *�5"Y�rD���t;�����~����e��N�D���h��R����*]�> ]���9t	���Mԩ�k� E�^X:V!.��I�=A1��W�9�7���Xr��_�΁4��ުc�"����g��C�u��R[��ҞKtH�x��0+����4�����A�B�^;
q�&��
���Z�7i.�Ld��LR�9��Ն0�dP�����0-�R�g0�����Ofb��k��B�K�d(�����A|���'%��f�9Ѕ<s����^�p�;E�.�~��LP������]�֍��W̦s�1B�WG$
���ʘ&'{f'�<'�t�&ר��xԹGH��=��l��gs���I�+�.�J[��;ik��.�X<�+%����1��s#kH�ġ��޷�A.����q��ur�\I�Z�r�H�2�R�8�����撜A�0�gV��W%hHr�'O"I<�����b�'*lNf�FA9�Z[�B�B <�{�0�A��f2����g%qg����gUY���]���,�Ūe.�ʜμP�,tys{4>\�T����m���Z��,�c�0���7�/���\W��^Lq��KM��Av��c1���o*�;4Uݔ��yιYk ���R��6���G�kW�^_�*�5��V�Ϥ���[p�t�p������i"o�۳�D��za�I:�k1B?7�a��e�A�ݵN�ǿ�/�hF۪K���KC����pd��X&��~�yl:�:����f�N����C`�(�yl#�UG	�Y[�����,tap(6�AL�YG��2��M�0s*���Jk��՚�Wh/�=GmX�SԈO[��Cy�4�HE,��&ݏL"��A��k��.<�Cx��k:�Q\����������gɛ撜@ITmK�#�9L���u�a�R�����_�[�l�J0�o��G��͐$�t��U�d\j����\�8��֣���H�)4!U�����T�8q���ͥ0�1Xu�95
͔>)<�S�[Ai���7�Z]���w����cz�1��^�޵��q�=���R3;Eu;1:�G�w���u�� �ܮ������:U͎�ۀR�:V�DY�-���0�uW/���;7��Z���_1�^8"+��@�Oe��!�L�i�槌h;����k�L{��~�Oߪw/X� IP2���S"$��"4�r�6l�����|P0��s�Jy�T=o�&�z���x�2��L�� �+���p4�t~��=�1��'dvK?k�sa,feB�.JA�"�I�i1��"E�삛��xi�rl���O�'#�����y�b�fֲ�n�6�ç	�UG=�t�����Aː���.Rg�ķ:uP&Ԋ-pJC�ိ�|���5��U�����Q}��].�����'4º�P+���ze:��k��wY���Y�l4X�TA�>�I�-���s���RQ�I�<�5�w��v%��EPfK��!_�K�]cv�s��x�!M�'wŔH% |��R��4!O;�U�yy�h��vr`��U�$,Joo�`-�j�/�V̔�d��u~̀� e��.���,���	Mr^x��팕�LZ�sJ����lY�M�ysAwa:�)G�[A�=z+*B��v�u8֝@l,r�1�>6؁�n/!w��Z�ZQ�*�~��E��yq:HD�I!�Ƨ;�=�/�����5uq�O�.{���8K�-f�h�'����ؓ� ?����2��pzۥȽ�·��-F�f�MYfï��6ֳ�ȁ���Y����ouVo��:�UG���Y�X��>厴9^��d�p��N��]�W�O\��CG�3�Z}�?`��fci���6rAe�+�����5��͈����J֙80oI|�3L��NB-��r��z悶Q߯1������:�}.O"�P]�����:� �a���՝*��WR�W��r�Ԑ i�1���G%�@�C���(�3M-4�\�#��vs1.
����ʇA�T��_�%j
�^T�$Qi�#�A`@u��{�-�ŗa�pwDE;�榯BE.�W��9�'�ItZ���hM(��(���O2iVJ��,�U�ӊFf�>B��I�a9�l���Q��3Pb	��a�?�!��"����d�4RX~�*��0flpfP�B����l��=�����{�
`��g�
G���tbԵz���R�v)١/��9�v��n$aV��W�s|=�
Q�a�!Ui�"����k��N�V
��m~Q��w�r ־�OL��_��b/�:4��ҏ��jW�������
�TC��1Eऱ@��itƷ�@���g��\rG��{�MO`���:,	�	zV���PG��`��_u�9�Y��oI��KD.O��&;O�1�F(j�E3��� ��L��F&=���<)O���<Uf[��_��_GG�g0&�P	��.w�b�Т��E�IU3N19o�d�u��~��G̕�G*�ت:e��)�pײ
.�S�t�i��"�H��Q���{� �9��*�p�.ƈ�u���1/�Ē�
m#nb���P�Y�����Ԋv�%�Z(��7��j������5������O����&�eZ\�"�C��7>�D^��y>n꒪����*���8B[Zu~z2�X��i9�B�G�S\$��j�����8��q-h?"�ŵ�rܛD���l�*?W�@'��T�z�Z%��]�[�[�R�:[���>��}X�l�9��lek�k۱��00K
Nx�����7��3�ҫ�X��C�@D��M�\eL�t=�k){��#YQNc$�ϓ7���H�>�8p�i������L����cd޲�}��d��P�Nd����A(x�.�>|l+����s9R�}����=�A���c�v7M���~�� r��ǁF+���;{ۀ�⍠]	�>��F������{�+(�]��hop�?����f��d��<���|ǳ�vH01�4g���vNXĩ8v�P_�^&��p�Q�r C�҇A��3���T�E:C�LH��F�B�ĺ%!O��&嚏��L�����}U����ŶĔk1u��������2k�b2ajx�taf²m�-����D� ��(.th-��9k���np��|3���]�o��m�>*�@����~�hV�b��M\�.�wK:�_����5#����_Jv�-����BAr~��$�N��9�Ўz�rOb�pϝ�l/n�a�b�j�_�A)����)km|���"p�2�Z�yX#�Ŕ"���U�L�)#g}�+B��xq��0:@�K�0�DG�1��z����jj5�$���%����UgF3$�c�G�������(�M�1��j�p�-Ȗ!�L�A�����D�(�G�;-�*�Ɉo�~p��Q�c-����5��^K�]�Zgc�o����oӛ/�D��|��Mn��� ����ꔺ)��Ҹ�%SEXu��1b$�m�4=SA�|О����G��H�v����]�Y���/� {�������z�Q�A����@`=C�˻�=��B!�\P�)5jU�~��n���~��$������$�m+�T�P!]�ğ����R-i�h1��<�C ��r�
#=n�u���kgWv�毾ݑ�K̈�`5��-�\�ӥ]���Wó ���� lxՑ�i�*oT�{�2�v���M"���5�� 8��s�I[�h�Vrl!N��ўE}����v�zy�-̧�<�f�q%E��*�?s�?����G��E?������J�V�!O�Qx�x��{u�6
���{KE�^�X{ZEg����p�E��8J�l
#�tdEb�f�iT�'���ڑy��I͂�c���V�Pl�Y!�y;�^S>+T p?l�m�Xz���v��v
X��ήm����kb�gẙ�(��D�0�L���iӪzI�E���j�ṸCm׍����;��w�������s�?Ȕ�o5�l�m���,9��]X�K�8��v䕎�@�}�:�l6w�p��cnM�D�l��>��W��i���_�r��/���;-�>�*Td ��r��$��Ǩ�R@k�;�����|w��� ����'��MѬ&��-��*�b#�u�W�Q����s���3R�g��I��`|{=+R\�����1	�����E���{�]�{z����P�l?�X�^8����i5E9���D0"�<޻��4�.�J�Kf� ��K�̖�rģ`l�R(QV��q�`�ڟ�2���ģ3�\�f����h8�ՃN�3GI�m�͉�ά�^bd|-��v+ggP���0���Py��ū�#�ɖ����A�N`��u*`>s9y$�2-��[i3u�.�#(�l�-��$U�sv~�ڤ �^��|2S|�O!d����[�/e3|t���"R��h� Mw�uKČSK��@��K�G��kZ�ʿ}Y�J^����I��?5��C���N�(,�s���5^
%R�`ɪ,�
����5q�>X�Zg�l�;_Kqm��QM�6}��k1�֖6�
�3,?�� 4��s.�'p����{�w;�����P��5�%��c	H, �dJ�<��>o%h+'&�t�W5Up�v�$���Jʻ���zXAXą��	s�
/���.̵�}9A�C纠^�,����2�`S���P�ήaT	t�^����H	�W�!-uK�*��ȩ�D���x^un�֘�f�g(I�v�=��7�����GC
���@�0|������h+�84jm��B H~^G_����-�d|Twa�檤kv�o#��/����������s�*e��\Xy#�S�9����bM��sz+�Y��L�~ Q��xw1ɼzvL�dt���N��8c����Ԋ����O��	��7�daʖ&�;�*��1=���9��MbvX�NY���~Q�:x��A���ǋt΍� [\��́��_d�XO�[��U��@�6�6�ߺx���3��TB��ҿ�)y�/�Y�}>,@�F�����!��JVb��귩��5הt�̪?�D?�u�%N&�(�V�]�F�g�t��:�����G�����:�]��)�L3	�H�1�[�<���C����a&�=��]\��X���'�.'.&�S�\�����	P�}��?9��%'��V۽go"�ߓ���l�jT�,����v(�5�׋��&Fӓ�񋊻-r�������y�}ip`'Ƥ���X�q�� C	՟Րé�oŷ=��Y0H�?��@?���չhQ�tiq�AAl�> ��Ǿߝx ����l(©f��]��u��"�)��6�n�t9��¸cB�>�i_N�ВI��ت_i�m�bo�3h�n\e�`�l�;w�p���Ȱ�\t}Np��85R8�> �8;�re�39�_b�eC��ߊ�uf~i�6�s�c��6V��$���9����z��r�)V�P/�/c	�����Ĺ�/�H�X���k;�4�Ԡj�qs@?�vG�&�)[ɴ���8O�x����/�����[@	V�;�"tv\o�\�7.0A�P6janPIW��jG镶w��$�q�x�9 ��e�G	�aWʁ�'3cm%��APl��i4����v���'�_Q_
�L�I���t��Ȱx.8É�WX��<)��]Ǎ��Y�<���Ų�]ζ652�K�0�PZMm�ͳ��INX39	>�|���e�A��v�rQt3�u��j��T�ύ���"/<�����G /���X�? S'�/12�<\�rf Z�k?*�u���I)�>�S��}J?\�����?�JZc'��v�����3M �
�	3������%��g#[�t'��V�։ɽLqT��4^D�}����n�y�|d)�!ja��1�QgZ|0fD���QK����=��r�w�D��E�E5@i�H'�s3�����SY`�}�=}�Hj�L�~d���j�(��$�-�6��Ղ�7	��;����1b�B$K��i�ұG�X��>���陆�ͨJ
��HG�v+���I���w�q�Ģh��]¯�1$������'v�������l#v�D{�_���u��$|Xq�.v�����:N9a;A";-�||�<�o=�Id��ga���_��)5Ӕ�E�{7w//��?9���ⲕ��Gq�n���+��$5�0,ޝ=#�|�����q^{6��#�+�^l����)s�vP��b)��k�T�I_��o�Q�Y�y���vh��3�Et��������8FƂB�5Mຼ�=�'w}�}���R��t�UU�nUw{��\.�z�(�d`s}�4m�[��X���P�m�k,v�Õ�:A��d�p+��n��WS�TD�u��I�7�"g�'Y������c�B�)s^�t�Y���G�z6��@�O�3k��u��-4[����(i�" U�^�Hy$�5Ⱆ���2�xb�9[��U��ۧ����!�;��x��{G`�͟`��c̍1��������1��	y�(�(��U��.߽�ȉ~E�.�V�� c��?�����Q�X�g���ë͛�ZRl���B� $������i`�����֛��b,�6g-��LO��bs�N��~�eU�wB'/iT��%V]v� ��FϦ:��_�f��V��ޒ�3E���
�s4f��eƿ
����B?�N.V�,A�ڃ���{~�}U�K�etK(?hdv
���Nyi��N�?��*V�-����u��Jf��BL"��߄h�ܡ�|�g_��{����֫���Ғ�{Bx�!����U��p�|�X������n��C9O�jn��J�a��*�NiT$k�,�I����+IJ%x҃���%���^��ӗ.�2���=�C<�+d&�1��2`�V s[=�TJ�P���oڦ%Р�Z��*��ߒ0�5���r�U��p�#�B[՟q�gw8�x�3��S���|]�>�kʢ��V��x��kh�G&�<+����v�\��B�6�҉?Jt�GS�8,ڈ0g�^�����(�p�����~+���ɶw��J�l)?�ʸU�"p˧��`c��2g��>?��ϫ56�k��l�G�0������{?W4e�����o�^��� �����[b��q=1Kq/���zKžx�)Ĕ���1LWg��*EЉ��S�K�[��j�!����	���	D�k�BA�1�M3H��G��i+�7R��D����1y��%c�TR~?j�e�h_;{�����M㹚��4�>��V������[>3��)�z<^��|p^��5����7��m^��f�7җ����HQ�M��N&<�D)7��)f��Nx��b���.��� :F|KRA����3Ѽfe��󫝑�-��f*�f�6���;�F+�ȍ�O�P��UMKFM���;Lqə�j��/�_'�ťC0���_��"�exn�� 3��&U�J��i��(a`������3ɚ�L����7E�俹R��DAD����5�;OcG}��kz���!�ˇ�$�X���c�#V&�3��R4��Ӣ��Yc*U������G��+2�9�;W���g.�,�+�] ݖ9�	�9��%W���*1��n��x�����,vD߬�m���~s��1.��q2l=�G��m��'�W6�r�yw@�U:J�K��V�V���ڰY^�> �h�i���5ރW � ߴ�ᚐ�!�L^iv'8֙�����D���L��[ㄷq�o����s�n_�q�﯄��������s(����1�W����\�l�A�rwy,�@:� �˘U�=�
:���~I��l��,mn����>�hT[G��S�]4m5E�]}m��`��(�P��X��1>�Cw�;�LKI��n��hN9Y�7N��[��,t�Z�?�X�#'&y���_���{Q���Z'WV�����_K4�P��u�;>�so�:��RȆ���?�p���Tv��%�@�ԉ<#���?m�clWF;��ɉ�k��1Ϝ�
���H����ЫoO�7m���p��6x�(ǎ�6�������G��;�7I��ba�rS=�f*: MN�x3�A�[0�J�����H�Dqҷx�2^�Vխ`���h�C�t�Z���Z�N�3Z�{�3�4�ʩ��d@�2�Z_�x8��UmE߶A���醉����rӒ������gv�X�~���ߣ��=_�a�>' ��V����pxx��LŒ� ��+��?IRe'Y3~��8S�LE��TK)�m�$�����Z����K3�転̦Z���Y�g@��Fض&�q��#ʦ���_�"�T �ƥ?d59Nt�[�:k#���^`I'��XF�E6{����2��q�G�*�e���b���;��4C�z�+_��{�~���W_�φ�&q��9:��K]ơZaWdpԤG^�T�p�ț#�����,�;k�����vE&Tq�t���4�g��́�L��>R��sxV	��yi4�j��39)���+�Ş��+��?�	��b Sm{k��=���{�=���=�!���J����1����H&���e���7���g:^V�o�[��p]v�v�E��Q����c*���@��,%��z��K�2���W��-XS�:+��`?H�]�nO�A�y#���ꗙṞK�4,����?O�%�떃.D���
]I�;߅t ���n�݆���~��������4��?���vn1�j_�l�_	�&��(<b�A�>�K"(�Yd���V��Fq��(4*��e]�w��\q������
7%�Thb:���AC��R�.�Ϣ�y0yQ�a|B��J�x�໑�r�˵��8��,�X���ք�|�V�I'-�:F(���;�}[s�e�!?�WY�l���R��p��r��W�93��Y�!B��F�rr �&e,�gT�;���5F�J�R�=�`|C�挞.�W�����l�vb�&A���O�Ċ��]��e)e~�ʋ�9z�1�Om�)SD�#�c�[�!(�����/5��t�x۳ cR-e{�*˱���aH��FD�wh�.�3g^���#WONt�!�e�j��k�#\�z&�Y��jRj5Et�+��9 _���oѡ�&!���5��xM=�X'֒E��\.ĥg��u4+�+?�R�&q[�����r ���R�[Ƶ9!׫N�̴�"g&L� 8>�Ѱ���!�x^��$�x%�L����ͮ�R	e�6F&�ЦV	���Ɔ�8��|5o� 3�.��Hc-Aj'�MlIC���ƀ�$$oP��~,
��|+οI�Cy��c_�o��pxR�)�z�cɀl)G��B�_c�w[\*�����/��=��

�`�*�:��x�D�K(X �"�M�0M?�B�kɧfo�H�5XY�TU'y��.����C���y�q�;��ϗvzR䓰O�ŭL�E9�WH*p�-hu�{9m��kl @���"�\������.�Ck�"E*�(0�tҥ;��+qQG�Yǹ�9�/��g���rBM��=�#��}�c�_�6���{�����W��P�|�B��:�x퉥�,Y��|:�m�O�<�vy��������:<�/Ֆ�w:��Sv���ԋ8u;���.-7�}!�<L<7������E��D�;�+mɏ���)�b(1�QA	*N�[��F<Mk�K�C�ZLJ��,��o�w�&�Vf����8
��wj��(��E�8D�r$^4����rGu�c�gŤ�ӵ7kԡ�}]�]���݀RB:��>@E�ીs"]�2�+��*0_��9[E�/K$v�R���vB�$�6�	�{%c>\b)�h0/�Z��Wb��E�X�z�ˢ�4n��)4���'4�O������g"���<����U+Y���0���0� S��4��L()��j��O����O���ǟ�2[��r�k�ݗT��@� �ehK&I�ZAG*Vv��3�ɸ���(��Ã�@�6�N@Я������ei-~�s�)�l7'�X�8��'o>�������2ƞ�������ç��b�$|U�E�R%���(~�Z ��նXj��P��m��2iO��nYX$��(B;��	0V^�� w��WP�
$m�����5�q���H�Ʉ%�1ǁ%�Sr"(4"����}|���;�ʆ-�|��1:_��/<:BRe\g�����Ё�&�<?#A��-7q�0��ǘ�b���(N�K�y�N�\�o�P+��z�	���@t���k���T��ReH�O���Y��Ԅ�dX�ꁬr������R�B�zb�/�rk���&���}�3�k�����9/�vQ�%g7����~��I�N+x%?���לA��Ss�؛"Mp��{���Y�@�4t�x�9ՙcO��ڋ����Hl���H愯�O�n�GUn!�^�����q;� �l��E��1�}��'�-W�}����6�䍇��������Em�L�9��/���%�.�)�|��zs�1O��p=r�}�ñ<�(�y|�f�luW$v$.��.I�8���-?�ij�s���O���U,C�`8X�,���	��Y��V�ا<m���l�?�K�K2��R��_2��P�����&n6�����Xh����?JW4��D��Ϻɺ�1�s	M�@�7UlQ��hs�FC=�-��lǎ³}�jҰ��ziU�t�vAߨ�MD�BpA��	f��bbX�{�!�*D���\.JG��9����U�D?�.p,��a6��,�P�P�Q����6�T�s�/��^~��[��xfQ�pz!.ҷ2c�	��)��Ag�VصZ�9�E��`�x}��K2��"4~��� ����|�`��;ͬOd���_ש�����R^�^��X�V~Fqz�&$��y-</߫a��D8AM~qeR�5gg^�N��<��P�� �G�0wE����]�{��
�ڊ*wó�~��Bn��z0p�b�աke8��Yq�����t����m��8��n�ņ2�LÝݡ�:q�}�|S�������q�ԡ��:JzZ^�]`^�����w��n��U�V�� ��������b����S.*��H��?蚄g⊗�������s����&����/����^+�?�p���U���`9l�9L�$`�x�d5�M�˙Du�y�f��,%�ɍ�l��A�����w��3�MT�0	'��R;����"�a���7��������.�6�F��]y�a� ���4W��
RLQ�l�^_*E��;߻b�.�s$�"N[�y��V	w �@���^�vP�7#��"������v�p�TDى���hˍ�q�\��1JN��		��ע|)��3t��u)�A� B�f�f �I �����<NZsb6���u��?��BQg���S�$���ch*����9�:ٿ�]�`jA���z+:=D�����c����ح~�@% r-���������,�  B��Mkl�ח�12���^��4;���V@a� P8�܌�~GR�U���uD���	��b-����;�G��L�$j��.���T$��ءCM���J�~�2����/�(e�;s|`a�ng� �[�m�LZy@(`���4��a:r��r��Z�*��-�|W?G%�y�y��u�{� �É�mh�'yV�j� �Ò�t�����2�����ޔ������
1��;�|�C�� jl4����^s�^�y�m0��>��	�E�8eJ-�BnUSy�$Y�)��h>��Yx��~C+�É�7�՚��+��>�#��J=6�jl@hh�]�����Q멎��M��6k�'x����.��l��UM���K��g>�vJ��$����iH���ت6�
!��+f ��s<��t�2;fwAFZ*��6$|��̺��0����Gs��9g����'��d���n��a�4�fXf@�9�f�@�1�q�FX��)�@�H���ǴMo�DB�1I�O�EyTS���J�f����@+����q�ti:`HX_�aì[u�3��kv#�r����\���aU��Ћ\��#�u5KG��]�}
���B��!��,�d�^�H�I�y��"�	T�8�$^*�~���(O ��%��Y1;��M:�i��������ݪc�z��Ձ6���m��E*Z8��#;{no]��!4ה�S���}"7��%��=��pc��M��}>��f��4��~��o�i�1�i���*7�оL���L�A%�1D�Oc������e���(-F�N������α_)�4���C��^�3X5^�%�B��X>�0�>�;�.V�wޘ�ZI�1 2�>9�Q���4������R�_4��Z�q�c{��\8\	�e��9���C3s�Hݬ�������D�:� ��N�z�	`�d �uN�!bX��Ѷ��m{��8{B���|�_�ͱQ�ge.��@w˛3��z��8�Ű12�l��z��M����J���l�[%����Q�E�X:&j<�u�e�}Ƕȓ.|���v�qT{�b=q�o �y;�F�m�h_&;&����7�ນ9�5&��������׭��%n�O튲E�-�v@�����7}��!��
�fr{�L9���[��2��̠���!O�X�M��h~w|c��"��\SX$�IQrfc�.�6Љ�;;����W����R�����N�U�f/��O��` �W(��2S|��#`�X�i(<>��ཨ����o�J�)�s���<���vĂ�O77��a�y�W�2}��	e�81�c<���GZ���3"Gc9�m�r"I9�m�b�X����3����^�����霂�BS�� �kY/xd١@��&��L\s��� ���>�,�2��I�;�N�"�=��D�Qz����U�=f�;�SHϰ|�����w�/Z*C����[Pq�s�V���@���DM���$6-��������O�'l���]�(�pk]�����dӲo��QB�Jf$ȋ�a~W�х�H<�����f<)�\4_Q=^�q�w(��J�[�&���;�8x���zz�P�S��~P��g��3�ğ����)[��u�sT���<�U9.&�>Ò��9�D5yd�3��u�m����E�Rn �~�#���( �K�n��}���+��/ȌMj�%(�l�ϙ��h��<�_W�iO:��.���J�j�?,q�{���?`X�1BR�cțT��67�HC`	�_+V�h�U��"��da�0��ik�5���W�$/� Tk�9f�lP�`� n8�qusi0�'��B�@?�B}�j����1υԵNXo!tEv��`�:چP��V.C�{�c���g��!
-$;K��Nb�n+�q��5S���������D��>���'c8I!���X����w���S��7���"Ԧiih%f1���d��Z������A����	�'�J�Og~�Y;ߞ��pIr�jr��b�+���,���Ǒˍ�"�U|����/}岱	Yc���zI1	
�N����s�����G��X �(�_�9b��+����(�l��NM���,5�N�jr�.e}�@��/����
�}�S\)J����^�Y�b���r�N�inA��ݾ��T���)~)hwm�����&��u:`�ZtZ%E��:�VJ;憀uQԐH���ɍ��C��yTJ�]�h�$nT��뵑s��U �l,~G����?�� g%�-Z�&�2z�o��L�<���qL�攔ʶ�k���!#�D(<A
[�(q:bo�>�X(Tl��$0qG��֗=܆� Ϥh�����v�6-x�E�����$��-����Q�Y3*�7b�#��t�0�`��F,Ʋ\Մ��0r��f�$���3��?H�36&=��G(�lvWS4��f5t�D�+����۪-�B�BJ�X^�t�R��B�a���^Ѷ��}�*����]��Rl���.)�����`�%��ab�rY�ff��S�~P��)�	]�hj��)��)��Y�A�$�N�hDַ�ޒ��D�7Z �w�,���+np�Jg�����[�ƅ*��u��e�ѐԚ�/��$w"u�J�?#C[jO'rY��_�i�t�Tr�����T�:q��l 7��jE�d"F�P�
�w� �W81��5�\MHB5h q�2XZ��D�_�6u��l�{�:����X��g���V�lv@�s[�K��صtd������|�^��7@�M���>��+�/Q\|2Oד�l�.�j��	�Aj��c���},f��+bUZU�DC�Xd;��FQ87���ba`��0D����?Ī���u��Bq+����Ku�۟XMq/�5�w��;"vR%X]+dr�@F�+w�q)� mə��ވV���c5w{2�"z�DpM��괩~�J0a��ިpr�b\�Pٰ1�+(�P��d_�3��i�~��_|�o�����RŶ*����� x
��s�c�\]���ԛƠ�:;W�OV�[�y��5hR���6���H^�K��A����?�DЯ0	�Jp�N����EO--\9r�	+o/j󚀶smvP���I��~�f_踫_�8z��X
����TO�N�+�����I�����>�T��R�@���8�UU���4C���zk~����-B��t�L���ο��Zs�)O�`Kd�"Ȯs�z`U����sHh�O2+��[d��702{�M�&�s�L)��ߢ���y).6�}?�����f摻��v�O�㍅i&�Jτ�$�SG ��<]�� ^��V_y�a|�x�1��i��$�.=��Ԩ��x5��AO^���m�(8���G�$s�0k��tU�%�eM ���e� ���x�!��YC�j���LՁD�J��WϹ�&U���������	��������ĽҞ��M�&/�������ZxR��c��gP(ݓ8ÿNDf&�F����PC��],��.�����w���G��B�K}'1�vp�g��hX4駗 �3��f~���Θ����$g1(����1'���Ta���k�� d���@UB�Ds������)02�$	3���,�.&���й=����f:��ߣ#���a���p~N%23KI$�?|�sQ�JH�����g�*hO��Ȣ���y��k��'y^�d�o�pOތ7Pq��I͐J�BH�=�V�j�L?߫�Wa�q��~�
�o�i!ϖt�L�ˋi�6����!�IR�#���C��]�E&2M@h}R��qMI��p�P��f���l��P��J�/������RL�;��NE�I`��+��]=ZS	{�F��u���m,5������P�Q l�0ye{�-���&=�i�^�/0��La�m�W,L ��,��T�֢�L��0��J�S@cd�a#������c,��U[�C�!�yf~���"�#��c�>؊�����Z��"d_�mmyN���e���
�̙��y�0?�΍T>�	v��g��3u4�FQ�?��l�F��9@�[Z��㊔/�4�,�3"��y�?�nc!h�mI���4�5R���N��ǣg��V^�>W�^�]��o���Ρ?q�q񲾓3:����Ŀ�L�8��iẼx-�Y�Ҹ��H/��s�4���x0&z9Øhb���&��܌pxQ�K3p�F�[�Nt�
�"�wDHN��8B��b�G'~B�1#������n�"h/F��s����+~�6���[P�;�n�L�S�g��͙�.!�.�S���T�w?=��ʌP$��>,>]׬xc�*��.m=� e#y��p`Q���	ޘmTFt�i�dK����{�����8�J��ec�'�������'�cی
���R1\�����i�*fN;7�+!��u���Y��[~�T����3ez~:�b������T�����1���j���~�(�1Ѿ3�xf�<:@�=$���!Ͳz,� P�m_����`�7��1?_�؞IN��<~�g�vșr�n}�<XK��P�?ѡŅ@�����oٻzV��\���̓�|��93�ieS������|XeOҫ��1!N	c_JĽ%W���ܗrqTH�\uR7�����uE� 9l>�3�E���{�+j�U�'�	q��k�g��X��P�(G�����M������<x�>y�<s�p�ya�ے±��K�6����,�(,��J�����zlMT��'J�y%�C�Y*'!+�O��9?��c��[,�ן?h��Q�,����Q[��wN�@ZjKk���0z�������ϬGb��_�&H���Еnk�?�#����t�p^���Y��f�f���=���>��J�⓺��[��;�������#�A/���t|���y� 81 �eN�����3�#+�]_���c�����a9������>���6�˂���t�8ǂ��k�|��}r#p]C@�ƒ�Ve6g���,��O�γxg<W���U�d��f�����Eo[��L�*�׹�˨؏�ڄq*�#��V���u��A�^�d""�����D9��QB�ps^���ჳ��R����������_:A�R�)�|ш�S�i���ₖl��,���{��-R~ֶ��2�26jF�J�-��BSS��?u��z�j����O(�	vw�񼃢lL�8�l�K�*>5�߱d,C�ul�)z_�i�0(P���>Rq���*�G��i�d��R5��k�8��fll7��S��!��Se%�����۝E;��� FI���1JV+<{6o��|[L�ݢ4x�B���,)�%��.	`# ��c��e	�1�4g%[�Fㆸ�h�a�D�r0�6dp���bޭ;�8�F,en��!�
�:T���a�|ۃ��w@Q υ��(Ai�RꖓV�jm��8A�Vᜡ�[�X�@d�i�ּz�3P�2��Qܛ[{�ET���9�1	�wx84�>�y�j��:txҮ:,d39=i[&����k�}��pR�%�9H],A;��V������Tn��K�:�(�.4PD��׸�Yu�
)#9�����"��"Y&��l,����K{;�X�@bqa2��p�ϴB��&n8��4��rw�R�����&����s栃��܊�V�*a����U���|��ۊ��7g��Y�;<�@���9#f|H���qѡ�c�7
¥ ��\����YՓ�� G8UgAKտIT
%薙�~1�a@J�IB{�zq㠆rM_B*!���Rv|��	�bQI��&�YWn�Ϥ�[��OTx針��qq �	���I۴�jI���`�Z�����sNAM `�4�@�)�Nt��6��z�_��^�<4~��{�Z
%��w+F��]� �>>������ܐ�}�z�3������q�'3<��_��!�X�?Ay��Z��3�_�D`)OVe'}7����^<�H*��Ǎ�7_��D���W�y��W��G��%j�i�z}�K*Z������ɀcp���r\��V�S�T��&�r��"B�u��q��\��)��U)�5A��m)]�����'�����;�%)�-ɂdi\_1�I��ҝu{]�Z������9|�^�[;WOH��	���R<oU��07�g}���."A�*�w%�E�3�ɗ��-�;:W��MwPgF��'=�ܰ:�Ho��3�~EʖP�Xj�V��lZ~�����D�V���Z�,z�w�O�CZ�R�B������y��i��Dq����ͺu�w� ������!тGuX�Iqg�d[�?�f�f���ٟ��(�&ŃU�����Ĵ� &���+>�sY��$tU� �U<(&A3��gB�cbM���1�4�l2`
7�����ĵ�F��k{9y������!�ܲ�J0��BƟ�Н#��L!�*<�A>��F��z���k����M�
�_�i��-�,P�{�/�@�.��6�)��WP�Ţ8� �$*I�g�Q��@��_��bk�$��������V����/{�L��!r�0�8���6��X���qK���fp�M@X6؇y,�4/Dp��c� �;l��r�5�1�wHf��[5־�Q����+A�-Q4�<BO�&��U�H���܁�R����r���� �)��m�v(惺k�&���bO�W�-�=Թˠ��w���'��[u����ih��>R��Z�����F.�k�z\[��b:�'m��|��T
���(�'68&���Z��\��-8�(� �L]�y�S�5N�a�U�"�����J�Dxz��ŏ��U~�إ��t�/ltb]���(}�,�mg�<��1�>����mOXS
xASB���j1<O��5�6E����(�/�/@�5��Bx�o==>z�ljt��!ڃu	j��QF}�wD�dƐvIQ��5<A�y�̹Ky�ي��Q��z_AɃ� ��61ߡ<lIƭ�ͥ�N)��b�f����ro����ˡ1� ���s/ ���GѸژq�L_�Q� zɻ�:�q��b�]�5�n�g���͇�g����W�������A�)���Ȩ;�U�B	�{.W$n#�<C84���y���7��}�}u�5�Axv	�����x��� ��'Pw�7Y�'���Sr"����> � ��Wk���vɱHٔG��QM o����a���Qȫb�Y��q�o.�r`���N|b�KJ ?���0!�UzfY��cKb���JPern���r֫��֐�Ƞ����Tc�w�,��`�mi�_|�n��5��*�`��1sc�&TԮw�Tx@�_r���ni��,�j����.,[�Z��Ǉf�.��-嚾
�s*�\dn�X��y��rl�v=�%WD���?�b�o K��B��g$��NЌr�m[5�W�|��9fI �Ì�(_{�d4�CG������vX�4ԉ�ڹvw�����{��+�X4&�� ��<���
D|��{��{�;�d�_�B��xВ��-��1B�U8G�Z|�֯��Jk-A!fI�ﵴ���s�y(��"�)���Q0����b ��)�;��?q����ⳮ���CQo0�`�tYv�Ս�]��7_Ѝ�:?�+G����圝Y��}q|�n�U��m{-4`�������	Ga���`�"����%���R=Hǚ�%Y��P-������F5N�@Q�\���w���v���HrW��<Ү1����)�]�|��O��L� �uS���sg�7{mW|l�g��4jcU�����h~ɟ_�R�q-��ŷ��.�w�{�=�7#£��m�^��;��X�2y�U�-�������,�v����Sŭ�$�I��&���%���Ņ,q���Ö9����Y���-��������`%)��!0P�wol1]�hA�F�>4�SA��E�QH���������m���10D)X-1���.Z���Ω�ƈ�k�������R�1t��Ӭ�W4��@?ۭ�j���)�����K�C�zu��2P��%�6Ѳ޻WUD��u�5T�@�o�ҵH#Z��<K%�>�Njm���C���+�\�$�yE���Bȸ�P����ģt8�:�$mn����4�I�@	�پ�WB�~�=����eB��W~�������>D����eު-[�4]������wב|�U���)́�z�L`Fg3-�*G�$�*��\�@5���&z5��im����	TY$tO[3�vU��N�� �n<�L�SE�Lnm��{�@�࢐����b7S�bp�[F3hx������Z�{RY�h��2�mr��E��W��G�b:5�`� �����>�߼��Y�Z��1�q޼iMm>�쁀���7i?>ʁR�Z��\X�/�5�p�ilk�u�Nz�y�@�����3Ov�a@|�^������qE�u��T��8�u�	���b�y��Q�A�áNeql0�߶���%�� _��4 �L���A[���:�Z�[yݡ �7�S���-)����!��P��B�&�����M�*փ�P��|�h�Dp)����y{�}�M�b�o4q����h�Kg�����L�f�9�
$Ci�8��g��%ﲇP:��p�'g�$����󭵪ّ���C��a�*�; �E7��ë95�=���%*����v� /���,L>K��p���ɥ1[���2���7�U���'�ѳY��@���2w���s��©g�Ԑ�Y���݀�n��>��L��;��:�FX�@U���E���|P��BnM�+�JX}���{t(��������TPl���V=k�b_G��9"ι�bK3��Kcϖ(��wl6���'�We�p$|=��ȅ���ñU8����7�u&b�y�1�E��.@(�3W�.��*����A�;��iK�aa`f��\����{�L�Zp��bΟ�?��9!6is���ؓ~}��Ě�}��.�*�C ���ǘT����2-���oDVd(r�/�2֢��ψʁ��Q����on'b\������6��lp_H�Qil3*�A�A���U�bg�qC�Sa����x,=ӍAb���l�q҃��B nTZs$�H�%�)o'ǻ;�-�i�ix7��/6��SȲ<�r��kAN��IMibp�bWe#�k!vk��|z��N�[�K?7"�<���W�:���Jp[>^��qm|�&W�)�J����u�qؕU���u;3g~!Ce����?`;w�9$�<㝧�Bҋ�g�h�ÿ����-0Fݲ��>�l���H�u��S�π�8
Q��LW�
���w�u+�_�Zo�N|��j'���Z���g�K�E��bG�*3w�/޾'Bz/�Dq>��b0�eî�f��k)�g������n�6ϡɥ�)Lg�. B�8��.6��39;�����Lk�9���Vh�jzJ�P�_�PE����4bqex��,QE����e�pp[�54���S��4<��_�6XedE/i��\?����.�La9�)T!l�կ@y-����` N�"-;6�EjI ���2�'�3RU�0�`�sO�iN kz������A�y���)a����z0�g8된x}d)��H����/�R���X�R�l9�ʳ�G�!�'��@��"&��K7'͏p,4U��%����6yy���<�㣙s�������{rbЙ �筃�h��)�<�8�巜��n��r�������)!pxlٰj���������Δ)�!V�<6c��Q�hKٱ)N��/�'9ήo�D�s�?#_��sW�����'8=�&Ou{d�h$Ks}���3��粈u�e�R�&�9!� (z��t����D�!O���53�_�h���r�	ã�4(cD� ���C��w���]��w���_<�0���s�![N4�'��s�m(�\i� Un��7>˩���1�h�wǳֻT�.]���x	�.ț�/�n�G��h2�O����l��)����8֫ޢJh��G<�:�}�EcShx_�
g��!rs$��&��Dzo��s�O�0�9��>Ȯ^E� ��#?>�m��Y$ߪVP�|��;Dށ��a���@~,(y�#�\h�Wy�Bi�E������2�d(t�a�y�wR�Fj�����FF��j�d'�a5]t��_���� �������f:�5A+�AL.�'�\��w���
���9Ց������,M�ɊO�>����u�&z���s�ި��]�&���[=���|���}��� �Jޓ�P}p ��o\��L����a?�g��ֶ��^9�z�#%G�^��&��*��b�LU5�g)�v���1g&�z�X)���xb�������]%�d7&K�7����kEqn۷�n���T���Z��h�;�s&�t�KW#͋�������c23-^�e5.\t�9�rV�dT��47v�,�y.����@����ӏ���Vp��9���#�:�l&g;Z+�b�"�U�k��`���U/G�g;j�k��um�Ŋg'LFaD	)�����9B*0<%�o�JK&+U�`Ϝ��8*�b��J�B0��mˉ���N��w"�AH�]�t�Ox)q\��e�'Ɉa�[�Ԋ*+C��+���v��~�+��W0�l �izg�����͋I85�>D�kԛh����Y"�DJ*����
��u[�k,8fc�u�89'���	? X��O��	���ك|���8'���d��=�4�
�A3���C�؛r�5�����������PwI�;�pD�a�g�!64�Γs<y8m֏�.}���ńܦ���%5�k����0Hԓ.~eK��61\��N�2?��� ȁUKEP�����%�LO�!w�_Ǿ5bƣ $�F�nh7OUUݬβO���c��xZ%�&�	d�Y�X��I&�rkL�,!6a�b�TXy�\a�wd!�I0��0x%<��!UN���������t�͕T��{��V�[��h'�]�XqA��	�$[���9^�r�S�J�F��>c��.`��":I<�����0�f�9^E��9�F-���j�~���bߞK)�͹Ti���6�]I��7�
:�y!j�**��s�&q�9��k��7L�`7������x�lw�:__b���z88w�(�R��6�9�1o��|��Xw�WF��n)U�`����A��,	��y�N����~b�&��B��=�-���8�Yz3֬G���'|ڒ��Gk��g S}IAe8�@@��:D�v;tOA?��a��
�+��x� ���F{D�c̓:�SQ�3�@�5��Cu�D�fD#̽�b�-�QXU��oX�<����@+,��ޙ;��C���r�����/IX�1�9f��P)z���h{�b�L×�⛞>OO:J��H(=�ӭ\m�=�H/�0�β����kG�ъj�̆����ď�]���B_��kC��?2Rh��<n��]Чl�)f�A�g�pb�LL_hRy��uQ�'��)'�%^����� �Ɏ��{Y�v�P�3*���ň�/�\����a�ŭ� �J^F� ?jkC��(�2F��(*���2T�6���I�ެ�E�����%8{̾���B��VMͩ��A�rn���G�8 �:-�3?e?t�\S3k�XfJhuXJ����q�1IO$��&�jR������-�'���O��e4�����׷�%�B$m�d/I'X�?���o��	����J�*�4��qQ�������Z�Y�E!0���0Z`��D�����E�ȁ@��P��hѕ����ߘ����F�1��Q�K(���s9��'�&�_��dN�}�>�|�cY�KN@zhw�ي�XA�1�C��e�'4����z����q�Ya�}�<kaAӉ��-��h��q��`�Hd�=8�K��̧��9�HKw���F�ѭ=Ɲ*&�����l��{�F����U��M�՘N�ͶI�z�P�s���I��4W>q�����,a��	����P��H#k��j�	o�h����

Ȕt,�tc���,�>�eGЎ4��|�H�f7�� �u?�xO��F��0����xʍ��+�g���� 2��/��2���!��w�]inG7tH�Yb?N��� VL�2Bſ.~��!������<��%�h��^������Ȉ}H�gG�zI�q��(|Y�ƚ���z]rD�����p�����.2�%�Q�z���G�!��EKX��aO���
��}�cߑ��9�ͷ���:���]�y�mr��xzg����G��G�$
W?�qF��)���%�=�cFOX��O����B�*�p5�?Fp��V���o�G;����@�cz`	-�4c�Z�}��3i�	R��d�Ip���{�~8c�/t���)��#���\g����VZ�P!1����}2�	���D��n|��Գ�_�J�=��F�Ց9��m2����h�װȍ��[r�郣9B�^z�*��k+/x�H9�>NI��zz �1!Ǭag�zYӹ	(��I�ў̅_&4D��V�aJ�1�N��@O�ߎ6�V:�ئrs퟿6-�I�׳�p;4z�@��^��i-�7Z�W#)�l��g�i���R�D��8�����d�f��wFF�q�����ۈV�^g<�e������&l�G
lO�����Sd���!!�3����v��W��R:,��U�;����b��0 ]USc�we��h�c�z�C����/�H@�d/&1pG� �Z�U����X8$�8W�ͯ�>͓�]�^�3�"��Š�2T����k63�����]��#�
��|8�fwOo��2��	��b[�1�L6{���)�6a���\r�[�h�k� a$3��������E0k6������RJ�tZ�8���?�Oh�@R���*�O��4IC M3�)��Y�\C�(jp'�G��xf�M���C� �@Ԓ�^Z\��X�ZNgv��Ap������Ox<l�,�'����v�T2D���V��\+�lA���[/A��ntOѨN2�vQ��,��>��J���}�����rm��h���I+�˹{+5.h��2-V��V���лm��5����U>���0�VcCF� ���%��J���%J�6@=i���l n�L~���b��}~��$���"�㙉ҷhj`�
�v��)������ �5���Ӯ�+m��.�DNP����!/ßV����/��{%������oZGl.����&���Ð�A��;!�bx�v:k
 /�
tV���s�t_�fS��,oE�����5�?�}��DضO��'��G�t�P �׌ �X�/��3*�1���K��GeCkP(Q��j�@���^����蝰�����mvcX��<����H��;��(�k�7iY1��D\77�[�=�_A�C;���r�.� ��!j;��c��
�8�*���!�@�H��ߛ�z�x=���H�Уؑ��;��nH����m@��Z��g����M��7Pk}���IY��
������4�9��淟�_a�2��`�P�"2��T�@���	��CY+�+�ȗ��MZ�ʺ`�{<���_�9�܋���IS���'S�Q��{�[ddC��h�+J@�^�A�W�&4��o4ÐL�C�/� ��O�*%y���~s ���BKo��g�=#��Y���l���qBO�CP�O�{�jCK`m���ς.�c$��az\Ȇ���'����\܏�2_�\-Q� ��XxKpC��=!VI�в�E�O�Q��ޖ������X̞��!	�%WT�-8���J7��F���0W���?�%"�&fS,��R��jD��Q4)�s��X�c�8`x\�)� =���}ԗ7��	�iR�B�g>�%�,fy�׭��+������r�|'�B�pV>kiOaծ��H����/(���ׯ�zJX�T (��L�i��A"s�K�^Q������v��=����=̿O[b/Pv�:>ײT~���&�<s����Q=;��E�)J�����)��7�M�(�t��+H3����2Z�\*:?����H�栜�-G���(Zu�	��J��LW��9�(E�|�|1��"�Ou�6���{� �̱3@	{�;�_�|t��a�yvSk�$õ��~�+��[�I�*�7���ݬ�r�����fc9-g)�2��{N=��G��O�@��a�}�����"	�e�"Z����Thjk��56	b��M�w��Hs��8������z �S&����$���;�A����	j��l+q�p�+�������UZM&>��^��5���8��O����3=Un��;E��lo.w�d]�znf�J�_\R.s\:(xs����]�1�Q~�J�.b���IV��t͜q��X? ��s��/�j8��`/�����o��+���/�N*�븕"WN�_/*4���d{�2�F�� ��g�ъ�I^�j�&���C��w���_#vmAiƔwѴXP#����`]�s������}Yu�zf�<s�ntP��'8�{pů���}X���pb􂺄ljd&��y��b�P�����ϑF�~࿹���S8 a��N��^n(�mu������@���Y`9|��]T���b}����.��f�T�Ȯ�m��Ɲ�+3�((̖���Wɗ���`�Ul>>�ڶ�K?��ѹ�q�_��`u��rV&��)�8=���l,T�a=z�=`����n�;��鳕����z��%�����ܰ#Ȓ�����eR�d�I�ծ�H��|�֏?��4
�c���D�ER\��o�#�4'�ػ�_�Gƅ[B5H];�[��o7(���wV����X��nk3dtOB�1�梖UL�*Uj&	�G� G����'�*ȹ!��,J[�#~듭��	��}f��������g��a��ut�/yd�Zm'r�GTo"���f�.#���m���;�ph\�
fͯ�'��U%s�	f���&s�����R"���9IQ@^s<��Bm_5>>ZA��uc�TI <�Z��#���
 ���x�Ӌ�V���l����t��E��� ��m��7d_(h����[:��B=,I��]xxƆ�ҙ�Rŋ��^�J�/��OTn��
��x��$?a�� C��FNAZ��9Z�<,f{
���Uk�E�,���ܚ���!ѫ�#×��k�`c8�%Yoۀ~������k9+x=K�.�zD�3F%`_QmB�du�������e�J�����\rr.��xoN�L�S�Q.?���YĀ}0�]�v��BSb.� �A�2i�j[�KI
�� �C����k�-�� i�e�c%�v5�D�p?@qM�q�*�����z��y'=X�\�
��A��p���Z�c&:��a�)��5 �ry�^J�2��ߡm��0�vinwU�c��5����C�a@%��N�Ɓ�%>h ,� K��KB�e��y2�t_t���B����y8��dL� .$jO�}�����q�Bk�m�R_�rD~���a��㱩���2�Z�WY�*������;W"v!�F��� �l2���b
�iV��VPRa�~���M�0?+"%�(f%R@/r}�j�� 6�q��Α���s��+�`��E��ڃ�����lv�iި�$4��^��yPt�����ρ����:����9�w�T�t��h��)|����f,���a�sY���}�)����`�'aKD�!N݈�,�J���AW����0Ō���`�ml
ۡ�@*�0�*��%����`h!g7."�����Y�i%���X��x/��_�:�j����aky��2^�|�41��D6va���(�J0A����J��N�GfX���33�^��/5$24�Y\LR.��:(.!��," �>�����데/S�'�}����7�܊
�u9���{D�� ��2N6��ԃ,IƴRBkn�����S4A�۫8Ch�q\������ �_�76B��a���j���e��-�αY_u�h���S�E��G-�NK�*��;Q֨X D�l_����K 	)ŋ���vzZ���G�̕p��Ţz+���ѱ��V�������K75=���r�2ĵӸS!�����`�^�5� �ۋ�)�{M���l�HW脙�V�TK�Eᖡ�y"��iq�!t�F��0@�oH��{{S,,��/-,<Z���y<�x�4����>��J2o��y䉅q�Pa�nR�>Y��q=*��Ƿ��r٩0'Zo:��U -�#2 f?~��D���<Ҫ�p�*b�K[辣~�Y�x��c�Y03�5�#u�C���^��n?�^�,��U9�e>�����($��]Y�6<_���<n�Z����2���%96��t�9[�A���D���g�X�]��S0��V�S����/�zP<���J�=i�6�㚀�`�8r�+gp����M����DT3S/?&aj���]��55�\
��d|��Z�sA�h�e���菎#k��)}4(:)3�����-�NVl��G�<���g��C�U�t�%}+-˻jfhXr|喻t�qS'�H���ɮ��_d��z�߻�V1H�v_Cv�#QV�t�َ2Zhm�����ԿU�K3}��|'�" d����tk��X~WR�H��^�7Sy���L`>��5�ވ�#���@D����a�0��&B�nj��ٔ5��$6v�}��Z��Q)3YuS�&D�Zg6�Ьp�{�1�m�����ǣp�kf��I%��%�