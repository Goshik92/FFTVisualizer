��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M��*����g#φ'����T��6%.^f��8{�^v�wK�T��fAN(.�oC�Yt���Ao�>���� �h�*��9礩[s�Tj˧��Y���oG� �'!�D!�#S��E3@b����}��(��ѣԿ���:+��rYV��;��6��!�iG�{#�Rݕ_����JkK�ݽ4\�(��.*�[{��+����3J��� ���J�S��pթ�`�]JX��X(EЊ"����sZ�Бx���
�Bo\Q�t�����vw�ջW����ccσ�*^���%l���N�rd�!����Z�q0G�nRu�4Q� ���������㜕�f{$u�6v���9,(�l�Sj�[V모� 8n1�.� {gwi�S��������  �E���Ê_b�JWJ?8���5Q`��b��$Wp�!(M��=Q��ӈt������SH�j��$�VL�d66W��#�9aԠW�okk��������?�4ёK���S��x���a����!��M�: T��Cr�9g���=�O�wz`�����Q��
��%2�ÿ��M٣�-�7��("%8B�9��if5�$�q.���A�@5���$Yj�)��)��7���<���3$�XN$
��ս��Y��#���qzu�)�L�.%�z����>F�ßMl�_aI��0ǲ-V�GV�_�8�Z/g;�-M�/� ���A�YY"���o�{a�I3��b�/��>XK՘�WX����"g<�����"ꑽ{��9M�ϼ�pP�z_|�	�aG���������^��C��'s�3S�+��!����b�lA��+naʿES3p��ޅ?�%I�4��Q:æ��R��?�zp(e�:��·,,�%�W,��O�\�?,ͻ��Aw櫼�	g�Г������C�ЏՓ���2{��f�E5Gf��^b}ȵ@�4|f>@h%�C�h�,�ݪ��h>_&�ijOί�S�9"4'��BDlRSJe��qV����V�J��>�(��|�(D�ō�&A���_1��4#�o�����z��\i	Ҡ!A�Né�a.���pqi�C�\׏f}���6)JY���G�s��f6�C3|���</��]����1�����L���.4���m�����1l�|6��<�C��d_v�l����x������Y���^κoX���'w���4��!VD�"Eî�=|Z��P�Z�l	��
����,�V\#�����TUI$?9z�2)�h������������b��t�쁝�x!�_&�.n�����ȳk�5���UO����0/sETNp�l2�/��YKX�	w��� 2F#i9� ġ.�̇�f��$�����4����J$K�˗Kv�#yr�T��_�X�li�� j�hU����($De�Rn~FCo���xZY��㫬���F%!V��6���,k������<�ֲ��?��/���;3��G��狟ZW蹚�(� � �)l��R4�Kp쀲������#rbS�1d2�!�['#Hr�p�/F�O5��sD�z�m�<�P���XZN�y(�W6b����4`���}0{�������\�O;<��>T���*8e�E��}1�#i
G�������;� �˪��h=�*�[��r r��D��xa�
;0�Ll����;˥K����6�O+�#�� �M)M)-C(�D�QjZ̈�t�?Y��}�{�����!���uCq��G��	ƝA\��Ǜ�^t�ɳ5٧���c�Q��p9��jD�ۋ��15���(2�P@��w�R�㳀APwS��3N���Z�:�ny�}ڲ�}BU��#sk�zV��\�A4��";��]}j ������OF~v:��*庽9�4���2�#�߈�Z�a\�A��Q�h�I��c������������GЄ�[�/����"�����s.x�h�X�r�"{��.�M���7]J��׬ƀgd��Cߗ:�C� >��|�J=9 ���s������3
�{��C�����a�и�@.�@�kժ�(�pǪ�ch��pk�����PC�,[�TP�L���A(v�`}Wg.p���:}�Bm���]�Zϋug�!�-m,�1����SG�K4������k\�� ��2U�]c�aI��M�����V�
U����vOJ�"����a��B	�I����7f#Zk���=�z[���
���0�ލt]�<LT��Vܱ�=?թ��Y �F@B�9�V���6J��tԁg=��s�H��i��(\���dt�k�{���r�U�>(�ߒ�Z�8���'l�L�e��,��W7�|' ��9-��ՆD�J���.��ٻ4��ov��n��^`�G�eŠs�~@l��ٿ��'�?n�#�=����l��3��.CB�Q�����qt@���;@u�J�
��������@y�(y�!�u|Q�k�7NV^�We@X_��UFb��<��@F���r� 9�t���ĻROX��{�W��Α�Zy�4M��[n�C�9�Mt.�*�tN8���?�As��,�|\��pb��(�)��K1��N"SK�y���C@/=z��˦Im �ۅP+����O��}?����§,42����{\����ޙ��\�v��x�L�2H�������pq�k����'ſ�����N����݋��J�9�H��.�H �e'�z�f�]�T'���v�{�A�~LJ���DqT|��;C���vz�!"��wk��Bgt
��U���B�V�W�A'^�_����y!f�	���m]�p���`���n�MG8��;�P���M߽v��x��Q�H����M�y��D/���dU�^&��B�������=-���n>D�ܤ���0�F�w7�D�1�M8,�2nbR2�Y�'oe�?Z!��w�{��	a�>��}��}2��BHʡC'6k���O�2���o��`��-�r_���t�C����9'�ێ�R�Y�흫q"����Z���2�
	��)c�0��E6�,EϮ�g�i�v/�HUN:JE��0eA`��T�;����Rk��ܑ�rt�?S��������$
�_p�;�A�t�Rޛ4#��Q�,;�?1`Br7��O�@�?3;�6gh�)���t^o����hT)X �j�;a>��Y~Dt����+��42�A�vvҍ�����Th�&v��!����w�K"V�_�,�@�.�em�͒|�y���z�C���Cޱ� �G�ENs��P��<�*�z��}H(��x��wXf�k���n>ݵ����.����fnХcm~i��4�88z�
T��@dʗ�/�0�v�Y�	R�q��)m�4b
%���S[
�Ӳ�o�,6bf%P��0���O�cדcw1K���ç��m/Mɐ����r���LS��ӛ�y��ro�$�ۘyy���ڼAu�ƙ���+��iq�����' �~��z���ͱ��A�ا��$s��.59\�A�u����&u;;����w�h����ʾ�`�}��'��h��B�ު7uL�j^s�&q	B�E�[�G���u:����_Y8�\�s*ǃ��?��*a��J���Cv��*���u@ER'_A��J��!��-�
����ːd��W����Co�E�g�w����w��	v( k� ��V��^ I� (���^)��N��9k���X9�Љg'�|�P���&hsK��f�X��~�,�� T�Cf@G�Sx�� h��Kr&/Z�%q�!$��T �d?�)f�_&����r|�^'p�Ѓ!��X�"p|���N����мOh�_�'u������zn؋j/^��H���D�jbv��M����5N��=�s�*0(�x�9eׄ�g�����#���-|q�yPѦ0%�R��"���5zQ����P4+f���mZ)�ևL�"�1�:O�<q����k�$Lk�M�����4�Xr�Y����_J�~��%�sʱ|bE���;v�3� �)"�]���[
��ǳ�$3e,¯��6ȓ*ς$�]�$��������崷���s�y@�D�a)L�B��n���fK4�6}�5L��U��y!�"[f�u��J,�p�+�)9~l%y�0	��7���En�B��z ]�	�i��_U�p���\�Anh�%d5�G�*n���˅��1��ֳ���<���{(�zapS�S���>}�K�����Ti�/A�7) I���
����/�9�WH.-L��sEs���9������͇;)��{���սA{ǀ��2��u�O�E�(�aw���nŷ��|������P~+$
FO���
�8f������d���@�7��G�N5�C�{�
٤e���.���WQ����F(�/ǖٱ+�ͷŢsV� 1��b�Y"�	h�4�6�p�o��7�	�]a:��3�WcE���O��t����"���T���f������{��v<�W�E���*$S^I�# 83i�P�;��Fp��!^_o��(H�-�ی�`���2^�#0�z9Ń��з�oF�9� ���V8�pA~����~yP<��(S�me��k6��W��2��k.�t5~Ă��Y�w�*z`��V�w=>��U��=ߑy��V��������k���j[�m�G�M�����bq����U��㰷��~��{TY����&y��k��<a�-ڠ��c�2�2=%ZmҔ� �W�z'��!?�e�{��DV�����n�	��6s�!�f
D�N�p�^$�
	xz/F�_�&�o��Ưp��S>��^w�R<t�q�y*��\�Ѳ���Z���j7�Z���
@0Iw�L�K# 4��!k�y�(�=!�9
r�p��8'"od��oZh��߁�ﳒ�;q\�v�0��\ϔ\��?�l��p��
������o)*?�����g���^���U3�p�q�� 2HS�i@j	�"GS���8.���Z��^������u���T[����b�R���}L���ұ�w�����E�;-C����vZ'3���t�>&�"(Y�:/�+��FV�M+P��
��>LRr�Ēy5�|U�R����ʈ�qw�AA�ǟE�'�p�̓��31̟������P�C�ypЪ�Uðѩj��F�h�{�����).�b���C��V��	�<}���C�K�8�`�4��ܶ�||�vRY�����^��_���4�!�-�9����'����c�_��:v��Ǻ'C�<�׷-���!��A��i������Jӂ�ӾL�q�C�b���E����Q������t��9���`�{��ڀ˓����5��ş���e%�������Hb�8��!�p�(fBq����܎���2	�P�WW��B3d�P���#W5­5'%�y�EE`���k.v �����{Q$�Z#�<��_��VFcoK��Yp�6\4������)k v�;��T^�6yE<���N���F��ڌǞ#��!�G��n��FD�.~�c�J9��YS:q�lXӺ��0Mp��夯3vܗ��(�����*ts���	��N���SS���K=6���?�K1!��̎�\��NcT.�l�举ߵJ(]PW*`�?pjr�C;ex:���9�������`���� R���t��̈���E�̺��ȴ�S��@.bn[Q1.�4�0��bm#WW�$Z���~�����܆�1�B������"{WX꒍R�7�9w|"�g�c���͡=�](����*ܻ�Y�j���3�-���6������"���I���Q�7{u���/�؛�"O�Z[5ڇ	n¨ zEY����_&���?�#�&YU3��-��p��d̷[4&������&?����w�l+�W�������\o�RU��Y��ON$t�˜(���5.o9!���ޚl�][i_��Ft�,���Ʃ5Y�+��2LE�n�cJ��_a�~Z�)Oz-{_h"��U��c^��v��KZegA%\X�v�;'�A̍��yi����q�S���M�%�J������1���L�Kn����^��|p�;M��+(#�����K�uY1J��gIyUy��\*�w�6��_4�/�lX�YXS��.?ӄ�=�l_H-��f��W@��2����2���|�rcyϵ���&H��h��Q `Ŗ���� �6_`���������2�5�������;��]gu>^[�'$�X>x�N&M��K����æ�ӄg"�qb��p����ӆm�3����!y9�7��ĺ��n���E�ov�{x�>��
�Q]Y�
H����t�~.�?�QLO�
W簬UDs��j�RCk�	�Bb�2�1�ȩ����zn��/#xI�s�F�ń�߱IIZ)�a�P@�zH����J� K��];��c���3�;G�����!�qg8��2��WZCؖ�G��,����a2��kZw��v��G+)��|��Y�k�5vM�s!
��`b]�";��|`��!q0��<}d����$��� �7If�7n�ƚ ��<7�X@�(ѣ�©l�Yj$�:V�6S&�c7OS����#y�M�gz����I�GklCN��4�F��n��2�;4��9S�3����������z�YTM����L�,U�,p+�O�Q7��?�����p9�T8��	�).ib� eQz������N�MV�(��\�!���w��o;zSPu���;�0Z���zyA;�6��h_>�a��|���Cs_X_����,�B�T�S�;�=Z�C�@��5�c�!*�����ƻ��%\O�6��:Y�l�������#n�� �����A�G��y^�ghP���a�6ڈ���b*f,�;�"��$�M�u��r��@<�ǘ��w����w^�fE���|��n3��D����Ն��wK
/4jJ�k�퓢���}��?��i��������a������A�X)�E�����}}��_���*�罿�J��B{���Y����S+��L�UG��Y���(�v��\��u'���#�}d�W�c���\����`���⬦,:��"�L��<\��nY�n�	m;Wȏ2f�qBntnǈ5f�B���R�xVD)�d��~�I�8x���(�jq��^�5��9.���U���g����A������w��2q��P0�r-���1x��8��Y[��Z�*~h�B-����=�g�,�1Dv_�Z+/N��r��	�����Oպ�/�l�r�2NC��`]}�`�-�}M,5Q�U"�RD�U)#�G��͚��w��g�� ����'�w�H��T%�Bt6Ml��֗51��C܋�0�-�0�6N�cX�_�>�A�
:2H��ư ey�w��RJڥH;W5Ah�Eט]��_K�œ��ac����*����.	/8�k�9�חy� �N��
����k2;Y�(�$ղa�s{BزRO�P���Oߛ�Ìuأ�o�@1�����O��� MV6w/��Ll�hq�a%����x�BN#����dы��	�_!��,k<���¹��%A�n��41��8�u��Q�Y�F�.�3�$�-U �r\�Y����L�qWSGKvv�l9����|7Z�2�R�[��g�7��#G�M%6%W'�A��g�����o~��&cS沌Lh)y� <��(X�>8�By�66*)Vy��W�̋�b��ޘ�ʵmcm�]�$Q�|yἲ�lN�d6&�f
�f"�L[qNK&�YG|Qs]矴Y�ؿt��Y����/��.A{��kW�g|h�>�W;o��6_;����g��z�����98��3��z�������y�Y��3����0��Mkr�1<A�T��k��k�n�!���k1���.�;�t_/��8��$�J�%e{-���˸����z�<�q���9}S	�N�<�g�����1r�k��V�$\W��lE��:�d(�2�V�}Q����-�C�o�]
�93�]�,��+Кb�X~ڐoON�Y�f��ro�}���A9!��ǿ�R0�U����q��e6�|�)�P���ڞ�ف;i�fy��B���$��YH�̔92� ����os���J���������t��=;y�Pg��2�,V�9l�{h��Xewxy3q�b>�{�eC%@�#寧 ���w���D��� 
���t�Q������;��G��s�It�\zz�)�rgΒ��Y"�s�i�<�t�£i5��m��/�V�{��@7���
O[�R��M�]8�jh�����|O��ܵo�� f�@җ-GZoe�:�(�M���'�5a�K�=8�UEsen��KA��Sb����ƥ R��r'C�x����Tk�Y�)��;���UFPD��K7ƮLV>������v۝��M�8�1��q]5F�H9U���6ĝ�w�AX��i�;U��a��$i���_i�#	U� ^�!})��D�u�;�%R��(�w���Id������n����SBV��7?{���n!p�0��\���v?�t��q�D�t��5�R��
*I[�h��g�vxdH�[���+�o=(�^p@z>�����$�K߼P�\�py.x�1�4��s�&Duop���ѓ�7&����ֲ�z����:X6Я��8�ܲ'(�khy%"�]s�z�3���ŵk+_XM�"�=d7`���ם5�)"}�D�G#{Q���s#�~��^�)��4��^�36,/C�q/�H�X�������+nj�w±P�7h֔j�V���Ih@HO5�jE<��R�T�
���\�NG����&Q`�%/����9y���B���t%t�]оHRu���(rN���gr5��:�)�"/�c7	��NT|m�'�ʨr��.!N��05�AЏ�̼��� ��:���m������Du�R�ږ��@$��A�"��P��*le��*�msu4�гL��L��g	ͨǟ�?����\>~"h"Y��D�_g�����P���W�������9��&*�~�����>�n�:�H_�Ӛ�w�u�{=���d^EIo�3��p�|�	J]��l�V��AdӶ��hҡ�c&؃�h��ذ8���	Ȉ����MÉk��U�T���b<�$Ȑ���~��z37MhX+7��k�#��.ry��zf� �atd��,�BL�i���wl��q���Fr�˅���E��50����@�u<�����bFUw���~~�g�r���S��M�˓猤*��5l*����?g ��,Y��2��.U�p^�sJ���z��-�0nᄺN�;<��m"��4IhH�i��h�w��z�����'��Y�b�e������4N/nK�GS��Wwv��Wa�FE�8����$q���,<L+Cw*_q_y{P���5��k�H��L��^HJJ
"�����#o�U�4J����*�1�ZG)�H*�C�K:\��y}��� ��&}��:��S�f
p��B}����J�JR�ڥ݃��_����K�9��
��&�O	� 3H ��%��08I�ӊ8FZV#�nӃ�6������{:h�H��
�R�\������iKm2�B��%�`m������Ҫ��tf����X�/$!:�$��eM��9��=�0��?�yj�t}���Q�O��0S>�x��erZ��NaJS46��jߝ�
��_����>b�l�������[�������7n =�d6�cx�4yo��L�Է��{�5���}��>��Lq�@�9�ه���$�N�Fܶ��w��~/�գlo}�z|Of=]-�,8pt%�Hz�w��Z�+�b�G�F�Rs���׳~P��Ex;z�Z�?Z=�o�������G�7j�9Go�#�&[1��I�ss�:�2���!q�Sr̳p���j:���D[����o[��,�����#snG����/}��#s��}�"��KR)�o�U2̩�����"#'�fy=�)��hx�e��l���gCVA��'�|�q��'l�"X�L�!,V���Q�4�X� ��Md�B�]�_���*���<8p���FOa/���2$�hפ^s���SQ���D���O7<F�L�5����s�u�5��j>��T^w��5Xq�x>�휲o*�����[G2H"<n����b���k>Gy[;�ӞNe��dV:R��,��~#Ĝ ޤd.xW�׎�c$7 � ���`�^�RG���5��A�a�.�;d���/��g��I8�y��i�z���z&,E�Vl,�q�K��ln��v��<"HR�x�ox}dyH�bf�b�Ã����u���$s�:g��;y�~{[��ȳ7,m�Ȝ+:ڱ�O��h���FRu����z�d׫f��2�O�����݌���F�6�"w��3��[W,(>���od��c�{��~�NM��� �U�eǋd$[�!U�n�d�Z��ɡᏏ�%���4 ���kc�?�+�6f��,�//�L�EEB�p<��7t~�D�8T��`;A��.zg�y�"b�m5�P;7@]� XXJ{M��9&å��DC|�s��u�����/f��Mg�:�oC_�%G5�s���鴐���l���Ԡy20̰�&-�P	����K7��]����=2f�,���5���蝚I��}���.�P��K�vl��E����Rs����1�$���X�8fk��
65lj�%�#A�6E��E�,��I�c����I�Cc!A�7�`�x.I��iN֌��Ҭ��<��l�e����-vg��Y��n.n�s6��e�D-
o� ���/�����5&��7rX5��	+Y��h�Oa��t�mݵX�Z�c��d?o8���� ͷ�� ���vo�&_�{�dad����7}�����ɟ�
Mz֍j����l�_7�T�ū�5>����
d�8]b9I��)�.<�wz���`�y�čbu�� ����̎�.�3(�+�irV\�q�l^|\`43y�H���׊���];�_զ��PM#�-Z\[���uAY6��A�%�B�K�`�3S��P��0����۳_�V��"�jk��E��[o� S�:�	��S�YSR�6���@n�80Y��[n�[J�fi�_�H��9]��x]1LH<�����i� m%�|��o*�n��"vW�8[E�υ%W۴fr�E]��qܪ��8�vk���r�1k��Lp3�����XZ��{_�ÅRx��c��ޚ�up�@���/h�Ĳ�2w|W�u�TSCӼ�~( oC����T�L�i�l�Q>�v�8��w������e���=���f��/�8�2+�e||�E� ����0	���s�J��N��$?lɠ�!
��r)��U[q��`D�a6;�b�)e�H(��Å}�X���I	�a?7&%p��|�W�ϕ+h�#'1;k۸#�}�����G��
sTsE��(hp�����l���ہ���F?��X&nifx���P���tp��VsH��{a��o�^�>l,gd	��;".���ɮ�m���57�XJ;���[
�/�w��hg�vP*�¹=�kT��Gw�x�`���Օ�QWu@7b�Zkբ+�>�A�?ޙG�mq�n����K���4�#F�+|L��Was�j"�ߦ��]�`�H�ٚGs�����Ov���H�(c�)*��V���/,�
ޱɻ�s�8�x.t�j�H1W��n;�ӂj�JO},�:ZZ>'[[o�%RD {i!��{ip��Ϙ�Mc��hOj�S�Tav̷�ˣW�[%9�@Ǌ67�s�A�̌�|rx~w搫�Q���z��<��'�_���lKӹ7���Z�&-3�e�j\e��jlIo+G�G	���V-pN�-Axg�X�h��1?Q<#R{�ڍ�>A�!�q�(���\F+�*��)
� 1}rV���e�s�
k���.�.�����,��������ro��$A	M�i6��q���Zf5�X�K�[�-}�*���<u��K�|y���t��R\6�i���4������X�mB$����w���\�ʭN�|N��:ک���f���3 z�	�?���V2�2A�`���]�Oٕ�)�� ҉�GK_���Y��|��}�V���u	4xi�(�96�0 TR� [^!��P�@���5�B�����PnH��H�/��:��os�v$�rfB]g#�7fP=��ni�?ߍ*���
��Fe�5i*�*ͧ��M��x�����{���Y-���p�4K+>ҁbZ���i(�G�Wz��yK�VJ&`'�BЮgW�7�,E���8aG���6�L�K��5֌)� �q���I)��Y�[���v��sh�����PbY�F�^�["t��'H��M�'3�1�l�P3�+����6d��r���r��R��0ٲ뷬�=�)���ŭ���k;g�+��5)�k���uм�g���)�-����#��<Æ#��=P�T5��Z�휷���z�R�n��R�0s�YD%�_=f��`�����m�VI�q����=i���q�l�n�H5��oc�&�5����VI������r`��LvI͕�m����̻ب�R[<q�ČZ9R��.L]�Z������[�K�۬ć?�`G�j��7V�DFL{n4�F�:��sRӄ���:.�vo3wV��x�c
���g6:w�����������R���RzH㨪�x�BI-&��H=�/���8�L12����.�%6*y�L}��@��<��O�_9W�bq:ܡ��`l?�D���6��n�� T�o>c2{���i9��gC��p}�s>�
ũ�,��;I��|�#���Y;�ה����|5N�n�8���<%���E^��F48�97ȗ�a�w��ݎ��Y��l����ԙ�]:v1�ùJ��f$:�چA�\�K��L#TJ'R�朩�O�8Y~�Hn����/xc{ٙ��DÐG1I��-��x�ag�9��?=	���l��[���	�z{@?�r2|���:뺎�}m_��Y*�&��c���q �EP��	���rS�����4Y��Y�b�sNk���HT����T�~j<�:[[������7 D
�u�S�D���;��"�˸��,�	���	�rAU�A��BSm�#��/�C���+it�p���+M�t�G��X���������l�Y��x�W�a�c����[�OY�v�@���=��Y1(�70�Y��{��.�����ΰ�M&��[Gj�q��|���kgzZ�/��<�3f�U@�@`�&,�ّ�Xa(�Nx*���J�"�;�wM�&p�����KJ���V��k�ұ�;��¾�yѮ����d�1���Ѥ�z�t�W�_'�� ��f�{�ڝ��P�7"���7�>��G�G�6����.�4
*m��ᬧ��}h_h(���!�bKe
Q��QN�>/O�p�]���j���Y�5����:�H�'0��
�٥������p���`��H��_Gѯn�ȋH��Rd�/�:��O>�H)��������0��>���W{ �p�
��z*�~k�9���h��r�#��F��ExR�{.ä�+G���۩�i?�0RU��W���L�:z�UQ�1�6�[ۿ��r�c�z�����p��jCP��!�vY�M��ڽ���uD��o�ubi��6�8w}+��ű8��+YZ����pk�k�3�c�j�C�&�z�#�˿v�̳	��X��AS�> �9n6��}��+���k�3-	�t����c�/������<A#��Yqb����Ի_k\��G��i,���0��_|�/��@ٮ��nN7��x�]W� t"��t�}�%�]��V��}���*�p@fd�������b�UE�$��0,���o�q�U�r�o��?�n󂖥W��5��/�pR�x��Yr$/(F��0v��=Ǻ��g\�"��ķ
�&��Ux�|>S@�+����6jA�)a
\(^֤��ϫ�����gO����`S�R(�mM��ɚS�|�L���U	.?���-6K�	��\I�T���3�^jƖ���+����3nʠmtPI���3:6OpVV�*���@U�� N�"$\\��L �g'hQgj���/�튬):E%��� cO��N�-C�a��g����Xw
��\���y�'D���z
:�~����#�]�����-�kCb�L=��da�֏��H�)�"b�)�aA+_�8R�ҁMWh�V��;��(9@�C�h������FS���nG�Q=I����d�{v�%X&;����0QλD�͡
�bɴ���?EJ����u!������2 7;��2��LՈ�&u�W�d=����Y�
���C(�NF��������ԕe>~P3K"��S��u�R�$Ù�2���L"�>�	�m�Y7�KshV�t�<����p��YI/��[8j�KDJ9U��m�Z����S���Pn��\~+>��*Ar*��m�?<�h����8�4��k���K�(�7��mp���D�	ң����`C�@$rj�D��p���0��O>H���"Fo�V{�1!R\\�H�,)&�&���G��J0�$NA_'����m�W/��	g�>���>�F�;��>�>�'�ߩ����M�����1����#�O-(�2��[-{�t��ISCm�h��Ӡ��+ ����{���U}ǀ�^���Q���܇T���y�ꬁ�毕�Ji<��G�s�����/.���c`�DD��digܿ�|4~�B.���������mu������v�|��DL��x�`7���ҹ,�)�^IR�7�އ��9=
1I1�7���j�覷��UBj6:��w��_�>�"�3�R�λ��#���#�#{40���\-���d��Kp�y�.<���CF0���,."d���Q�?$��
�|^�#��6�##�ܩ� p���C��a�c�h 2^WL�l��:�;�*
��g�11$��N�NȌ%-����fb�
B^y*�Y����+z�W�xI�ap2�ܮs|����R�*��͖�ۗG�BP4G�tZ�Q�J�W������.��y�������e0�\ނ�u�A9,��m�wY��åV�����
qHkg2l�]'�մ�M���>�q�A*gf�`�_����=���ڝV8����U|��Ӳ9YM/��3����f(2�>To:HWF�)�f$`n�E��������g�_"�����Bw�p�	NE�L T��W��Gy����O��J��σ7��*c<(K �r�w��1��Fǹ�_E��Yve���?f*`�_�p�!L������l6,�P"J�[Pb߲��]�G*9�9����ֹT���������ȡ� D�m�`j���fslz<����%���1%�H叺�>�n�:�G��x�Q��<EC�o��2:t��RܟP�EE���i�Ҕ�˂�=�.`���Xa��؀�T{�8���i���� ����;�b �ȗ�m���}r�( u��q�Ԕ�J�_2��'S����$b�VS�/@�<j����a��(�H�F9�m�wDU�iE��	z�כ$�4��ힰqv	@����-���"2���ȭC�T!�!�3�Ĥb�ƛ�N�ў�����w!8T�W'^���B[&�\JU�a��'-v|F	�G�dpe�&]NVH�uzc �( r���I%����)��.��﬍�L[d��x�X��1@���	_l�����@}���mϟB���)��#��+�k����T+e�Tp\�+�ւ6Ym��a�)��1d��7Y�m�i{g��H�_�$m����z1<5��j'�Ѣ2^�W?�	hZ����W�f��ʺÂƕMRWQHkk{�w�f�����kJ�(�6��g�>䙙y�==�v�IR�%��`��x�Wi~�Y�rm~��9J
���'��l�yY<}���?�!����Ӑ8����%�e�.|hBXU:�/*�ju���l7"���+���2�5�f�4ЁP_�c`��A��g��\�C=��֛�U���f�e)E�we����~�k2%&� )Í�ӵ��W*�^2a�"�Ի!_���ޓ�l��m�-�h.䫄�W������Т�B�ꏖ�d�%[�{t�P��H,�P��6���I���\CO�fN�o�����G���, ��X�Z���r�Us��޻LN��7�@ÀEVB��0NXmoҽ��,��v�mC�o���/����:��6�Q��sdW���u��TsK1�T,�&��*����e�C��8�s��0BU�;���OB.��-?������͊�Y����<�0_+v#C���t����0�g:�m���ڜqi��p���v+���R���\�t4����Ř�r�C>����驃h���~b-��8@����b��
�М�(�T�az���Z7GR�3��[���E�b�>���i���?�5=_T3x�uT��/kD�b������dܲ9s��r"�Q���?�����c��^�vќ L�`t����
��[���B`��F�w~��*��x0����XOdY�=H�U�>O$�O2��[��!7�_�ɺ�����YRƵ����@�w��oQ	/{����Y�"�m��cr�P�L�C��T#��+WwV3u�9�.C��Z���I����r�]Ҷs�)\��?D*�f5�����Z<
a���|+�")���;����l�VWǘ{'Ҿfa�<KV�ϓ��L��,?�KB�}�;"_*O�q/�`Gs�n��B�;VWƚ�"������p�#Z�T�F��������P����2��ﰜC����9ʚ�����f�Џa�E��+����K�݀���81��z�z�høN��j�ք��ԇ�e��g*����xB���8��^�n)��k2�ٍV>��M�!�o�CGD���N�%�%l���\*���=f��2'���7mݓ$�.R�q7�a�=l�?6�U �,�xu�~.���5ܪe{���S�m��s`�"r����O.ɩ�'&����e��gS�"!��K�����&��IVq��
��7s�If3s7[��tF*�KAaMT9�Q�,Q5�+XO�*|lG����^տy:J��y���C��MsA�����.ͨ�ޮ�N���%�Ƥ�a%fawJ�Ϊ4�<E�κ|�S����k�t��.�=����N�Փ��Y�7����(��EZ�N�9�zK�LۊW����BQ�H3�<@�F�~��`�O�o:��b�����V����O4H���m���Ղ�o�S���Z֣����CA9Dvv���V��r����*nn�24MN{w��#��S~�'H��7�ȝr�@<�KO*)'�P���w�'��P�ßF��~��d%���e����#��0j��ѣL��(O&��j�n����aK�I�)�De���M��VI�ڽa�3p��{Ӷ+Ɠ�9������{/����8N���b=~��!t ����h�� ihL�U��ac�Ŋb�	�����p�˒(�`\,�r�j��$�;X�/	�2�f/��苜[R�!~�ư�%�,�wb-�1�;��)��}��#�sS0�2��}o��e�%�Q�\f\�fy�]	;�B�����7I���W�>��3V����-(L�/��_�H�Y|ߤt�Wm�SD"}A� -��D>����G�e�ܭ�ͣ�"I��bļ�Ϩ N��iĲ�Kހ�P�\WfP���k��,ˤ@r����쀪�J��\W�d��p�y4uU�W�Ig䝡� z��rjZ �!�yu V�L����]wq��Ic�Դd����">�~
r�)�D2�J L"��S>�7�!��Z3ғ��ȿСk�ͺ��-j�2�ʹ���X�"�nq��*� �(Kuæ�q�`]8��W�]Zұ�%�U��Tj��Jj-/.ɋ�2
��w4�\;��݇��v���q��L^�@."A�����+����ҧ���,u�o�BGD��
�N�����S�>���u+�S�\=�Q��];�ؿ���	5,�v��S%�`$`J�I��H�$o �E\:t� ���9ŚC�?�xM��'����g@���x'�D��xtM }�?&Ӛ�����Y�<����� ���-�qW�+�cE6�MM�a�;���psb�~F�~ԈET��8v��S��+��p��x�)17����ζ2�l���=┡�_���85��7r�\����9&�/ƫrC�u���+	���W׺����CViLd.&SQq�>DWYд
1ػ�PNFڦƮ5��FDi��g��Qk��k�̖�C��m�-[aT�ĭ�+P�G-�o�[Ά�6)Մ�/��y�^)|�n-Q0{L_�F��P[�T���F$�{1���<�-���0��"��1=Ue�2M��t1ˆv�6��71�k����-�@EE��_��78ˊ}�03(�S����X�k�sf�@ǼݏPg�>{c�\;�PYR��׳a�>���w�rLĘJo:���o��[�A�#���1��n���A\�)��=��5�to���B����d���hά�$<ʘ�E~��=��ޣx��s�I�*4���t��7�=�yP�MP�8yM��73�Zm���/\�'n��4�̉��������}��t�,j�r\sH��Fvp���Q�kW|+L$Ŕ�b�
(�m�[�%���h���JxA}C���¡'���y\�2'��A�J���QV�Z˂U��0ɇP�y[���h媯d�̹��9�Xa�Fy��^3���;�@��|�`��kG���V�AB(Zn����t c��ny�jz�s�Ԝ�#��7R���۳�Q��_|�x2G����9�4��L7f5���N�5�p�$�.q\"]�8�KL�o�����q��V����a���d������bz�Yʓ(_1����k����-�"���)�Ҫ_���mӥ����&ғ}�]Ζ�eV��xm6�3�9��b��nYW�D�(�nC��_M��X:�Bˁ�ғt���}Է���9�'r��^��^���m�d׉�.���$&a�;&xDQ�=��
��|����n⾹��2�P��Ҁ�%l.gs{�-���6�)��t4�P��VX�q�Ξ}��NHD�X�QR���oG��(;X8�.��VN�{D ��zY���3|���Lm
�gp`�e��l��|���h3>wǒK]7�3��0�	����ˆ���,��s�B'mWP���K�.�;%�[V|$HL>ݺ�h���NY9����]�i�'3<V D��3�y��#nw:>�6�@UEOU����*
�8ߛ��s�^��i�Rl�>h%��Lχ����L0���}�6e'U�TBX�v�6�6��ChBf�!a�W/���_�'��E	���CҰ��k_��$�/����F+��7Cs�Qρ^6���&�u���5'CW�A���xB���)ܚ�<�c0$�Đqa;$���g^�4ű0�����G�MzT�^��8�4��Ko����*'})�%����Cv ���e�/TfX8N`7�Ύq�9ܴX�Im��`�Nh	�y�On]�嵚|�`xKg
fzo�6.o�q���� ���I���B���AU�R�H�$�ח��?�w[P*�s�&�Uuw���CH�`B�<�
������n����
3�)��8�t�b�vW���p4�? � Y<�"�8��Ď���a�±�~�#7�އsZ֎�#�d�ӂ�`aj���/`s��{�G�$�D��޸�~�ǩ����� �y��GS7Fs�`S5PV�(�eRR;�΅�Y��z�Hq�;�`��rgBr�\���\���{�����*���J�`�ɵ�mc��l]�(���=��=��Unˎ���{��A�v�XtA:������a�����⹟��< �L͊H����F�+��hO����h��5�vK�OwtP�pm���]��3�w��e��'�%�*dy-^sAI����]�L��D�8+%O&��D'��5���:,HO뒖Y���L�7q�o!'%�Ѻ1l������E������j���!h�_n�W�3�	x�����vR9c��������@;�^&�~���?�7�8�s�qb���m��7&
|�����[s�l/ç��Wl��qPi�%�:����M�ݠL�C��*��nc:�c*�	IVx�^�� �f����2�[��)�ıe*
l����̯7A��9���l��D���0?�>��h�P#'jVkǞ�������V;��Z�h�0��#ɲ��y��P}	JU=,{��&� n�
 �'@jO�**᜼gi�"�Lh����`
�9}h��9=|J͂��8��3���iiD���8������i�Ӫ�U�yhYb\���Qe&9�lɬt��"��h}��X�'�c������j�����w�Q��fA:)��O?c�$�bB!o�����O(�6km�s���;�$�=����X��ེ�uv�R��D(i's�$��>~�I�͚�,Ĝ��:��"e>#����הsN���C�j����Ϝjϲ�Is̘�hOԊB�bN88j/)�-eI!o��ƹ�v�+GLY/ڽtB���� ��W�XB���pN6Ga^������cW�m��28C���F��@���?V1b�i*������K"1�"hg��Se���P����۝���#�0c�$�rZ�5���	�5�)���ě��*o��sn6��0��I�6�Ɏ�;��r�Y���"`�zx�F�T���~�$%��{��\�=^��4�%X�Zd�ɺ�5��mt�䶚�H��E��)��o�*�Kv��ZZH��JR���G�L{BI����>r�C��|�X�i�s�y�֎}r�����j�
h�LNJ���F��\>�~�ܥS��Bp���8^�ҥ�&Vl��9�6<
Q�(=_:����2�Cm�s��������)�]`-Lm����۞�J�Z��ڭB�V*����dz��:��Zb�B�O�H$/��u��!ɌSH`3�R�o�?�N�2s�b}�LlFݒ� <� \�����C�����m�y�!pfK��*�!U�)�pv��3������8?�>Ce"�1S��|�,Zd;"���!~t��O�Ee��9�Ϡ�w�XI�ov�O<�3�Ly(}8|"p���_��&j{��i�Q�����d����*I�2O�~rx��B\�����,u���F�$nk�e�� D�2ƿ�r _q���~̹⚌�A�r��
�RP�%Nj}�����E%5G�Y���'��+ݿ�&�K��}���F��T���b��4B̣|�F�}go*�Yt� �c��[��H�G$�0Šؗ+�,�_pm�*��wFQV_62 �Or�H�z�����_�ex�<;���b�9\�Q�5-�ʿf�<k�������m�c�s���6(���2��ދ5#��D$�8��׿K8?�c~�5�*�x^�"m `��4����hqz�AAo@��*;�~p�)�S(
f;���T�Aq#�p����)��k��s1��Ud�JΕ]���5�,��W�d�<��[5��A g���<�����Njճ۽�-U�=���Aa���j���y�H����n�B��3cY����9�~�����]�Y��ѣ�����b�T?�H�HΒ!���\���xb����h��s�dS�J��}VM�l�Z�ԇ��S��'̻b��
�Y�;���%�����7X
��w��O_J�ɞ
��S�-&!�ׅĲ����zcc�>��� ���>V`W{��O+�E{D���g>}�;���r�
)E�B�Ǐ4��_
�.��`��#n��.���"��VAR}_����`*%:#��B��\�u�|EM{��Z�eH�N�!�Z��;b@|�i�e��	]�F��i��=���Ǵ�+iH�1%xr��w&����F�I���JU���1��0���P�L!�6*9�����e�u��
�]?(����	̟L��H�+�D��v�p�b�#\��#Ƹ Ud�X��{Tڕ��V3�%g<~�d΀kx��'�L�jr���*�2@2�����������P�.Gb����hP�f�\(�X�
��Pǲ6=� �����x��ӻe1 %�ي-��9�ޟs"��`fOAAM�|P�!�
�"h�M�J"ʊ^�ɝx�#�Ǡ��\Y���v�tlR��� g���'�Zvʦr����=��f�����:�i+�q�̘�*�vYƈ�� xɲ�(e��o�tT��Aοq$9W��+?o3�?��Jv�Hcc���a�)C�S58��N���O����dg�#lkz�Ocƥ:��x_�0��eÕ"Zi97H)w0wDi,A<��E#�����._�mv�|��E:XE@��R[YI
�eL'���,f�cӇ��δV����*1m�� �ul���(T�7�H�$&ɇM��5��c �k��[�C��F��@V)M��֖Z�}('�'��r�X�v�a~���B�䣒F��ԬOƠ��2����W1�zv|#S[U��N�|m6�^�����
����(Vv�����u�A�;'�-�3�]0�_�Q>F�s�����2k��&�T�>�uK^3��G!Q��C�>
f�"�,���n!��!r�����n�Fs�8�!%_�g�i�u�d�Y�ߓ�ez�2��g��a��T���ue��b4[���H�L����A�:�@�o���Į��4��nua@�.(з���>����3��{t1,���g��h׳����v*_綪����U�Hg.׾�2����q����+�f�����|����.�~��;�N�=|K��+�O�ڭbQ�Ͻ��Lc�{)�3..�`X�x��h{�ݚ��Hf��Q�т��ְ�F
�*+�����*��Q�q�y.�5muQ�{���`�U  ]��0��+�a�Ai��-rT�&��:���zW�]z����*��#��uA<��e����5չmV���3!�;#U���s�/o�w�E���F�@���ᒟ��m(1@,��������5��$k�y��
8-!��i' D/����q��9�;�Iw�@Y���~?Љ
���
.�??�r^�\����9`3`]�m�����34=Z�6��ܾ7��O]��;�?@��(5;��GeY�N�8/��9���ǌ��ȇ�s�lr|�<=�U�ia��8?�8�cI?.���X]I6t�4�^SK(2��= �\</&a�-`S����:
gu�ƀ�H�=@��6�M�����Tܭ��ٸ0R�B�n�3�M��3��m�b���Ad����
��@t�?q�G�*~�=ʶ�v��;����m UY���ځ&�M!}I��wn�ݗ?r�*J�.��_�^��[/7��:P"���P�ǧ
�&f� ,�Cz����ch�����ކ'7>O1� �6x<�Xw���4�j�Ʋ�NEsq
<�/%�B��p�-w2��/E�+d���m����B�psP�8آ4"�z��P�c&Tř	��/�BYk�č�UJ���g��tDy�x�v!c����=�K.זB��ّ�����O.(]��^
��7���o�QT^����I�� d|<tD�J%