��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]����j6�Jr��*}����^��f�,u���0��������#�ޮǘVtA�=�X���F�a1g�p7��0=��Xe.%��y"Hpas�����,���൷I_�U�SI��ZK�&���\P�4�&�=h�3���am8�F[sb��v�{q|�W�r�L�3�S"̪�*��7B�K�"��sS��i���{�rg�.�v6X�矲�J�C����%^c��͡�q��|��3�ED������Gg����7
�M���C���|��e���!�h��s�_c��"�����xp�U���.V$̽�_[�_ݪ�(���t�Pe�F���3�T����ۨ�
��G�=�[�G����z��4)�L����H�}������:���Z��R
�-baE�O��V'�� �zN�t0����-���Ȋ����U�&��9�������H�����,v�RK���P�.h���9�A��;*�]��9����2�4O{�㒞�a�=��x��">E�\����!��cpP-Ձ��@�.C���$�ӯ<�x:d4�ƱY#�S P�?�Z�#��+T27L�rq�K��{����G~���0� T�V�2�=Ƌ��G�>5���*�{z��!g��}537z�	�^��B��O+��K'��t����o��Ĥ��6��.�[�����aC���G���c����g�4���$�<�ڢoH�:0s�'^cY�t8:U|���'��W	:��8^*�e>+;�7�W�`��H2"�>�y�a�jN_\�]y1]��=`���O�@�S�aª��b�V��˂ ��U���G���}C��h�s_����"4�m�~�,�am�������!_��♷����^BW�����RBM�{��&b��`���/�t��B�w,�W-A��c���tim��$'���K���
	�o ����ӑկ^+hU�
�&I�Ww}�k�E3��}�*��>�d�t7�F)Ԉ�v�Б*g�C�HY�B������Y�#�B9x"�=��9Q[���_�B?i�E��Q��D��6&��ГX�/6��pm}I��\C�Z�B�Ր6B4�7m=Y��3�����
N����zj(�{�S�%,�x标��/����Q����
��{�a���<L�4����J�F�
��R8N�B�2�%1qɄ���X�c��ң9M�f�����#0� :5��4�Fc=Dr.��
�ʇ�A�UB�@#m�-��x:z���Ȣ�<�1
)��{/4��1-p�m�s&�h'F������'M׊�I�pT���BT\�g��dJ.��վ�W����_�����m�%#��h���umM�s��5>�I�@��|�(�K[DQ��������ڍ������c����8[j5	�	��Z%����΍�ţ�#�cpL��c����*v�I����F��ݛ�*�2��8�
m�$�[�Lud�EA+E�e��|���[��l��.��S�yGU.�N��5dD���<A��,V�|ܽ�,���7fat�8�!����#ω����<M��
� ��}V��&ds3q��A�`Ļ����)q��tD:�я|��T�0��QO��&�� Dܵ�UU��Ͳ�/�A�2u&�^�ŏ���U���פ�y���qxH���
du����"0��x,_�M+�
8��ת��[���� H@��� ���L|�7o�B�\_T�K,�A���c�_QZ�g��
�w��SjeQ�S�Dg~��hL� ����'��.x�7�'����$Km�Bb(X�4Ę#�~'߳"�Z���@�Pz���η>*�!�lx��@�}U�}�:z�;���tZK��4e�{_ס�3�V4�-G�;�:�<�) n@��3�=��s��3�FG��P����g��m;��#lDv���bW����Q�5+�(?�9ZV�ةs�(�sǤ�� qEl��8\b����.VGx�P]��N�hf�J�1��������/�����;�b�X7�6qh>��V�3-E��.��60�g_>�'�H�;o24������3�*��|J�Y�>zw�?�8=�k�cfW6V�G��U�}n ��Vŋ�N���X���{l!�3�*w�MS�_�M���2�D�V�2�e
�i҇�r����wH GG6���n>ߘe�,���L�O�#�����*� �XfD6*��@g?��^W]��3� Oِ[����㌑�+� ��d�
�JcLE1f�Uǵ�{b��}/Q�Q�/�;ͽ��U�e�3J�����QK[H|�4^��z"B��øŋ=�/߯;��qs�d����Y=��l�:GP��Ai�EI2�YMB�����O]���J ��Ń��t��m�R�Fc-:+&� WT�#����F�lֱ32�ᅦ�'Y��[%�ZF�B<����E'�*�7U_r6�?�����j,�Y/�⢩�L�כ�1�\��� k�5�9͓��-�R����Rċ��S]�����6�=}ؒM�>�D�C~�o;)�����%ow'���?�f�+�	nMu�(�K�"�׌�u��J������Κ�x���\y�d�?h���~���^�B� ��;f�e�}�����D(�aC�J�'�jɌ��K���B"�P���M?��{�Ә$���%s���SK93K+B�&&s����;���/o�E�DF�ga3�%�:�����|��̦
RG�;���I��W����f+���}����|��W�nq�]Z�w�n8�a*�B��(�:g����>�{�a{�~���հع�7�`����}�}(�FY�r g�Z��~A��K:$��?�˘�-.�����$�\���A��Hw] �5�z�(��<|�7M�f*96���Q���ϥ�������?{������^�[-�fei�<�`��!4X�ne��κ�U�n�BZ�l���}�д�$���dZX�z�p�}��[�H�An�g�[M�y7`�L,�hn���^�C��� �XUqȽ	.K��ȶ�Q��D?D��\T� ʷ9	il1�4@�g�In�W���,��m�꤉vW6��n�H- ����\4]��>�b��8#f[o����lϗ	伻�QX.�Nxd����c��w�� ��g��׈#�1~I_-��r+�u�:�LW0��酯��l�JH����)2�]�{��ڄ�A)��ޢE ��0��3��kV�x�@���8 5�j�aƄ�S��(;ja$Ք����[��Ԙ��(C���?��T�t3s�:����$X��J��K���͐E}l�{h#M-�o,�!��
P��RQ�,��[�l�Mlb���}%�8���́���qf�lF �k^�-��/���y�O��0]���U�)��/o+��:�y�����"Ǿ������j��v�=!��P�! ��O.�7�1�����[DA��3�f��8�l֝����jwn%f�/2����r�8�K^K��'Y�GS�8 �8Ad�z�P�����`	����Ԡ��t�� f<��RO���^�� �x��l�M�M�A��B;ik��}�3yQ�>B��2��D��>�i(D�M���+��_�u%��j�ݙf�����]���$�v�/��K_�1'�嗅r�?G�}��WwߏN�����I݅��4�4B�*-�r�q��K`�"��\�m��e���>J6P�r��m�$M��x6��A"��YU�K�,ɞ���A G5�/�x��|�e��Ho{ČDݑ�Xeo����"�$Y Y
8Rr��Ƈ��i^�B�K�"�
2-E$�-^���b��toT���.�gx�&��+P \����
�����I2����ㄸO�;6P�$O#��}���Bm ס�Oƽ�oM�Ux�~����}��n��P�]���4Oh�h��1��x�J[�q����kD]���E�E�w��a��L vډNȒ���f0�d�R��Iq�����T�^�єDg���VD/Y�adT�ԏD�@�KS}���X�~�����s����6Y��U�=����ZT���4ᒼ8&�VE�a]�j���%�e�zv�eh}��L��~˯��{%%~6e�|��ْ6��w����70��!�����r�x�o��,f�|7js�[����g�25���3n����r�]���5�D���@<�׀V�3�;�Ι�=�RV8]�k�;�;P����TP���H�������=�٪��Eaj��8wd��go�y��VV���J:���u��t��Y��9z#�˖YJ��I��'RP�8"#�l�b�^��@�<+��9�up����p����
�Sˎٓ���JǺ���ޗɦ��ON��a��:�z�����摰*�7*��t��J>�8a�r8�A��S�^��?*�X��p�B[��<���!�o�*;���Q��a[��0��}�CamX�M�����F��u`6 ��aL���m�����Y���g��,�c_S�k� ߨ�`���#e0�.<��	�[��=:3�ߡj-n�9 �k"cv������!��,,(�5U3���1��#	�k�>B*����:%r�%��6�&`�Sg#y(�L����Σ����yD샺�G��o�2��h��}̜;��٫���w3"*�f�&X���@�Ϝ�.+xd\�&~���>:���9��kn|����ZP�+�9u�~��v�('$ �P��eQ7��YѲٵ��{m>�:qt��<�N��0����w���E�9���$ `yBܑAߛ�
oV
��{�F�ah����XQ���oN���x|�X
I���("�!����I=���<�u�L��������u'�^|��+)mo��`k���=����D6�J�H��Up��~�/Kr����I4m�8�ֹ��B�3[��J+O�ˈ��B=t�yz
���wn������L|Q)�7���)�>�_2�Y�r����iЫ��&?�~=Nov4�b�`h��P�5K�=�X f|<\���)�z��B:�d�Qߠ���|����%��Mc
�K�|VE�"�K�(J���8��v;?_���m��{&����ײ z�������ʛ��B(�,��ѧ!�p5��a���\o� VB{�-�L ���ue>Ul'�������l���h���݅p�~|7�pM{�S��'A:,R���;�����+�4q�ٮ��2?��'�-��ϯ�$"�)���]ۈl��;�#���c5$�O�M�;�u��/���g�S��g~�~�󫖛,I��F �.2.��V[Rrqz"��[��dY,�<T�����N��XR�/��Y�2��f��v�o��>�|�ͤ�<�S�@ܚH�-�[�N��"��J�{%�3�%���:;��L�s�ԏř����L�vØS�O( jC~�@�����	���͛�;Ӑ7�7��M�30:��iiǲ�H�u]njX�9Ie#[l�ov�ms��m����x���ͱ2��6q��kb;g*��3���^�|��	'`���$�y�r���Z���>5����I.'���1=KZ�KRMt���7Ի�"�__����d���.�U�.�Q�,ڇ����!�s�o�aC�R�Uµ4^,ZA�������L!-�K�ފޖ�)��tqO�m��m��N��5���s��|�/�x���E�$� �sj�����;(�Hp���Yl��0���)7��j�;C�հ��v*�c,��Q��<ߙkhei�AJ���I)���Hmd�����D}�u������כ�5.�����ގSX�g	ׅ��b���a��W�sZ���K՝7�g.�Ù�p܀1�f/[�^�"��[�,��}�f'�p����ɳ->k�q~�������|E ��kc"c�N<1��P.ٕXㄠ�V�-��Ҟ��oҢXm,��Uʷ���lG�e��X��T~�Dq�+�iI��	q_msH#H���v�:��#�y���+/01�<P�B ;�(�e��Y����`cR��AxCT���JJ��Ux�	���l��7l��#��[TFh�W�y�߁�2�k5�ό3�pCz���jx�NA³�A$�X��w����o�}��#]�P��pݯ�z�	t��2B�bX�ng�e1���v�c̔E�����W6�-$�dѾ~�,J��/љ� �wQ��W�$��ꨟ�b�7�#��H\G�����Q�"��])�RX/ E�PP\��	6���d�!gz�U8bEyP�_�������e8�����x�>, �r6�0"�;���zo���ܜ^�7xMә;���ȯ!�p׌��t
2{#�[�B���,藈���KsO�Kx�+f��k��q�N+�H�x)R���'p��4��`6"tө��)�땂��y�M�[	��҄}M��{{3ĝC�S�6�]��nmKHPZS_S¤W�S�D��g}	Z;��S�z�-~�V�|���?#��>��V�K)���ׅ����W9ҭ����k~y�,S!*l�� ��4W����8�^�7;��0]~���
�H�9}��C���ΰ�m8�@A�$��$���ve0�Z2̛)(G�5����)}!a7X�靈�����y�B��y���01��Y2P�ސaRB����~��"���z4��A�3i[<};��B�q%��~y3�$�I���#�G��@�+�=���E訿1�U v�D[��>���ߍ��T^�(�j$�g�I(O��=��3��!/��0�s�[�M���LHVt;�F�|�V!8�Z�#i�7�ޕ )M��/����~Vm�֫)jr�ߋ\g%/�N;�N?Ug']&KP��f7��LL[��Y�n�,a�.�y4>��]NJHW^��D����l4���n��1+�?$2V���V-�"��U�����:���)N�q�~���������}�V������V�2��tzj�)bp��f-����o�K�SG��P&ǳSU�j)��v�W�a��)�X�@�JEl_/9r�k[���u
�`75e(&���>k�&9_��Ј1J���0�헵�#������BӖƇrn⫠�=}� �������vNbZb�1��Z�ӭi�t��������j��GdFp��*-�yHk�K�?��?f��GQ,Hʼ���G��K�����ä2��R�b_���p�'�^~�k��1��S4�upܻ��C�b�)"��� q���Z낯�N��G�
��'K���,#�������iŤl���ڛ�60yK�����&����CGf%oM�!��3z�^b��K�cg|*���ߪ�>��C�a
�'V�m<Q��7�E��Kn\ w��C<vf>�[�xP�.�����_�����3rmD���O.��� jB��l��H/bY�����+|#�$�1z�r���Ns��!�{x'd���h�lt�9(솸3aݕ>�oGa��dEd�h����B�&8f�f}�E[��L$xS�-9���UF�^��Y[0ZZ
���=E�]��d��w�̳o�ب���JS^�b�U6��W����؝�s�6/lg��ɔ�=N���d��3��(	�r�;�y���Jx�_��q���ht�!wC�K�n�緑'o���7i���7�I�wk���@z��K�Vg��dt	�?}c�l��kki�I{�\����z�h&��	��@�7�k���'�( �s�<�Teˇ�;p;�͡+X�2�K�2������� �1Bz�C�X�]��ξQ~~�˷�WO�Bwbܺ�ʵ�{qU�����}���� ˈVb���^3��"�?+�i>�g/l��ĝ�W�*aR��M����.�#�Hgn�j�����%�������ʨOɧ!��Հ��삌u8f@�j/��8{�xs�F^���)|ڹ��F��n�vS���zs  �x���4��#>;��!O7�s]�h�9�f��J���6�a5�A�.Ut��"WT�?M�9����\U���=���K>"�}�|��NK���
�B�͒�����m4Еr�_U�|=ժl���ϭ}���9�����ܞD:;A���'hTcH��U��fa����m�s Xs]��@���՗�i���#&ח�7�ی�ZN:�� q%ߑ�~�^9˫��{�� ��$�W����`q���Z�*p�z�~0:��͔Do̪qW�*��>R�rX֧���)��UM����`�Ho�:��G��V��jfi�b%4�����?�x�	��l���������5���y���7Y�~�(��f��|_k�OZ)���>?]$����H�㙯y/��Z��F���Ǒ�����I4�G��4�C�z�#@8�[�^A�~�67�����"l��M|�����#Hy
T�☴�8c�$V�^\���բ
o��%Lo0@��+��K��A��4����m��&[�՛$�"�ٽx��Fƥ�zG!l0��齃9q��Yՙ����V�}�JR+�:Zh��~� t��8�47�����u�Zq�r>J�nU]��7�c.p��`���t�.�ɛd�il�a���[H����2l��
��L墶���s�>��vǇ;I�h�N�;s��ϡ6�����'�t*~��p�%����1G��9{����5�*�����N'�vw����� t���և�ꐴ��د��X�]y��ѻ ���];�?��zay����Tm�*��=_�V�/��@&`A��\6#Cf�����<������;<�A%m������<Mh1Y|�wE��6��� �R�� P�IpQt��{���0z��ҔK���=?70y��������qo�ٽGeC�0=2���M��@۹������(<NPȩ�h8�`��=�d���,��A6G��9pL�y��y����O�m�S������BH�96���G�,�� �,�'�,A�1G��m@��D��=pe)�^$�h2����s�ѧ�2�a$y��+��d�!�Q��V�7{!�M�uF%��T�A|.�L��K��#1��6��I��{�����