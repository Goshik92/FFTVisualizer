��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|��&���i} Ĳ?��O?!��$v�X*�y)�ޔ�$�m���o~kG{��cn�B2��d�f_~:���f&n�d"j�i�5�Ų�x�����U��*��]a��
5i�&����Ջ`�ɿ�0�0H��9���D�P04��M��b�/hrxD��%�:��xd���2<�V���l�M�r����"l�~�nT��a�~H�(��r��U)�v��j��:�ǵ��_�u��z'���"���Ѽ�����.w�����N�i���߯!6G��e5��B�Pj�2���3J f9ݪB������/ĩZ@�ؘ�b��Z,���L������Kti?GT��Ϳx�.�M�M?���d^Ӎۭ��r����$� m&I2��=	�,z\y��G#�M����4�;�N��{��k��h��N�����9���B���o<�!�xN'�(W��m���a�NZ���f)	'�Hv�@;�Kw�WW9*Ug~�ɄW0+�-�����\�և�I��M�@EܷW���w@�H���V���˖;/Y���z�f�H����鉒}�]���λ_c������ru��Tw�����d���d�`s�YM�����v�D�J�
��tf3�[sk� ���߳��e)2���(��os�تm�<)�YV{��m�L�O�����k�y_�9�0�X�v%y��ՠ �(�ޢ�C����Hu���'�rܾ������<�ä����ц�m�S)z^�Tf~�oeu��Kw�#DKWy�+R�W*J�@�9"2c��"57�5�YLó�c(^��Uup�Bꉫ���<���S�뤸C���0�j�
F�����̈�
��H"(��D�8�ƾ�H0�/���n�G�s�Qە�L��#��c�.^ЯٷXwb/0ͬA,uh��a���2���v7����p2�LM���Gb �"-���M-98w�~<̩x,�L��*t|f��4�%��4s�B���J�KC>aHlf�.?�5�rc�����$�?������Ы?M^��
Xc�3b+C��k>�P�8����7a����B�I�G'�[��\���䳆.u7� hW��������Ѽ���d�lM�8R�f.����@F&��k��s5.T�X C
�Rh-o�ȡ��p�DK��F�%r}�ѳN�a�ˢl�YN�c�X��C�&�T��R(yY�mѥnƈ��h!b����6�/�3ҀQ&�0�#�� �P��{��z�o� ���Aԍ<oQ��/�1�����P0��G�x�N9ʠ2E�O;¹ ��\J&���mɈf'�T@ӈ��,Hba�3�7�t�Vo���4L�q�xcOJy�jH ��q>�� [Z(L7�d��ӊ���`\���vo��Ś�@C��J�`H&�s�a�U��vt'vD�4�֞{�(�~�<�0FY�w�`�q~7�R��IO-���7�
N�B0�v����3j9�(*B��[wg��En�!8��2>�獷��*
�@��>Q9V�VQV}��ֵ<~�o�f�aL`����U:����EI}@��h�(���g��UV�%�0��l�G���d���~�%�@,PvHq��鞄�=_'I��,�'oU#��y'-���-�gh����� ���3t��,٭�Ԡ�
� <^%���Gߛ��>�rgx~T�?4��ԧ�o���ƓIQ=�͙d���K�yF))�-�퓥z�� �X��.���Z�wۨniv�H�
7��;���6��\J5+���I��!����;dM��[��ԑOS���9ѽ�>j�έ^�K��Nh�+ʙ3@$r!r�JԳe�:��6�Ю��kk(�L=�y�l�!'q�v�E�yeS����j��Տv3���|\Zy�0Ka�*����"��GP�ڍp�t4>�ѽ�4Z'/����
f��W�ZZ?˒I��z0��S2~�B�ݽ�� ���B�^� G�$�Q�>���nD��e=#`�!NJ�@�\��e�6l�7��U.�bx�A�?
���v"�C�ʁ��=��;`���C���$y�{;�68�m�F��
&�ݨ��4���Jz�9Tp����/�xLEƱ�}�ƒ�;�P�rأϵ�?b����o�m����o�Qҭ�o#B�z�mm�V�����Z�-0}�֒�s;,u�$��BX��bؕ���X�h��6��e��Q%�l�=�Zyz7���3	�Y�'���E�� }y�'��T�%�q�z�=�Է���@����������І%n�sЋEE���D�m/�x�)�ʵj���0v�����)E�@^Е�]��/�}�2~$�g�x���b%7��(5'��b�;I(I�'A��Y�g��r�̤��p�y���6Ĵ�ǩ��$T��
nZ�P���ܳ�2qK��}y�.TB�ʾ��{მU(u�	!�����>�
o�k�_В���.�KZ`�m4j�scX��d�ks�w4$o"��q]����wN3A,']-*Vr�� ���k�%�'��/����qPLmnR��His�q���{�0�}?W���i�-���l�K~\5��p�I氝韎�&a��A�WM+׹���j�a��ך�b�BbPZQ�C�l�p|���ս��Gh@5��3�uF"y>�ܗ{ρg�n�=@{ʳt�b�l����~μ��v«m��=F�]�2�F��.�Є7���?���m�,���_H?=��Q��ď�'	G�W�crg䨱�<��S���mW#��?�����?���;^*-���6��	k�B���q�8��O�J�t�T����~j�z�-�ڄ��t�{A�:����·'�N'��q�`��L)wD�r�.��s\8�J����$A���P_���*V`rtDs�`ro?�����3x� >�&�y�7պ�"
,qG�r�6���`<�;���t+���&�7$���5�|���u�ꛘ]�@s�[t��Gai����ѭT�6O�K����9���d��S��� ����ǋ�h�r��Z.Y��n������NT`���|�~�Fw=V�#��~BSʭ���am�<&�6k��N����#��!�E�8R�����9Eѧ\"␟b���>�� ��622w��=�@
6TF�����3��$$$�E��TC�hfG�"1N���9FeYO���C�	 �[�B D4_v}#ב5���y�y���Ǡ�C��O���qZpԸ#>~�Tq��˞����^A��ܥ���U֭Ntݡ_g��_9����&���{���+U2f����,��SB�SƯ�P�6]F("<�E25Egԫ�_�wq);�S�u�۷�A��N�����M�r�<�4lC�|	5�7�Xz���o�Z�f��[�Ne*��տ�cyR**�x��I �V�f���W��>�f��?�F)#�Q�}�5M���G����+C<FIZ���2��GfŽj8��R5Ue�����Ū�������U�Z�:yA%jP�8�T�#��}x�v�}PyQyL�ߴO�"U1���+~�	������K��e�z�~�2���I͐���i.�/N/�L;������"Z��I��T���_�V��V2瀘�|��@W�*�u�����Y�_g$�Ҍ�0�L+ۯa2�-��==��!K�܇�t�5dJ<t�q�J��QV	�'�3������<�(��ˆ0gܸ���,��잊�wKbd�S�eVd��%�c���-��M��?^��F�T����;���N��9f���d�qF�yz?�ě$w�7B�:b"RN��⡭���Mт����H
7�Vy�������K�.�����P̤��4%c��i��T�2m�8�R��5��ABM�|�E���7�2ʜ3{;7�si�21`He���`��:|��	/�c˦\z}J�	�.��ah��P����6��[�w(G���mX4ݼI*2{ۿ�pdP�ϬV�\��x�H;�N�"J��%ae�U�%�C�®7����F0yp1�+$0f�� ��jp8h��h��b����v�Kb�9:3��&���#��ݎ�1n��g�5|��63�V
���������GӖRiC�v�J��ط��E�W���\x��RG=��ߊ�+l�\h���ڷ]G�����*l�/ޓ�C߉��t��YX��S��Ul7G��>�;kكqD�D{r��H��B�m��*��t+��=��;�C�_�*�BWV����@���@��ԐܿO�sJ*��Ty�yϑ N�}��S��@�I)'�?��Zf+�|�3� ^\l6�ԟ�Ӳ�[���
;G�H[���
sE `	��f{�l���\�w����c����<�Y
��Z4<e� �d6��4���3·\�M�%�\�^@�ʵUWW�pc<��7�z B^?;�s 8*�F�Pm�vI���(;����֌�G��t��c�P�^!��^9`U+^M :��ax�?k��%;_�̠�%�没^y��S��=��1͛4��c�U=Uf+/�z�Y���d����5vk�iwe]�l{Xɛ31l�p#�^ha����];yݟ��a!u��>+�2�J)6��yŗc�<
�� ^�K�X����QUe�B��0a���n�c�eVZk`#��hӱ��쎌�@�b�zSǭ}�w_�E�Z޽��c��JQ|�
Z�I��ię9���^�"8[!�`LH��J~�Y���T�7�J�#Y�"#�i�e)����B�W 
8�*� .J�U�y͹DA�a�I�'�= 1 mr;Zu��~Ě�s!���ψ���	�p9��bn|���]CyqX�ث����Z���ȣ{��Ah-�Fq
X��#6�hNݖ��W-��}�R��zܥk�	���qk<����M��qa.Pd5V�S�{�A���/���6q��u�4w�֯��jJ��;Q:�9a�-@�5�=;�sج%y�UZ��f/v{}8[T�Q?��yn̘�;w]>d���X�_r}�B�Ωѱ���{�Ky��E��6���r��%!C�'	�H,��3ՁͲ�0 �eN�E�f\�� �<�b���w�=��lDЫ H�WH!E�t�c�i��j�d	��	�=D�}�\t���l�
��UX���	R����]PMw[���?d@*��H��k�i��3�;���c�A��b6�m�;tV������C`J%3֝�#����s��zC4蠗]��a���B�Iq�f�	"º{��x�UYa�#��}��C��f���ɦ��ZV��C�����. 钥���&d��cs�e �3e�.��v�4M,�$�%{����D�N�M<�Aw����u��G��	S�=׍�H�I��Փ5����%z�: j��ޖ��Ϲ6E7�A�ᬣC�r��	�v��-y��~��:O���j�J���K1��PYe��;�LB�A&S�ߏ�<f�E���ܫ��m!�9�S��%/~;7`9�(+��|~�Gyl�t���7v~>z����[�8s��q�X�@���|ĕ`�h�Ð���ѐ��[�T�2R3����i �<"xI��\�MR8cES��}�1h:]m�W��Y��k]#Ԡ��W˷y�'��N��k4�fqD�V)�iC52���͠����@��x��6'����Q���<qӭ��'[9*�~�Ѣk6�<�S�g=d��͵�f�`�~\y� ���e|�s�u '[�Ȁ�C��emE�a�a����B�����}��g���c���RBz�ɠ�j�1u��v����*\����2�`��j�YW���L�%�9ដ���7j�����Y����"��j�P�Sh?��	q*LE�
lH1R����ը��#nq$��D%�5�}�w/��[_.c��Z��rX��T�ї����(	����PZ��X0*ULo.���,�Vi��,Y�����f:=>��AUO��1�TkM��*r�Ǝ@�8/w޴,��Z�g,[��yTmd(hC�G1�O(/c.f�PB	T���ݪ�����gsVĿv	֥�(o9V��¥�mu�ꠒIS����	���U��	��k ��ᒢ��^�o4U,��Y$�-�9�JN+z��1G�A5��.�*�0���)"�=$���m̓��0���.���ŕBuɊ�Y
@�L)&ޢ6���*l�ҩ�����,W��[ka�I��#VÂ�e�+l�:�N]�����C���5��R�zU�V�s��Bf~@Uk�ޥ�Cr�J�qD ����ea�����4�B��s�l����1IԈTD��g4ErDC�dRB��uN�v�� ��/]}?��r�ʜ/K��T���4v��c�Y:?-A�!��u�WG�~c���c�z]蟕��0��M<�l�(R�jG�gO�v��_!�|� ���8,�X��bXdSdX�#�]Ӈ���E�8c��~�����2�o��Sr�ܪ� ]v�V�y�!ͩvK�,'�LSJ������:��jA��:��hi�ħ�[���[F��0��6|�/���D��)�o��O�I����[�>ᢕ�z��LV5d�oh��_�!�8�������Iyzn������	��x��_M�Q���n6T$:�-����~��Z�R���g*�߬c���`6D=O��ĀW	g��*��~b�+�B9��L�)S���&NN�/Q�	~A��)f%;�kq4w��<��¯"��_ )��������A��X�%0���ég�J���$�����N�ER�����A��w�fX������6�(%	����_E�����g[(5<��&�%�flM����F�`hW'�"x;b�����Ѣ��*��y�b`�9v�����8E����?[-��&nf�~�G&_[�>�,Ӝ;>�F":���S���ojخ�X?[ʩ#�yt�^�.י�D|{o������J��.�
�y Q1�&^��G6�}���'cob
�b�T�R�ez)6�[�h���ټ�H��Eee�����|X�m������K�%��7�K�Q�����
�U��R�4�@}<
��Cm-0�݄#S%��Z�!�yz��u�;��p-�H��h�%5־M)	�Ů56�����m�b�Ը�J��>��	��.q,�{���*Xi�y����k��İ��XB�F�R�)4����}snr"�ëg~�i7*���P�C��	���(�ثP%܂s��0eCXf(��j$�aBd�H�7��W��I��=E�m2?I����_��gSBι�����&���)yߡ�����kS<�d�Q���6(��ӖM��|f|�m6z��f��EԢ��=��r�U�u����z��B"��0MB������ۆh���,j#�p�ϰ,�Y�#�m�N�}(���6~w�`(Iq]��V1�0 nSn��M�G���l
i=C822 @,��O�_������=� Y�ш~��'Z��3_fg���j�dX���6� �Gg_���7����B������M���,��O�'�W
����o�/�ִR����*�m��o��ߚ���SJ�F�v�p��"�s yT�2#7�^.�%��x%&c�D`�0D���:{أk�!��QUh��d��җ=Ȝ���uPL��g3(��
�OF�%�|9��iW��>Z�GB����u���Sƌ���n-�1Q�FŦ*����Z(�GOm�2��RM eyzU��\c�?�+���6�t���xQ�`��z�9�z�&��j�*�.�TD��<�Ƚ�¯��� �a�]��xb&1�S���0��z��#��lC��jz��5*ٯ1�h��������Ld�tMFaG��&$�j��l{���r�J���`f}�ikQUJ��h��\9{7��<)Ud!��m8���D��D�.N&�ංX����#so��T+��0B�Dtr̟թ�W�� !�4)(qPH��sN�"�n+#��J�[|�ܩ?�EX��Z,��i�*J_
�w�kE���l�>�^�9毧0�!���.���kr���ɾ���L� ��zs�dNg!}����,`$�S�q���%�2�X���X�.���?ԅh%`J6�,N��>�]��C�h~E�H$G<Ω=E��n]�>��7m�g�Iq*�q��ϣI�[ ����<�e=�}�����,yϔ���aS�,rʩ<iX �2(��}��T��7���q��~90�	r�ڡ�~��6�Ռ?�%�iL�_��%a�e�������V���4�,%��ݱ��>������R~\�؞�j�YX�2�����^���u[�r�0��}:scR�2c=vj��#�xv��J�zx^*s02���޺�^m����d��|	U�C&�V�ߘdo'�}{I�9���z�4%��~��h����l�~�T�|�>�MkH��NfY� �)Hoџ��ի��)h���������[�?*a�1SP>n2�!�Բ�_R���q[�s<)}����fj��o<؛�}6�h��;b����~�D����5������:Q�qwlyb�&�7�5���9�d�_�8���F������h�/Rv��9Q^����j�uX֦�,ܼ(���X{E��������&�r�ѭ�z���i�?.wq������V�H�-�J�>��k�D��̮n"L<M���{��<*
�G��5ю%�о CQZ��U�����g�xF��t��L��y��kY?��{��O�"�ECF�c�ھV�IR�:êq���J�n0��<L|g�Pc��?�c���
�r^�*&
���ة����xiK���8١8�1�3�}XE$�������b[���Q�;a�m�c4����������w4� �$�S�d�}>�{S)h��E�R�\#�籼cm����7J�%$PG6q��j��Fb��d�A>f!�/Q��w0Ą���ռ�ۂ���4��!$h�k����NӒ���oj���1��?�4`� ÷��~d�\�A��E��?)�X��t4���l,��X�4�"#%����1�x��\����#r��C��&���C�N��UZ:�_���+�h&���9�`�ȴ�����G����Bo��Z(3"q�]�xh��Kh$��;�%w�t��e�)Q�l'�@M�4Ϣc��,���r��nP#"��Al�t0�Ɯ׹��70�A_#a�N���#(�؇��۰A�����i�����D�=�Y��>c����ɮ͉�J,�T�,fэ�]Ő�={}WtV�.�ݍ1�}�������ptvZ�r��U5*$��ߣy%}C���#���j�q�z� cC�B�YepP� DF�S�g)l��}ݣxv�È�y�\ω�d���$��,�L�d�:��W�89A'-���\�t<������oK��㔶p��Hj�(�>��? �����71
�����ĉ���B�b7�ǳ`��t;�^t�WPI��8��Ǆ6��u+3�����41Ҩ���ӕP)mYh����ұ��m6e��/�1gt�J�1#k��^�*�E`X��(`�����X�~w�DO� ʅ'p#�����d��	�{���/�H��$��){?�A�=I#���lç��7�d��~@ �yP������?��FfO��ɐN��ٲ��G�c�8ܧ�r���EGUD:
��V��/�2��3��3��q�G,�����*i7 �lX��<⏶QK������nm��~��"||���_��v�RCwx��Vr8w垄G� ��~!�d�5�!�}�p�5n�T���e��b�Gd~�V������V#�����f���!8�ۄJ�۲��#�p���C�AD�9��-�I����[�-�ZRD��>.T�e%r�_�7I�5^�!(dv�C�+�9'�cX��琈 %2�O�͘#�VP�.1�C>ɮGL���n�q��*���ɭ:�m��vU��2��J��[�U�{-�N*�Xk1&`	Y��fcDq�����<��]����5�H��h�Qϛ N_��FwͦJ���~e�_�{���|�
�����C�?�z"�(U6}MM$���熖�qL��y/�>Q���:��r�Im���:FSHR�J�9ޅ��n�;LJ�Փ1S��Q�m�W7���P/~��(��X��E$�r� �������~^r�z���!�\��)���� ���F|�i�����G.z��r�W_j7|O5�B�<����Y��@�9�;G����h9�$D���9�����^?����.�Iʄ�A��q��PӐ�Hi=��j.���F���)���1��+�o�� v����`*%����r5�5�E�(������<��b�@�n��>-}�	{�aު��m&|JW-T퐧�&?e6���p��0N�ʶ2�f��M�ĺ�_HG�*5�${]ߙAa�!nR��Uq�A����u���F+1g�Li�K#�ӗ����A�l��Y`��f&\��̺���F��X=�D,^ۑOս�z@j�Z���>g؊���H�_p|�N(
����� ʁ�C
2�)>�O���~W�d�o{ar{�$=c4�9`&�x���A^dY�3��u����}y���<"��)���&4�i��7T��2�[��e�����gil�LVy]�5�>c�r�v "�R/�S�׌�B�O2�b�*>�ҖbW{X�dWThM��}�����|�7w���^$�!�W0��ߧ�{��I%����:�w�e_�$�s7Ji�d��bvmb��Eɱ���]	F4�N�(ז/���J��3��ה|}C~2�Q���TM* {�mX[�f��VեsL�#��<ϸ?�Ó���0`E,�Uy�~8̳��zIA�b�D�?qn7U��B{�Yy�(����w.f���#
�$�N�2�X#�A��3sJ檗p��3bҝ�ޞ1Z�B���<��G�u�)�m[�W������o��i��yMJo�K謒�.�A�5��a���]�286�Uv�sA+���H��?��w�Oކ��rm������լ`c| ����`��q��T��UOع��R}rn�^ZG�@�G�F|h/�}�9��a�cD߱Zr���� X�H��A$Hqf�o��O�ӕj��׺�R7�)��74��N�t�%�n]`�q���u�����x����[8\�)_���:ܳ!"R!����aP��<�{+��<R8�Z�+����!��!l�_���
�.����[��T���$�]�᣾���� uϕi�6[_7jKa�b{�y�C|̊�Mм�����jI���D�ؽ�_��3j�ܫH�::;��EV
-�t���>��)M7�Ι{R~J�o���%7l�_\a��7࠯�(\��꺠���Ԗ������ȕ�d�'[Xdd(��U�K5��3`�;nb�|���ȠvIwŝ�]��#g��4,R�����Ȟ-3�K\�w��I�-�J<��?ɑ� �K����g���T�>��_��#`��� �S�n�đ��Q��"�����Z�8��q��NԌ���T�DX ���1����4��{���U����d���!x�?�o�*,��k��7�(Y; r)��I�
8�7��?@�_�\�&�z��7�gBq:�/Dd�K睚�����eE�_lN��p�.0tU�r�lz�O��͇����E�f��{K�اu	3QCWB$�m�^��_{�+L�&5����t�|U�Gn�����y��K���0�Z�P����;�7=`JcQ�<�J���m����\qF踃�lB�U�2u�.�I}S�[V@�j&���4�F�&�}j/�/��/��xCA.�Fˊ�����5���"?#p�+ztkb���r各�18�EWꫠ���+ ""u2�)�6G����r��M�|H#���V�1��C���9^���o�(�"�}�̓ؠvU��}$��dk'��� f�r�m�>t-Έj���$�Gd�&���Z��@���FW|�tQ!ˀ�Ntr���/L�C�<{��.�)z?t��q���:�����C�!���)�7 �.�	
m��ك�98��sr���@:�7��-�������
e��ܩ�$ܔ�P�j�WWí$gH��Т�km��d�����b,��m�@���!�{w�q�zs���^C���CA�E��A)A�����9ڴ�b@�tJ��qK2}W�h�K�n�Z����{��|��SOǬ��2�m���?d��r��Rɵ�@~��;���B0���7q��]T�,LX�f
�|QK�Z俁�@ޣ�6훲�y���_��bZr��D��`\Cܳ���ھ}TŶO���=N��ߐ��W���qY��Mݕ��X׽E���8B��c���*m＝cr2U���㫶w���Ǻk�n���$��� �Y�����~_Xg%E�A�'���$65���!-�0�wY��������Z,���I�4��tܥfsN�ȯ�u7:`-��S�&�赮c�r����p��U�}������m�0	<��H��,D9��X"[ol>�r�J~��VT�3=,�(�~���%bSo�������bڼ�#�#.Rq���� D<n��\3�GUm	#O&����j�Y�a wM���b	z5��r�M�x�I�>�V�z�N�B�Z���|�.O�(�3k�C#�^.ړ�t]N��V�Me,ݪ��3N����n'R���Ȕ��| �-==�U���a*5���?���w�[L�Q������@��dp�Fz<Ly���NŚ޳�� Af�bl������D$=p�Y�MUp�h�3���	ޡ.��]��v�[�#�)�:�9(�(�[��v��9v�Q�{��;҉���_j�yVc�> 7/�����G������z�&a+�U�;�d�'b΅U�Q���ʺS�q7�q�г�~[tx���LD�(:��#���|��[Ã�o<õj�i�6Ǽ�]An�k_S�jN�F�?���+Vtp=} ���bX8f�:!>~&wQ�H	8�ɳq��ЎS�ꯋ��oU|�sF�~�G����[���V�1?k[[իC�qp{�`�<ii�N�����W	�6��P�'�����#uUi������H?��~���"��-R���B֌1f�x2�@}��7��ݵ<0Wv���T�H���Ib�S�fo,[�b*�Ø��J寰���z�2�Ǩ]���^M��H~ȮGy	1�z�G���4����NU�nr$_]�O6v;��7ʮT)`�D��o���b�NKUv�u2.�9k�f#���
��|���ʯ�������r�+���6�xY���8���
?I�z"��چ1�+�b�a���L�k��J����
�T���0�x�N��[�g��, ��i�Jx]���9��PF��Jc�d�U���ȳ�8A��L)�d����%R�'�^�{{������ʟ6B�&�{������{�v+&�!1"��� �!�.9I��N�#�˰խm-dI"��y�w�;e����c�D�~5Kns룹=DQ\�|������!��V�~ju�Ar(����^����u�x������=�b�u�����Vݑ:X̿i(�%\� �d%�''Ri��Oc�������W�:	���3Zqx$�ǐ�{| �uI�JfhҖD0g�jN��KY�a\:�|��V���h�ޒ���m��A�5l��:u��m�0�j�%�y�dR�Z5u�ʹ�!���n�#.�ihL�GF0}y�>�I�7�*��.���g�Y <�n^{��1[ܩ�,���*����s�d��`�L�i�����e?Y�U�W��X
�%����tn(_��&3�9�v�A	�@E��~/U����rs#4:ɛ�ٺz�[�4wQy���4��UJ} /�XQx�>?Lv�Y��ȵ��&��G����\9�y���A�����h�{��X{Հ�N��U�v�R���8\�G��������b���=��گ����S;�a�F��:��W���(j����{�ro�"��iN@�tFC���&�-�oq�_��7���w�l�b�(=���)���������-?ݵ��8&�)3��+~a�u��Q�~��Y�eb}o���f��I��]d���l�s��c�����~>F܎"o����AJ��
Y��?c>?An��KL��dY���d��E�E��yh,�I:�u7GE�2��+u��$U�|K� xP�̈v�P_�+�u�d�wU[X�E���F�(v$�`Q��h���Hh$�B�u�l��I��gc D�ku�,Y�F��t����q�ffRWƯ�6����;}�@ȕ^K�O\��0µVsp<��>�G�J���+G'�o�ZA
GLf�ǈ�(�rϰ�8�A a#b�F��Թ2l�qs�i�^�t�^ҥ���b/17=֋�xLSCW�=k�]Ԥ�o�2��@r�� �2����!V��0��R����-�3[ko��s.y}�A4B>'�v�t�����&����6���_5NX���.���У�)~�~�����U8�L��(!=!�In^Dۮ����Z��'��8"�U���7�\L�ei�����T�>�y���a���C����\�:|���ԆWUo�-*,s��(	MW�RaH�B X}2Ŗ����𭐘CLl���*5R\�쓟ǟ�eW���^J&�X��&e2T M �\_���q��w���.Kv��+-�D'b<�2_@QZt����C� +�zk�E���h�N��>�����liH��(�¾&E4�R�e챑X�f�a�6����^�B�V.*8~���F�c�6��u� ;��a;U���Ǧ�î7gVk-Iz��r���ϧ�?o$�^ilk �sv�^�w����+̱���H9��*�~S�ݷ��q����6=Qa�>��y�%qi=�2}��0F�(8o��$͖���������vv��a��s�~pmҀ�a�7���Csq{u����f�]�EL+=^��Xj����X�;X��z%$�J^���8����S�O�Ϣ�%�R3����J�
�%B�ĕ�(�����9v^�l_wbUu�5U���}��Į�¦�
���n�!ȤUF
ek~��/��G�e��F���]xk��f�Bs�7qT�l[	i����Rs�JG?�*")e�����8(�M~��f�;|�4ǜ=�`��m>� ��\�O��|�;�.e�Q'c%�z9C���}�Z�+&Q�(Ή~#���γ�V���S�P@��S"*< ��%���p��9h��Ӻpۺ�Lw���-i�������M�|O���R7Ȝ^s3�{�>SH�G		�B*g�6Por��w�Z3�48gj�����\�6�꽫���6�b����Mtf����Ε�V�W!�k��kO�+�o������/k�����K82�����]R��r���Z�o]F��[f,1 ͽ�IX��r/]4��ǭ�iFdg�U�Bt�z�ô��6~���%�jo��KͿ�RI����^�����4��?qB��"S��R�9��r@]��y����w� x�u
�7t���S�e�wL�z(�VD��;MN�fv�%�2��������n���TZ&�+iF8���9�>z��!�k*��������F�:9KZ�Q6�C���D��τ��(!d����#�
��%�Hd����
()( KyJa�];B�R��تC��s�1�{�X����` �+�pyk��-����%u�lw�6;�o�����|T�{���xdǄ������t�"_0sȪ0�~
=եHK�����	��@���Evj�ˬi��IyB���8i� "sv�����փ����)�T_��y0:�]Vi��1�/��$��,�q+#�5�axz�}b���3o�3((לRE>$ۣ�Q
���!�oS�~� ���̤�6MPE(|��!�M�>!e�;��K�Əx���j������"B����!�>}=����,������j�3�N+�=�?�a�`�RE���.�w��x�z��xmP� ���5� �W6cv�Q�G7��h͚�U�G�.�����p�t��g@��f�Xv(A@�3�ltw��-ǈ�saZ�m�#��l�`RV�� !�K�t@[EɃ	���d�X�uo�R�ӝd��'��\ѩ�����E(hrpǠq��Ȃ��`��^	6���w��O�#GS	Md� ��'���]�ء�*z8���Q�cPU╂@a��"�/¯��j�ly�-��]b?�n�E?st��F
ʹ�L�e�q]�pH��2oNj�����f�0 ��q3��_�L�D&W��dvw��������~�Y�P����Tq�'� �Y�m��W �_���SM�ʚ�\t�P#J[�K��պύ�ȡ�3Wڃ�4�1x���YJ����o�����{��,6udj=Dj@(>g�>�_��O��	��3`�S�D�Yn�.���lX��pE�k��&��z80�U Ou׮����Nz���3si<A��ٝ8�ۃ�q�g����kG��!敕�p�7θ�wP
�������K�ԕsO�3�:K�M�V=C<��h"����B8��C�g'��V�wf%Oip�@�枞ڦR�o7�6�����L����~��3�O��w 
=/l�>� �y�ڎ�����!;�N�V�>υ���V[_�Ipu}�U���*��-��6W�M��ϧ�b`�8ň3�O�7b���h3O{6���ڭB�(���G��=��}W�r~\V��_�l8��R�}V@�m�zܸSGJȔ,�K7Hȯy"帬��SV}D��_�t�R��-�_�Lg'�s��ǂ3���3����;Pr�W=�|(%M��R[�� �.+�9\�:�Ih#� ��ȗ n����1"�}�7����I�ܝ�<U�C��vM�C�#S�ꚼ���y���T�ۣ^cB�`Y)������Xls]�"�e$�\����%��H�1��G�n��p0����%�JY��NQ�R�% 4�q�$9���k���oD��*
�KI���h�=�8y�8�^S-�:�v�7�'��Qv�Йg�F��G�<q�e:��gM��L,�m��NX�GM�@TE����S��-�ƫ�\�Ug��������_&	mޢ/���슖�J��Aw�m���z�a����p��+=l��u��3o�[P��Ii���L��pa_Z�)�#�dS�ǥ�*�x��*��_sB=��6��p&6v��z,��s���m������į �^Ϣ�q��j d�mT/��YeAE(�F��S���J����1�h1��>�	V�W:=
��ΦM��"����+���c�,�:��]��{=�Fy'-����q-��O������#�.��nH]�G�k���鷧\<�%��������Blo�c^pe�m[\ژ�^Cm�Ufu�(0��E\�̥��#f&�x�ݑ��!}B<U-���ɺ��U�hxʆ�I�f�3�K�G�A��e6� ���s�W异�L�\3<�1sN�����]b��]�7`X��儮L!"��`!�J��e;��&y�0�\���FM7B]_����,�Bqk|�4�ů��Ȯ�אLv�xg^��>Go��C���k����:Ϊ>�*���f�G�F�����j��@���g���,��X����d'�e���퉔�'���#�q�GɄ(��$����B�O���I�O���8ׇ2�Q�ר�O�Z_���>�<�o*d��@?]s�԰��3:�C.��Ld'y�����:�bm�@<}K=� T�? =��}����FZG�{�CO��lǩU4�����;$~IAw�RpGa��@��C؏7�d^��`�3�qą��ʂWHi��U���iZ�7����B�l�2���5�h��P�ᢧ�yĘ����.�c�j ��$�٠�K����>H�v�GEUO+<l�@���yŠ��O�Ϊ=I����/AL2cqFK
Ml(��W[{�Q�$��/g�,e9�;B��*�j72Cղ�Q3���Q�����#'�6­���m��%���/�^����Y�|dG~�ڰ&��#Ξ�ޚ���Q?$�}��Ь:�/n����E�x�He{O�$���h��.[�a]eТX��B����u���=�Cᖂ$/��ʭ��
(D_��8i�m:k��ff�Z\�X��q9��y��L�M=��K�0�PjO·�S�N�%��C�٥~�{"���U�J��/�m�ܺ�L�7%����!�(n��F[��Y�L�����&Y��[T4��W �3��yQ'3�Z�w�
S�B��aw��=�5W���_��?RRW_%�A�G,�3��b�{�Ƽ^�� xk�1�"lZ�#��ܕjA%\٥�*���?�U��HN�(ܗ�lVT<�Hirf�i�8/�Λ1!4wv`ܗ�Đ���\�h尭)ӈ��*�RJ��ȲK�t7��c��_m$�.#]����҄���[i�����A�͟!���x�T�;��҆�3�l␌~J��*�\1B�;��f���]����%?^�d���FZ`Y@��������VN��@�u����k�%�]���L���S6�	q��������7^�����>����E�-��S��̏n�3��?x�{� *O�!"&c\�-V���W�l�P5>ǹ�J��7RK`0b���᫸���Ŕ�T���yiW;<	_����a��S$L����{���B3��q���Dr ����B%�J��j���j�QFkR=�n�r�wb�+�2�u#s�5��8�	���rL?��'�Y��Y3��`0�"n|����}9���C��PT�Q-�x�Ru��VP��/]�xG�wk�O<l��g�b����
�%3��CЏ��՘U�d��?�ۄ�dՠ��Ykν���H�5��?�CI����9�����a}E'�&�MBao
�l%x����=窷��Y�dx+b�fYe>���tM+v���n;�\�A^5�K�DN�;�Pp@�:�O]0�Z���s��p=�[�@G�G��9h	�i?H�݁E��1�C0@�P4,2[�'``d,ӾQ�%�-��nk�5�ɹx -���c����h��9i*��V���P=kd֝��7E�f�^���(�ɇ��h9`�
�T�;��n%�p���(p�\�C�벀�hA���hkt�9D ^��nz ���o���y
=ER'��NX(9,ZM�OD 56>�-1���k��unWϿ��o�]e��QO7{��(�~DC<P�T^�{�B3e�'��-����J��on�zH.�[F�	B�8"'o?��\�[��"��|��
�3�n�� i�$���TGn�C�!ŮQ�_l��N.N.��X�^�_nq�(���U])0�����ο<%�t��ib�5l/��r�5�`�WA���,\L�g��V�E� D,�bI�\̒s�`^w�ן̻'0	$B����t4T�;;q/��)��4��cm_!i[��d�,���� ������%��/�H����`�^(/������Ȕ���Ki�*�a?��<\���*�}��~#L}"p���p�aD+1H*�^�Ӄ����y���'g��8��9��7��
���O���#���م��R�3�uť��'��"�)w��p�e�Y�9.t��T<P)S�<�쪕5w�������y�C�h5rG-���y,w!۹5���v�~8��{%'���J$�WP QIDn�������{���Ff��{��k��M��`����{A�_�L���Td�@;��D���6�q���G~}%r��x±C����r
��2�;��d˷�k��>�E"I�iH���/'���ŧ�¼%mȄ�u������&���ldcqD��d��O�.;�Ƿ��,l�(Xy�3��x/�a����n�\ʦG�E��vF�����!�D�fG]j��L��G��-�1���J�Se��v� O����1�Ǝ�07D���<j'2�!��r��j錖nzk�n�k�7��&��@��)�
lL��m�\�_�0��*����Q!*s=dl(�O�Kv��	 ����l��㖒`������t�Z�	v"=,S�Q�<\H��;d�ɗk/���j?�y��2F�z���K����Q�a�{K��P�C�V_��QeK���Y�KbE���#ݒg���V��)7^����y
SJ��Q�� �پ΢�7�W_�ށ^78U�G�����vBK�jvn-�߁��eD�4$�;U !z����Qvy�*$#ْE]#i˥ǀl_dT�;���Z����T��,]�꯼�B��)���H�=G��o��W��.���
���������AS��^�j�F���N��������Y�#Z$�]��g�/|PWॗ�b%�R�%-�Z��Hݡd=zbV����o�6�R�:�'adw9D�l�=�O*1�vb%Om�D�F\D�˺� ��e�+F���I��!�9�j���ZR+&2O��ñ�Ѵ��A�����<۹��÷�ɳQ��Fď7���Rje  �T��eD7����[cP����H���˲��
���t�9�YNYJ�h�>�b�P�,��p/E�~[
A;�
ͺ�^����2R|�M\�债���ɋ~<;"k���K*�E1k{�q�n:�q�/��b����p��L��l��H�C�>=/����\&����N&�>�׳߷����
"C.�3�y�vljw���|�����{�j�#��Ϝs��L>ի�N�C��K�Z��J�p����]����̫��� �3ݶ�j{�@�hU~N[}��v���NV����I�1�8;��P�:��(�=���s����QR�4���!�mbA����w����RW��f�̱�z 73���	姐��X� �Ε�."jT�jf.�L�"��[b�uRF��/��|���>4��ԅ��i�'��9�4���V��t>]�
E\LP:�By��nJ>I����x��ͯ�zz�Gl.���9g��N����ܫ+���CG3�Z��S������Gc+��ep#�נ.�1E����W5����a��C�z�4�F}�I�˺c�*o:���faC_@2�i6�8@�y������=��{T��m�Ƒ�U~�'X�9�m��N�����Ҡ>�p����~��D��]��7���q̑�.�<��ˢ�o�4�ԃ׼���D߂Ҫ5yi�~�X�0��X��i\I�R.݈
U���:JT3À��a���Ǧ��늲E���ý�� ���9;?���[�+�I�����L�P �7��D8��}?�L{5�1��<��[Q�/%�FZV��)r<J��$E {��ɡHw'G���΀�˟Jw1����G�)��	-���j���,N�j�za63����?X����d��$�]\��D��K@�����(p!^[�SȔ9ѕr	\�}Bb}����-JP��C���ƶ�j�"v��/�voq����1Q�p�d)���a��}Hs,��5)�ɒ����r�Z$�?��zW���@�v(M���^w���a�|�h	�ֱ����4��o�����w<o�!Ajd�t${
���!b?���4d��1���M��_���Q��7�,G���M"T�븪R��Q�����9�U��������-��֎���-כ��M���dk��K�\��W2�ۑ��{`@r���$������Jx���rN��.�z%O{�ϻ_�Ɂ�gR|���Cb��G��!*�ƞٱd���"T�ka؍�T.�h��,�Д��p(}v�Xq#o���5b�h��)L8"d��v���&�v�2edez4�P��ݪ��{�2���I�e���)�٠rl�K0)i"��<���^	�SE#,����8w�=K���m�"*0�����N��{'�;"�]���Ә�	�T_AB���mqz����v�m�˽_)�Y����C�����w�p-��0㖜+P�W�':\ ^��dO��B�]E��fLp�o�b(h���i�u���w�5tJ��b���b7w��"|,�%~��v#�F $Gtl �r�� B;�<�Ǡ�NA�v/!xP�b(�������FO�u���5���rW��"OЋ����w�3h�)-c�ʔ���- �Ve8��á4cԄ�6qE`�sj�����-�̪8�L�Y��4J�}KX-K���0� �-�s��Ko�q�"�� ~�S�Q�����þ�'��i�T�,{�9{��K�L��*+~�:�HF+����X7�%��U����/U�i�A���u>f�8�1�n*b���V�����r�=zQ[��>.w}�N�t�R�]9NW#Of������.0!i��<b�Q��@������ި����%��kZ��W��*Rޟ������0:`��4π�B����~��]��X� .*D;�i��-�zV3=.jy�]�Wt�|j�(<�y���a�B(C[��I��j%A�-V�h�XP�u�].�e!6�8-��g�T���*�|�>���3L��92.
�ߟwsި����?��'�}�?\<�l�϶@�n���3���"OG��L�AX��Ci�\"�_4��n={6�I[�d_[qb�̓H�b��zsۨ��q�լ�/�Ri�;���T���?V�/ �{*���k^��b����!6Łc��0��"��V�I(��?��Җ�VQ�E���=��G?�D��c��\D���ג�D}��O�m�HN�O�n�� |�'���U�5‾�Y�1Ж��h�X�s˹�ʡm��;��a�q�H��bHU�G���
�!;�fhG8F����0
e�O���u���̦Ѣy��-�X�a���Q{���[�7����T�}��g	�]?�;ݓas��i�IE�Y�����"��Q�rjq����؋����<�(Ҳ%Lt����g�6�+/<ۍ�!n�`���jBm'�aw��e�����{�:�/��[g=�'=]�S��Ƙυd�.�	8�PCiv�P��~�tM������U������_�H�aD�<�hnW�HN|F�����I�ԕ�?z� ��?�B|����qНV �8�r��/��B>���س*C�N��������Z]:�$������J6��0��M2���%���5�>�4o
ykSs-�p�����6e�BS�:Q�(0O�0�t|r\��$�Ϋx �ll����S-��>n������*=���z�&�;��V�G;�+�����w=$X�`����3�0�Rc�V)�OK�#��Լcv�{��'�4K�iW]$�?��ߢ��^׈?�8h@�T��p�Î��v��!�������,�n"��ig)�k&�[TX܊�|3$�*k0���s�&7 �p��:)�k���s�*�q>�UK��A��if/�p�4u�  58u�@NK�&�9�rg�rߥ��e��#���o0���ϐ� �HYH�bKF�,��2v)&<S[��'?[zA6n}���3�Y�V�W۠
>��s�f?����ٚ0���|D[}+�)ҹp+6�MoɧKJ��YVS#�v��6_�2ی	���$R�����[Q>��B�m/)�";��� up��O�qz�*5S]�"�H