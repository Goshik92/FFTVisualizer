��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�uwC�5�b ��ϴ�	+�
Ct� "�J~���z����<
�����'k�z��ߵ,d�.��Z�Ӝ��2�x$ҟdL��h��ʔf��#
����;�;m�ȋ��[F��E� &'{=u�3jg�b�)��LA�u/5{<	���ʂH�__�>g�{fԛ��
`�[A��Q��/43r�� �K4��<��{u*�b������� �^��F�?)�ˮy5�H���<Y�"u��Cg��/z'��������(�pr��aI�b%l�������^�F������Y� ���K�����=�:xjx}e@>��r"��UY���3���ݘ��"ͷȁ�z�� �s$v�����g��|O�Kh[�ceq)�"a��4S�p�qj�M��]��|��'E����Я+t8't�떭Ä�:��%�����^<�Q o�Sh�r��,��ifs�>�I�PG�u��l-�,U�W�t��z��-�I�$x��U-�s^�?����]߁AF�P�����ͱYJgG֊elg{�M� �w/�ӛ����euG��+�qr1�/����q424��ˉb�zax��J^iǯⸯ�YK������>z����\p*�q���s�e>���ϗ'3�ǅ����.���B��(�9�3��=���d�3#+(W2�W����a;Q��y�x��28�on�P#	:b)��bL�� .��5��,C����'�)m�ÞO��D��u��T@�RS���4�*D��os����u�X,_��#�z�wcM�İ�\䡟�Ʌ�f MgU7z7t9��두��7�����V�J�ǥm��3mH�+Z�����:W~9�>sK�*��a`��+��*ܔX90�S\�Xh|j���Z���^�}V>P%݁9��%�t"2���29g�@q�M�U/�Ra'�tj�T<?�����@�B��e}h^�e��*ѻM}�����D�9t(F�%� i�Gc�0�����*����jv��]�T���E 롅~��1��H`A�9m�n
L}�Ó\���Ѱ�����2�$[2�WO�}�3F��<���߻W��E��8> �uhN���f�UZ�m	���O�㈴L�c����ӝ����k��K���r���8Q�-��:��� ��{ ���/ �9�);��.S� F��!_4�h�y�_F�~��6e\���rk����~}���r	�p<�������
k��2X�pUQ���`�y����{Y���N-�6���H`x���ہ����:�|�~N:Ci|�3���9E9i �����s4 ��P������{(N��|��'��Oom����G����p�}S)�]v��1d����kegM���c-)�%K{��g�/�O�q���t�2=@ݝC��'~H����P��-����0�F�甗\O��r>2�"�ݚ�'t�	kGזM!(ᷡ���Խ < &c�	#g��5M5w�9V�[�ӛe�MК�9s���8Ի�� �&��aUջ�8�i|_���{�h<�%eod|����iG�
�So+�Y��>�)e�аJ�w�z T�����v|W��դ]��UjGfF	����79<�CI߫5���!wu�Ch�e��NCr/��)�����C�9A����>�W7Cw%'�b��m�D��o�3�PU�u��6Ŵ~][d��;����)�W��t�w~�'oJ��q��sD�����!J���G30�P5���ʥ�	��f~=J.:��ƫ�uW@+9��$�]���'Fѝ���\�sS"�;�:��ɂ��",�M�E�䶹��m��I�blf�H��I�S`ע�М��2C�v�s�FΉ�M�f��[�@������乽���[�ù��0 F�U�3s="5_-)L�>���J�Ujq!�p��h�$���O�����R_4���� �%2�;h��m��T��a$�N�� 踊�$\%�ۮa�W��-*$�' �e?L�C��u��;�2��V����ԙ3���U�?;|gE������2��S���_�o��ۮ,�2���/+,��C����y�ڕ�xZc��[��g2�������8��� ���Y�.`�p糱� �E���i�lE���_�Ngi]'�X��aM�q2Sc�F�D��Cq�Nw� ��=dv�������<������ D�g� B���w]��0�s�;���F�ɲ��}���ި~2m?Ӻ%K���{��؇��EXt���(V�������A���L?���߾n�^,˘��Q$�D���C�3�x�fM�j8��s���n8BЊ�=3ݡGqú�	(u׿,%�Ȝ1�z��:^.�!~�S��e�`F_��}�q���- ��<��$���5�1�$= �"��̉���O8gJ+	&��&��m�L�|��[��4�gH�a��Oi)�Z �e�(vjP� ��2��K�f���D�~iRH���i�(���P؍�����S�$�n�f��c߬�TR�f۽�J�!�y�-]��>py�|�X�����؃U�`�L C"��'��S'��
�ʜц��=�0������Ay��������q��~����ō�� ��2�dn����ٖ]a��H#��x���w)" ��ᒴ�	���NW�����4�@���ɻ/Wnq>})�J�0��ϱ�O���	�;uP]�h��N���h��ЎϘ�6?߮�����,�G�U~r��	w�l\>��/�_p��l[�i
Ā��Wt�^G�᡽~ȉe�aG��
=Ɵp5��sSzdd��s�e���+o�pu�J҃�߅���:C5 2���$
��MQ��ԍ�$-81�d�N2���
Ob���1�X�����!8yE c��W���A>=~76���h
V~'�?�7cۂq��
���8���-L=��n�F{��{q}�_�옱&p�#t|�-���;^�"=ӻ�W=�e�[�R󠩘W�*V�Kxk�MFl�W�P���1f�����~�$��c�y�r.�C>��oa���)���`'�����^�L6(�a^2L���V���c�B���!�I�9R�D�\Q�Xe^�ɓ?A�������z%%NMpC<X�)��I G%Õ��2�b����a���fK�����Q�����f�j�u@E�S�����u�U�l��|��>߶���x�~�-#��T��xs�V&���]�,<	��H��������p}X�(;p��u8O����%5���
w��gf��44�0�m��_6�Y$�W���|�YbI�8_CJ�cEx4&�CCxH6���ETG�0�������C�@�I��w��p9\�P�o�ڒ����I�c8xL3
�#���!��)�������'�[�-́�dq�@��£��b��~��uɀf�DlP��0גL�����%t򋐦���32����s��� �F: �Qw7�6Q~Z4p�p��>a�$qn�z����oMSО=�sq;����	V�@b+��Ζ�Qa����|�nU�xX:�ڠ�#H�3�����F9�ڲ֫�ݸ��إ��k
����#R2��[���+��V��zȇ��S�y�R/�`W~�0=q�C�%SS��}�ܰ/Y	q-�'Đd2Ce��$��4����Y�*j���y-ط�c���_��mLZ�f�����n�a�	h�]:�� /PP�������_C*�:kN���A�ȕM�@��}o�rv*Z��tC~��@��-�#�H[$��V�::TT��hέ 6�Bb�7C��P�$=�8y�4��ӂX�)�_Z��������.D_^��[����_�_�<��\y���#\��������ʚ�O����w����oX����e���2d�ߢ_�� ����ߤ�*"a#�/���ϖ�L�K�a]�iѨ�ў��46��CW������¶�A�lM�w�tNu�\ �:����f�kVa��jV��WC�U̶�	��m\&���> ~����+wX	$}�#!��*�A����6{�_�rR�y��W�sKl �G�o:&��i��jC�����lQ�A�?�a�^C�-μmL�RF��ơ��z�܅�t<����9�w�$"_����`��ݴ�?)S�>�:�j�vCNs)ɾ���u�ʑ������ܲ�~��L]zo��*��3�E	ϝb�1��x����)b���TV��kC]���y�։��t�`ז����_0Hz��Z���]r�.tM&J)6[5�U8a�D��E�gf�֎_���:~P7�v�?[�L)���?� �y��#��&֚�� /bMwݫQ^������ń�����1��8W�g2��ET���D�FtF�����t!ڼQH􉎼}A,�A�gVaD
�vϒ��2�����G����@�qL\�g�'�jy		!�Y���6�_r�PVYJ��^�
2-�$�e�p��Ьe�|+���YUnY�+rv�,�J�X3�z.u�=vE���Sq9*6�K�9���jY���}*��\�h/r�s��j�R,�Wq�&���q��Ee 'ϡ���F��7Yo|�7���C�D���n#~*r�yv_��KF�Źcg<3�.ܖ�"�P����lq2��ƹr�3�n�aXG�A���M�r�9��%|�-F�&�����gd�Ő���q8>���;��4��`#��#%b����N6�c�Ⱦ�d.۪d���29�i��1n��A�*�L�l�2������������5�?8�0ۏ�΍RMۈ��`��a^nS���T\hr�Ԇ�Oօ�����ލ��#�V���#O�h��h�����XV;[��?q�6��L���Q�p_�r��+*����sY�1j���?�5�>�5~<w�_q8���r|��wG��[B\�9]~��Q�����V���y)��t$2��-�k��P�$����[�����b^<��Hp+}x��
Z���Q	��%^7��>�wIM	&���z7S���b�~�W�r��1!���\�T�3���$����z�a����#D�L<:�>� �����x����%5bsm4�k͝bUeu]�G�?��/>6S\�v2�(���jgM�$���*e�k�3S_1��I�ڼ
y�H��y�>���?S}!�1�0���[
�<���5�t�ޥ�j}n�K�kY��ި�,�[­�������5���<�e����~az�&mO� _Cð�=��I_>��_�F�>�vt��^w��5:'���p݉2������Dc����`���{u�?���Tu�����8��,�Q�
\��/���J��e�~��6 �Vٝ�1~����M'R��Ptw�7*�U��1�e��Y_t;��ܺ�i����T���<+S2��Vơ10�]?�/;�!��>�����QF&�@��6�#_���[����P�[��4-9*Գf� }�x�F�0ƀ>��S��Pr@O�������Ž�8�ғG/������b��s��4��W���c�%�
�ɟ����?�ƚx��YF����Qŗ'��V5Ɨx��"*���Ҽ�!��⒈���@�V@�p;����׼��/3��-��O��TN|MF�R "���?0ei�NX�Uz�����v�^V�<�7���ߑY���8Ҭ+��#ý㻬�\�
ynt���u��ld�]t�a��¡F�F�:$xp7�����fG^2����jjL	=�)�*�VA���������-]������:Ҏ���N�˓��M�fo�C���WF0G���� e��yW�=k
���+͌p�V7B�H��VR�sc�j��-Z�S}�"��}���~�t\!8⦹ഁ�z0�¯C��x���,���(-3����/E���8krNi�zi���Z���,ۆ����x��e�)V~��&^�����\�MS
�ޕ64cS�!k-g��b�s0�U�pn�1��q�?���S���A�Ƞ�&�(�ҧ�&�	.��`XiB�#-㢫l��Sj9�
3 �t�k�0{\�RU�d
�d�#\�%Kb�ݬjp��hK|T73d݊PRݠ���b*���_����H���@�7���;9�B�`%
��Pl��j�W�-'m��b}jb�������H�=��.Ι�M&��v3�!D�@�Q�k�B�����[�J��ʸ*��${�Pf<����v����-��t���K�N�b��>r!��:6,�O��Ǳ�͍JQG�i��S���ۃ0�����5��X�?5jns,>w5�����38���ˍX7����*i�5�"xȔ�KȰx�K[=m��3ځ8���F�rϠ��k�H���2����љ�͎x��o��c��^X���Ux����'G3�������Yz��-��� C���t"�T����}r�oY @P�!��i���́]�ԐL�խ����0��=��[����>Q�vQ�`>�=K��e��������P񲿉=� E���j[�d?����睯|9>�Tk>������N��-���'|Jt�r��P0� �=�9�I u� r��(�v9�K�mF=zy��v��"��x�l��	���6�뉣�EFB�=�~��$�0��4�}p�N��qmJ�(��g�>�f�鬇�m��rD�Ny������4�ԶUkɄf4P��y��Ha�I��_�8o��+�zz����
$^�4�.*a7��Nv���D%� ����qv5u|�����b��CA,"5T|���	�Gj�!LV{��pG��`����1f_��=��7$�\���H+���l8\c������F���cr�������-�L�[�"�W93���� x"C��?,�b�Y����ؑjauJ�{���QV����ފv6�������RK�-)��?Sˆ�ژt��w�����c���e� ���/V4�Bx�P�9��-��g�c���K"p	�塚K�B��L|��M�`@���r%�����!�7Q`�"`�o��O.i>�>��X����pʭ���@�<�%?bMm��*>B����>���]_6�L9Mb���
���@�F?��y<6�X�=���l���-u��Ϫ��uÄv{�|�/.�v�y
|FT"�#69�vBr&�>Ч|���/�����@N��L^ZZ<V�������FpƹT�;��n��|h�M���h�)S��d�1{���\Ã{Ah��[x%�&d�V��2��f�>�
��0���i������ͬ��u�<{�� ��y��#�@�_#��kI|�RZA:��/��4o��}a�-G�h"��A|2�>�ɽ�ʫ��N�>�WY�_�uy����*�����{m���Y��u�����#��r`��7ߢp��=-`hI�tK�V�j)��G{hߞ�lc�D�=��#W
B&5�`���4�V��s���-���A@��o�ԯZ���e���崝O,��|h����-'L������Tcq�Wƚi0p�wC�WmxH�p�!=I�l(UG|���Q�֒�f�������Q����_�tKS!�1��oq5��b����*�{���j��m7ѐ�B���(n�s���n�.K8:[	N���(=���"���W��ht�[ҕɖ��{�55�Y���;����c�y<����];�LDu��D���~�P�AY{�2�d|y��\T��a��e��ǶL��ý+���*�,��NW� %�\�������Q<il���=�a4j;F��K�`
���2��dVC�3�j���m�硛W_rЮ*q�OQa�"��E�h#���d<�{ԙm�CfI�B0��C��6=��6��ˎ�mӗ��dv�D�+�XB]�-)�F�M�Vnzo��	���n��L?����:!�~*2v�]'ǄC���g�ڂ�@]�D�lPM��J�Y�7^I5�;��K�D.a��mƳm���i=�}���8������
�5! ԍ����喐�,����n))�n9$.�/���j~�����[�x����f�ǯB ��(]�_�\�Mc9\����a�K��J'%d�-ʓ6a:��I�Wǵ��WSp\w���;��~��g췼�?��ʀdtp�����LHQ�R�bWaW�
���%Nt;mgv��W Apx���G�{B
��e�F@��9���j��X�)���E�<���Cc�#1��Tr�j[ٮ y�e<�y-k�p1��0>����9a���9bb�����[��լ1�E3M�R�ku;�$?&~^�g���Z��$��$	���4�@lL@-�Q\�̟a%(�L�	[��(�ë-�'bx�R�
�����l�r�����;h��;��w�9��$1��!�r���"�:��i-��/Bނ���'���ϸq����?�Ǆ�{��(�x+�W�{��Mg�p5��De7i��P�Rj�m���4/��&����'1;,����*^�N%�@D3��@��#�<�촢!������5�7!��m�#�G��M�u�2
�P5�SZX�e*�q�2Uo��MVEgw��]!s��Qsj�o ��7sFq����~ �X춥p�w`�, ������fz�� 5>��(e�j-�`	�����iB?Un�(fX�^Yp�� e8��"
 ܕ�q�R���+'�`@�f����?���zͪ���8$�m�6bT4)��jZe�V'�i�I
a�%~�v,�]B�V��ל�)��B>����Q|��m��A���ݨ'�(#�^1����&�?�rݶ�1��A�]7��ύ�� ������)^r���=��tzz��՗�N�+�-�F7@TtŨ�Iu�J����Fu����ܣ���XR+^~[Ȭ&- �L�[<�>@�Ewh�9G����˹0M!Rs��l<c-e�k.e�����y�A�I��l��x-���.8�}��	@gNIA��,�R�e��օZ�����0�I���
\�BU�ߑ���Z���Q���FF@���݂��
.8�[)����
�5�oaIw�ӿ:�Q��X��ط��wB{[,d�7[�$e5��Y_9���	�Dh���q�P��C"4�����������:6���Be:�Ks�ѵ�˔��h�'�>|6R���}���V \�_CC�Y\�H�L@V������?"�3+���`���?_��J/����3/�'�y�2�x�y>��?���m��� /��?�4��֋6�.�w#"�ā�ϧ�I����6;y�g��ɢ\�2wr!ѯ�_o���V��N�u{^dr1��0Q�9��v-'&+	'EMk������$��ED}��\S���l������G&ѭ������3��﷉�]#)�#���%���mjR�7S�!RL���@��~ñyD�� )S�3W���x4��������� ��`X�
�Øko6�D��H�8mT��������l�'�Cv�X�9`dɓ�8,���#�]ZyGCk}v���	��6%o���LCmB;\*�g��P�6TGo	<=��G��p@����ּl�)}�\�h���H�ˬ��v��'�c�톂��.]����[N�Z��ĹL���n����:|�������%�2�9�]1�����QR\��H�J��n��m@c�j{��eS�&��[�:�%eW�4�+
���s��ϤxTp�G�}�eBB��p/�R	���\��w�=�mɴ?�g�I|���lo4�ؽ������@ě�OjJ$E~*��WQ	5"�fi����+	Ѻ�A 0"(o]7�z��a��C�9ں���²cpS����Ν��A)R�8o�Ul�<lN[��̿�1$�t��B��{������B��-���'�E\�ž�uز�v)MH.��6�ͩ\L�L�><$���k
�1;�K��=I��ܪ��ovjv�Tz�s)�����������j���WF% �����=�0��Ї��>��5��]�)oF\0��
q�ǡ�D����mX�G:����y�/6{7-�:m /�a�*/BjSI������h�:�L����r����<D���.�����AcE�����NJ�v�� ZS̃�I�f���< �n���nÕ(�F=/(�L�G{����<�������2�l�<�B����B��CۡD4�Fg�E�|���ak��[��*�H�Ub�ݤOʑ:����]JN���E
���o0��Zz%�#K~����v>����P������|LB��\���n"����U�����j���þ`�E���r���Z^i�=�ˉ��?�~Msm=�`2�[k����FU= 'B��q�D�+d�M��K�j��ܚ�>����#wR�f�̢��p<\x�Y�%	���)�p����x���6"	�ȳc�ɰ�2F�Ʌ̍���h�#��F,�N�X8�M���Н{��^ !6l�C ub�@~��O8�T�9]zt�?���K 7C%; .A�G�:q@[�����1�iקL�k����_-GE���fq)��܄��Q~u[_���fY'Sh\���*�=��� ���yi��x�������4�����'�%��§���H4�Mkr3:ޱXh̫��˵�?��+%�#�W���T�x�E����uAZl2���a*�����N�[Be��X�ц^+8�D�p��k-)1˨F���%`
q7�s6�p�x����1̎C7d�E>����;��[���IP@��ܨ��̽�ߚK�#��t}	�����V���(��"�a�}�kB���!�Q���W�.5�j��� q93�+Ź6�����0)�Wf�)_,u��V���p��E�-�וK�̮���(�y�L(~�Y�ڽ�L�eA�,q3�Ҝ9��v�R˾�63v�n����S��϶��ń�CV��I�������Ma��!����[>c@/�>��Ïnt��@RK�]Љջ��,�am�G� ��;��v.�Ӽ�����6'��6�c���dDB�{i�qɵ'���Jfp��Bl��f�^���k?AD��䱌\��z��*����-��*Lmɠ�4ԅ1\xdH��\�}j��7-$:Z!pw� ��V)g7��n&W���Z�M�az-�8�H�:Y����jzά��¥�[c�6,��z饡�ܥ�_Α�U��pvS|X�md,k�?k4�X>�V�⯃bث�T巨9n�V˄κ-��Rl�%[��@9~@vש��Y�J�a5h�ej��؁��k�TwX�ؽ�+'�&^O����Ͷ���q[L~[܈����Hݮ)�F����*���Nѝ��R���r���Y�^�N��*�'n�};��`����@vZ�1*����fmoȪ�w1�z�l\��4`%~L�C�M�3�>���V�x~"�
��>�ÙSȃVv����G�O!��e
`	BDX#j˒�M�P;��	q�˾\����t��qo9 F��#6����2���Ӟ���9N��W&]�7��ƴM�C�u���nVG��Ec�I��Tq��)�j�H�B���3��,_[���h*#^2�kA�:�>s�l���lP
�l2ͪ�����g�Jt��<��e$�a�&A��Ip��"��ө\I�r��ŋ'�L
�����٥u1�2�L=���/s�6�. _�	$�Z�R,�!�5S�M,�-P
id:D���^A��t ��yJ�\�����9�`Kq��*��QH�2�\�_zS�c_bg��5;c� R]�����q���"= 
�Z]�	�S��q�:���1:�˯m��F�ƙ�^n-�r7��&'����F�ä��Zc���~�W�9��r�.�xi!��
��׾��WՖ�����j���N� �[j��o/?��ʧe�Cq����/Ꮓ�	g'z��	����Ne$��b����n�_��,q����ޑk���|#�X��H��tz߽|u�dq-rzm%�d[�� �wc��Ae	c����8JIS�',~�0���`��CԨ����hLy��_`j���f��c����m��v�f�>�mQ��k�^�v��6����zVɤu���-ѽ�8�yd����&C�W3hpV�,J���~�FN|~9�rʻ%Uc�
0zl8��Κ� \K�rmyD&bl���1y��rz;g����K6�{�*�N�� �~�2��=�+��n���P��v��J�g���!��$h9!�x~��ն����M�@= X��="�W�����A�{��cPe� o���,����Q�V+S��� ��u�[���ZE~�������g�Pk��dͥ]�J_������-��^7��3T�3y΅��jڝJ�	����XE�A�*�����i�-��� ��gb�u��Ps�A ��aP= �T��ՠS<�ƬZV�������M0�?�L�q���:�"�0GĴ��mT�r�w!d�<5��W���_���#�]1���Y����(��؎"B��)�^p\�BM�
�}Oz'j�����iǝ"�����TJ{���?A��|0#ӡ�XV$>���������7�:����+F��x97"*�d���\肈I�{_ �7�s��<�]�C�	����5���BTj���0 O��a��H�%C?��;�S�}�-U��I��z���o�aϭwµ��7_�ʬ�
y���Q� -�R�`���Ķ1x�}�Sv0'�!��?mv���2�S1���vZF�0���T(S��1gV�冶dća����/�lz�I�V��)F���7L�|�<�#y��Ռt�i�6M���
�W�v�q","�=���r��)}k�<���M�4����WT�h��Eg��O��r�ıqʳ��z^�v���S
���C�OpE͝ҝ��yi\��ڽ��=>l����p�;�Ju�]ѧ����^�?����l6_��l���9�~�Qz>	Մ��{���B�nM�MŚUX!�f��Űy��<Ė.�o���k
��%E7*��ؘ�ʮ^]"A���]0��&�GH8>zz���Ի���n�(Vt[�!��)6����+r;�"�c��Htr��:�A��&��M���t)+��]���{�����wo�� bu�$-p�qu�~�y}M��y6 �Ι8����yx+SH& ���G�_e�n��!��v5��w6Ŵq]���v*�vl�# ��������cNٹ*���UWϠ�)����,j�3ܙ�A�y�	��wbL�=�?��!nH?�y���*�q� :�ʆ�\UR	 �T����Z�|�Tz:��B�
��ˁ&�Ou{��A��S�==np������	�����1MQ��=sD���V�&baTh��_���
Igk+4��Ȅ�ᇯ#���V%g�3ִﰍ`�B�5wt�[�X�n�\�����(q��XL� X� ��K��s |�7�Љ{�%�J� �j�KUh�ܨD��\o���_���J�D�`�y���\��f�	�������U˱�:�4:����O)���ݒ(�{�5xt�s4��5�2�Ҝx�����z25?\nw_�E���͞��W@�׈����Ã��d4"��Bqyn�/��eK�v��u0�%2'�)��M�c?����3�h�H{ۿ���w��/���(B.�� 0B���ӌs���g*�4V�V�5�$7U�1��R;=#�8i��;� ������� �ʎ*~8�&v�ˢ�袡ϣ6
��v�2͟A�ş��П���@�C��j�ݸ�a!ׄ�;@
;�e�A:��܇�iÕ�<����$q���ӽ[PAZ?����Er����L/*"_Rc�&����7�>�H01F��8e���>C�lW���i�_� u��pE���8$��\E������d�n���E6,7xA�'4O���ѥ�8;�
�,>��ĉ8Ėn3�&;�DM4�4�թL�eptKv42(7l�`�Hiv�wr��j�H��ӛف2�@�e�{�:�f!�OT��:�]";d;m8cl1���?��P��1�*�E��-s�B�̬(�
�Z椣�|azA ���<2)M��G\�ڇc���z�u�y`�s�b���sq=	��ב��8����S�(��j�,]e��()6R�c�1�nzgHf(��?�z�l�FN|�̱����p鳝�[�8��^�$T�>� ���������J3_�ĕ>>ȋ��Fj伃%���Ĺ��mM����o)�	����S�H�kx_|գw��J�0�6�K���t_�"��|���/H�J����$m���^� ��2ҕ�g�޷#.g��}�d�{��E��1��!�As4�6BC�H�:�ga �~P<v��N��(h� ��wnD�z"0�J=���v�X�|�"��2�?d�
�����F��m����?bn����;TE#�5�͞�_��*��Q��'f�v"�T,�;Tnv�[�e-b�kW�J��]�a����V>�[��G�!�+ys�Ҏ��ܼD����PBü_ [L9<�_r|@8֋p���]I�Sሯ��#�"��/v5�<;�+:���"��#��FڥT2��c��s)C1p�J�����J���k��%�@�(rz�4y�o7>�)�r��1Ě����h�R{��1'fi�� d~�8�Y�N!�/��3z)�x7.�`Ӧ�U�\ۣ���z�T��HV��>�Mh���Ё^Q�4�'�q���
��J�,*#S�.eD;�C�0%_�Ey���I�'_�h����[����3���y�V??���/�%	�fx����~�@�;�x��*7������n셜���b����Wș�lZ ��d�)n8۬;�I5yſ�[FGI�O2,�[���?M.�we/Yj&��ݬt���5R�Ate��݄��n�����=�Ds�RR���X���H��AcO8n3�����s#|e(b�Ng�Y z^����%�:�OUE����u��Ӧ��Em�VYI�1�! RC�������H	�h��R��������A��Q�\�mt>/�ַ�!���<ҠrV�p�ҳ��<g�<����9�8�QJ��I��R�z�{׋�zYr�o9A�y���<�ֵ�cP�*� CO��w*�qB��O̗�FG a"������-�C��z�*�iҮ����S���v�����Y�,�1)!"�\f�X;y���%vw���ڤ��
�1o\ͧ n�3$�[��pLV�D�m�m%��7M�g�g�ˈ�T��wcx8�G7ׯ��̺_��@[�o}b�K}�4��Ğ'^���"�F)���Ȑ��h�H��d���P��O�����7���X�	|i�5e���0��qբZ
���آXf���k�5��Q�w���:>�>$q-��[���a[�7��cM��1�E$O1/�=�	gp���Y`xV�-�����:q�"ԪY�~�*��l�5^���&T ��4܆Ee��uS��ܼ�$�-�1Ĩ"���-8W5�+^���73 ��_�*�k�	T�'X�֢o�;����x�lm��鲂�B�]_/��bI9)qBK�df�k�����ە���Ԇ��`C�.Pb�SI���=�՗�zM�|�G)��G?5l��,�~�>�Þ|A���:�e�?���?� H
j^ۨ�4�7$|m
Q��#�ǋ�����,���"* �ps��3j>�F�A�2/x��̢���Za�}�x�X�YA��GW'�0k���qp^b>�p��|��G���.�ٖ8�7j.1��o��_?9 ���ɪ�N�9������>��[xc)�d��Ww;
	�]A�Ը䔽*By�����9���d�^�L��"�']0���#H�T���Ǆ�������@E��ޕ[� �f1��⠨�{F�멸�N=z�f�07oN4�h�X@՜'��W^z�@2	�-©Qً�,�y�$d	�]s)?9њ��Kk���X��y�\�}ipRN����EV�j��m�V*����M]j��F�RM�U�P�;��r���jA�u�;���3�,�4(��j��A%#�L�Td�5eAO��&׎��rdP�X�G4ܺ��+���3 ��0�Л���s؇�㒻T�^(�����:�9F���5S�Ei%��)�lD���8U:�E�.K�c?��7���xB7Хl��US�3_��(xa�w�N)�����k���U�.Tk�_hm��e��mE�K��<N���
>�5�h���Ȝ�5z����[q֓����Lp5 /�:����^���q�=��,��V�x������Od������ˆ � Fҍ��!�?PcF�Z!l�d����m ���oʡjJkV��9S�Ư|��mx�������t���0�e;�����2=t�9��K�iz��.����G+�=w���տ;����XԶ�9v�Zg�t�-����\��-�pw�Z꼶�e>Yk���j���e�0|E ��h�^�}o���Z
�>��]5D
^���š����J��Gi��D���׼���CHǬ���p���V��1?�3�<�w�X��k7��}��m�>?��e��U���Jd?u#%�UUٜ���0��m떰���	�ᄌ��ѯ�f���jmm�9�����\g�&<�3�oŐ��K���&�8�2�襾�7�tz;̖]i�M���|��m�EJ ΈXuh�W��f@W��O<t8��|#���[�b9��N�{����qš��>�C����r�n�d�l�!�$A���1Ǣ�;[ۚ/�᪁�p�	v�漅VM����4��[�ü@��L�LmQ1�T�6P1��IP�>���Nz˵c�WW�����T�D���sVrM����X(�+crQ�A�M�N���Γ�A�s-���C<ѥ�"7��K���ٛG�E���%�N#1�����e��#6��:Mj�7�N�oZ'�<����OC'�m���j�Ģ�7�a�Pz�����V�d�{{˂�lZ�AO�YuNd����*K�>4� K-2ꄔ��Y�8��<��"�1�g�r� E)GD�a�=�h
�DY}MH�p���)�W Do|�2�X928]I����{1Q�T��4��PYh�T`)�3�q��8DZD�������0�c���?z�o$�&Z�:━��Z�#��J@�!�D���E�QUܜ���bm"۞��ěg\/C�M��?v�uR��W����� B�##�*�����'�[�D�s�Z���.�oGWؘ�
@̭���	�tV��A�T���$���^��ᛤ�J>�Uk0B@,>mU�(*��]��CIC2�zBm�=�i!�;cx8��%��r��"[�=��Jȑd
�&h����NT�4�ǣ_���{���F�z��N�g��B��%O���E�8�y���Λ
 ��*�V��*oL�����/3Ǖ	��CV��j��y "̈Y-�1�J|0
Q�Q4Z|�Gg�C"pbF�7��3�n]SZgy폓]�'����o8�Y��1+(������tf�=ԡ�|�?y�=~j��E2� ��=+���R
js��T�֔Ͽ��2�E'��jYQ�`e^�4lo��P˗kZztr�3�*1	w끁Q��C���Eǃ�+U�#�'k��6np#oR�@�"����r	���5������HM�N�,�Qj����7�Q-��MA���h	hx���8�\S�-�������9�ZrF��mȮW�%�fmG-�y���{�ן�%��hg��Yܿ�HZ�Z�c��nTJT{97���#K����~�_���$�˸Ζ_�����W�R�x�f��ږӶ�n` Vk6������d��Ș��wa�܍�"�4`��ZB�6����9{��%�:���I?�c�JZs4=����&�M|��}t�"�dE���]���s��Aӣ�;]��d`~C��&v�z4 C���ۻӔ�JXB��d�J�ys3v���L�pe/�dF�w*����^��AÓR"�g&�{��5Q���A��"��L��Ň���̵��'Jw�{|x@�>��U@<�@�l��
��l��i�d�J�VMT���X,W���P��y��S���z�U�[!�/t�{�/lhnl��Mu�(��,>�T��	 "�.0�Ӏ�F-*j�����(��\�.+�Lp1���^�!6�l�iq����Jbs6(�;�PAKd��WBQZ=�Ur��6uBo���̻
s�`��(+ya3�ǟqf5R�U�y��#�(��G2ì��(�IN<ڔ��6�S��qᰲ�XC$�A��;z+�zח��8oZ�;D��z��_][O��N��f�R�	�ffe��[���3�"-�1	�3�
$�����`4��3?����������z7Ņr��G��Z"�/�a���\��NE��9�N� W}i^W�Ҷ=W!E��S��Ǭ3��)��q7��	�z��G<�)� ��f�/��ZѳB�8������֑���A$�]5:�c��݇l�3`��/g�&��L@rsO��;=Ĉ���7TB����K9��C�=�h��@��'�ſ�&6���3���g��:;����
^���q�����%[Z�H��A��`�����`�-�!A�ay�rN�HY���F����}}w�5��ѺB�wL�Q�^1�/�1��Mͯ���=��Ǉg"��	Q�V(�Ą�-L�=lG�[�b�H#�6!�ݐG�,�^�< �v���C{pc�����I�i������<)�a���� �g gǷ�t��#���1��d��?6�~��;�ļ"m��e���4�c�ZF��N	�1u���ܨZ�f��-ei�aa��Out�zS-�Ll��ɮ}�8�dD��|z���.L	��gH�]�1̝��O&��o���t
X�<Ko�t��YkA�f�S��s=Lqu��g�f���,�s�3��d_&<��|���~F�p�"����!��+{I��?/1�I�B*�
3j�����}g��q8�D��I�9,!��ng�����q�C�2Q���@��,���/��� :�b5�K��Uх�c2�j�����8� _���w��&L�H��z�8�dqQ�0��~թ�?r �򗑥��Qr���m3�.������f�)����F?e����pư�	;�I�ae������t�Q~�s=4,e����Z�R��(~�^� Ov����9�lv޷����B���Ө���cH�(o�'�����w��/���y>��-�{�Y(a��3���_����!�d��c��Q���Y!��E�H.�a�
���{�3�%��>k���i�=������	�Wĺn!_{bK � n��N��,?$+(���1��ٵX󎜥����*�	���$ƙ���*-1�H�L8��D����ѹ���Y3�)��+uo`��LM��ׇ�z����m7t+�Y!b��]�5�W��>�#�x�50qK�zv�Pv清�s�:�Ȋ�PAceD�h��+\3�v����)�57OW��Vz��qP!/(C4��j���g�V� ���ڶ����\��X�[:���?�#����UR!������F:��U�豂=�/i�ƅa�����aFOc�q�Mw�_e΅3!�h��H���G�Q���H���B�پ>$ڹVGj�j��s*��o;pO�@~\�kS�쩞�J���?�w#5Z�¦�֒)���r&4A�ƩZ�;e��h���n���ɶ�њ���Y���g�/�o'$�T��_"�־��g�t�/3
s���Gۃ�%:v�-<�~�M�M�7���P�WSD/�ש���7�ִB���}J4��i����]�#��L�*�ʤ�����C<�$��Գu�>;x.����l�GE��U�vT�J��R10b8���_4y?�|J��Ox�bd'��D����<�އ)��˟���N;�'c��'h��8����n�@�`9d\U��(�^�U{� ��Ԝv��9���X����I��HY㑴��K��dO����`ӻx�� �8m�Ա�x����ˁa)Y6�׎PP��ew-�������,3ׇxe��s!�L�G��$�'@7�aH�0G50�:��8bBk�9�Є��|�4��~��5!I�uћ�f���"H�0���U�"���� ��Z���H	Y��3ؒXhZ\�=_��1���� /35M��}2�V���Y�s�DIK�ՠ ��-ѷ]�)�ieK�4���k�_��)�2���_(��r�y�?�Q�Ϭ�����vۗ��c��h|b�@U�A�����\i�=����4���ھ	����"{��Д��F�E�QhHφJQ�S��
�1��!Ĝ�UE��������|�b�}]��7���2�"�%
8A�'��=��c�.�e�a_#&�P#IׇF�";�j�N<{yơ͏� {~��M�	G1W�W�,�����cJ�:�:���x%7q,���jkK�3SO�n��]��c�-.2�ù5���t6#��6k��NA׶7=�ј�r�;�M�A0ST#��9�=���zs�o*�,_~��j	t�&ǃg0�����3�A�`����Sa5ؤ�Kj�� &��7q��u8!��X���,ei����HH	���Ԇ%വ�!�v�)��"sK��VZd�*�(���U�|�S{~�M]63_Ӥ�e� ��G��ˊ�|�bu��z��1����D��1��L�M�!ajO2;��3-#f'o�L;g��S,y������e�_u�7�'K�<����}��>	*��>�������<�rcg�#PYx�	�}6U���N&Ek@t{V�I��'(�ʴ ��!q�j�jÝD�M��?�g���˺�Ǯ��m'-y�h��"#���%X��F��A`�j�4+� e��<1�\7����ӓ�]G����	�V�2��ոo�Nh�☮�dE�T�4����§i~��x	�?%^fNj�8$c��j�c>ۭ6�o5����H��m��>$���;BN�E=9�ђ�Ŗ2H�d!�з4�e�Q�d����*����}n����`o�����ు�6o4�b,2%r@y�R�/<�/�$�_��3�ޕ�m�R�}�"U �t��?�F�K1o�d7�b�h<3�~�F�WE��(�W�D �g`����%������B@F8$~���6�ex��O�g�c��";A�T�Һ��5~�!r1o�ۈ������-@��iTSd����Ƒy|�ND}Hfi��� %Rׁ�z�h"^(��A�=��N��O�(<%ߍ�8�~��N/���i�P>E�.�������[�[O�i4��^���*�x���'js#ˢ�8x��w����~�I��7]&(<�P�Z������G-	?��{҅͆�g�Od�0�fȄ�.ϦI��[7�
ޠ�̛���m dQ�1S����=d~��*U-�7�9�O���m)/�6$����GDZShszNnE���q��b"��Zb���:��M�.^�J
�ݸ���z�H0���$ky�������x�����c�%�yD����U��۪v�`q������z�_������_������n6�kK�B���]S#�7������C���0pl��S�<��^:ǯ416�YL�6�	e`�f)E x���3e���]a01�P�f�;Ĥ?9o~���S��G��-�Z��ͭ�aS=��LW�ǩU[)�X�`�+ �v@�/�0�y��<W|�H%�l�������RqZK_]oa�f�����`���TdJf~���<� �M٠�Z=� O��Q-�*�?�z�F��}�O�y3�v+u�-V����T1�C�؅?m�zУ�.1�Wq^��do�y#FF���Rt���m�N6��Uz΍�W��&|9����*zxB�ds�-�&ԕ��	]F`����y?�P�����NX�#���Y��0�ѭ5gX�h]~��Z6��!BB��졭LI��v��Yt���L���jvӺ�G�H<���ʤ��m޽"�r�'i뗏������L&�_�<��}�f�u /mo�qE�(�;]����}���}ᾳ��y>ɀxFF}��2&8�O�X�[��ְ�8���m��K����g2�XGk�4:�WE��\YݟÈ1-���Hr��*,H"��'��QP���Us!B�T��"U��y�;�e#�U�aG�Tr�d��#�8�mÚm�߾��k�R!�@�KO�8
5�q1��{�@PHG?�M��39+�ۉId���7MX�J;�ٙL4*������N���/��� 4�KQ8�^��H<���n���=�����0t YcF�N�oo/�D@kF\ͫ��h��A�!E��uCϲ}#X�����?9��a[��=�Qˍ@�^���D&��7
���o����7Sn�o��R�UL�ѣ��Q��2
zm���a4�"���"U�֧�&�����J��9~O|$Sla
���1|}bp�{N�2��TvH�
%��[QC�%_u��-���p^�U� A�u��P�!������,i٪�tz�J1T0�� ���rh���a$t�m�PB5/'��8��B�l�R�T�#�Z��a-C����X��7Y���˛P麂���2N���~���U�٫ s�̻o�`������h`��ӂ��e3��.���6kX�,������Ȕ�\�4��?��
�I�w(�E�W������}��)��gW�q|+�hsoi�S��^�	����l�.���y��̹`׍���s��h=4:������������Jaa��8�-���\��7v����'|���kI
���8���ej��E��Y��?x��X>6
0����q����-�����D>R$"B�E�[���G��te������2�JDV�vR�N��PSa�)5�@yC3s� )�9�.���~M���F�R*%��^py�~�U��|!�
4�M����l�Mܔ��4�� �bو�:+��֡`��L��Ӻz�&7�  �@�^
K���T��<��j����k�4���YL�,���ymg^�Oa3Z�iRþT�oG��S|���tJ�/�3�h����M��1f��N��K[b��Ow�{���Y������v�ٶ��x>[�������R��p7�p�ӽ]�M{>`P��>ڢ���%��L�1��Gf�=_�!s1��b,�a���vM%KsZ0��V�)����,|�j��'M�hmBǕ("�ޖ����,��P��󎢧 :�����xn�m�i	�DI��qs�U�-�*�vr)� dɬ Y%%#��Cߌ�g5��������@�.���1���(;_�q��9ҁ�����4~����7������I�N@)�θ����4��N��*w؀�!�	ߠd�U����	�����r���l$��?�
��1"N�� מI�F��Y`��M=��)io����/�A������e0�QP*����9R�#\p.��'늅s^��,���Q֬"���#�{���1��!�u�T��ˋ������}��ٱشՠ���VG%J@���; D�d�|]0���>��b�YrO��|K�	G��s� *�xX�*	+RP{�Fa*�l��T����J����QE!zR�٬�A=����LT���6��{k��k/�1��Ĉ��?���TS����FY�f��:���[�x���0�Э0E�wv(����U؞˓m�)#��N.0�
����wWQ@��5�/���81��:��m����F���6_����V��S��U�)�*54�E���)
	C��R �~S�Unb�XM�#�s���?��7���J@���#��a�Hp�T��8T����I0���!D�J�CpK�![iұ �@�]t��{�㰮�����)K�b���Vܡ���{��2x5��PBJW����x u�[m�`������#~?b�E�6i��������p1�^.N�\8��/�0�2����gy�3�5l�	eR��?����i�2n<�koh�ғ
�ZHN�
������B��v�^�#�j��$e-�ZI��#��m5G>���ü�O�/�,��U��;�3�/O��9O@C��w�H�G͇~)mvK�-��2C��+�}9P|A�%ȶm*�e{��@p[Ä^��#���-1X�I!�%RַMަ��@04}KL���iW9�a�r͠���� 4�H�@�&8�G�މ����>���ιg�!��aẬf꼽��5�]�NM��o����<���_�w {�8^�1�|�O���ڢ	��D#,i�;�dkō��X7|���>K���qX׼�������MMp]��8���hܭuAC��'	�g��@1(���C�(��*"��=�yO���V�]�n,���I.�K(*ܐ��y!�#vCS݋��
t� �k&�%Õ��I	�f��[������y*�/�D �JjNj��M�j
��o�J	@��HW�x8�2�,큃����@��D"�[^m9�ғ�نKe��x,Y������Y�4�N�� w*�����GWh�Ax^����;�n�r�~�@37k�I���I[+-��+��.9�r�� �Ǘ@Y~�N�|�.hI.N������ɺ�,�vciP�h֡�ֳ�� X����<0V>���ղd�� Z׸�X#��`��4�M�İ<n�E�D.@k�,�.��4���o%����gr�ӊ6��G��˞]$b�5�V��n-4f�Z��N�Q����#9���a��,�"�"#E�!���:.��3f���!�Rd����v������Q��}��1n'NʥY��^��ĕt�H�ٍ��´��=��Ұs@�]�S��-F7 �@0�Vg^�%>%D��b�a^��.�.��Ť�����>_��D=��Q��eCQ�������j�"Χ���>ţ�oC��9nR;.���xn���M�:�-�7�ߺH.�/Ӌ��/��"�=�ڕ�s���h��]�l`�P���[~t.33��~`�R=f6<	l�fg�!�y�f6I��?�8�dBqZ{IY��`BOy���u#��n��{�bb�z(0�ݻ��4�+���(ɾ{�[򃖨<�\x�G�`3�3���o��#�O�1@������#@�T9�K�!*���CC����7]ە\V
OZE(s�M����f��(`s8�W����d�K@{z������_�@]`�l�&Ok�sy4h֒��vua":��)q�h�^-7P3Iщ�
%
l	��AOy�����7hf]�u��f곔6��d�v�V�찿b��\9RᓈǕ���R��bOҀ�w�����=�0�8��m 9,=���� Ϋ��L/����`6Q8�<; V?]�DѺ���1�OQi�lׂ�B5�Qw���ٕz�����C�\�<9l��Z���;�� �$���0g*Om��g�|�FF��l��D��8�� >�3"7����"M)��)
�:S��ZXŞ�:^�k}����`��b��l#��V{����o�}���݄cr肒^�h:i��,J;+��[�:���ne�͈E$I�\��( �>[��V�� �[-����	��d��u�×܉��џ�|�{�̤F=y%�g()�5T�8W�)�Ӕ$�k,����0�����Fn�UP)��!.;t�H'U"M9�'��qE	�6U�h�%�\H����y��>�������G�"?|䰷��?.�TU ��~F��V�tb�e�Z�9� ����>�@�N���/��Wv$����?�(QB�{w�AOX�@��Ip�qþ�f��M���]�>��9_���
�e�!ҏ7�]��#����s�WV@tr��f1@q�2J>��%7J�;x?�sH�m�?&ft�w�X�>%�����2(|p�F2���ޜ�9Nt��/}�\��g:׹b2Q\�\�P�]���SV\w��N��BR\y�Ĭ��\�V�J��3���XŪ�#�q@�����gr�t�;�V�Bd��U�qA�ݱ�B>�m�e�hFG�y.��+L���G��{��1�E����z���׬���S�xS�re�@�/3��9e�`�F��~��������F����
�rF�4unp�J"�=�n2�:�6�^�!C��f~��&FS�����&�^m��Òo�]�QPtx>Z�&
�Ur������g7@��V�_[��ua�{A8VY ��#��tH������=�c�(i/�d����
�}���U,�Ho�C����#��`"+�X��h�}�KkV�c @$"�����@ԑ������/�aJ,�!1r����$}f0���O�����F����<v�]j��W�=�D�UV�䟢8���!�Zݫ�o-W�*�h���W쬤���
��H������,C�h��*r���I������A���d������^�׶�x���o�b{
.�h�I��B��{ ш}s�.���w��\��u�ɝ��ek#847���P�$Ƨ�EA첩9`X�bao�I�Qڀ!5�*��3:z�_���#֒X�m��?��"j1��[��1�]\S����o��W�z���WZ�O��vi����Z�3��t�WIOܣ��Wi�
��I�����&�1l�v��k]���yu��#��p|Vo=4��#��"���R2x�����$b���jK&/!d�α��+���t{I�Y<���1��p1��͘������rZ�j&���Зː�P�ܺ,狆�9&��#�I�4�F'�D/��Tp��~W)_�2���P���1�A�лc���6���2Ϧ,)|<̉<�(f];���7�D���ф�%��4��T�ع�>�X��M�O�27��h����s}M�-�
��-���b���{��1�|��k�WIl+��|4g��zgզD�4�K�.��;���d�K�1T?'�㣡�
�u��\Zj~�2��[��b@C"$%�
���Sn*�;����pt H&P��I�W�;I�S��sV=�2(�� _;�nmxL���P�S}S�mS�Q߽�Ja%	��;&�����8R�J���A���E��I���>�Z��E�k�v�re�L_�;Dt���0Ѵ�f�$g�Nj9�ʝ�4k�t�G�I �,�������Q�Ǧ"���,�f&�QU�:n�����g��4�x���� ��:���Q(�]�u��M�@���>��@uN�w�'&,}ܶh�2��,ۆ�M���hIz���!&7pO+��x��/�JQ��o<�\f�3&����E(�^���Q��+9\D��}���P+yL�����@��Wh_H�:���8]���?�l^�-g>�d�L��J���i�'�a����%+��Q�\�\k�GFR�S3WDV����J�<Z���EW N�w��}T�^bCn���u�%�b������rDҩ��N5�(���#;)�X��߭�ŇרΙ\*'` N��!�[h�".����i\��F����|s�/E?Unʹ�m���Q��s���!Hu���.Zk�.�����"@G=���a��`@��TqcTC���9�>u:�ny�.�3�Y��u��y7M�w�sMc�g�&��3��x��(گ���*Ƶ ��~|x\��s!�V��)�B�0�����(q���{F��0\���b�k�WW]�φK:CI�=���+O���;{�7��â��I���b�T��}�4��M�Ij���H�����.Eb�Y�\�Q�˩��3V�[^�w�AqݤD���������|q3ӨR�̓�ҏ���F��;�c�ހ�����O�l�Gs��0�A��I�����S	#�Kls�F4�yYגE�1�o�?7���[��p.B��+:�Z����7��ZX q�m���{���	��7��.�I��0@(%E�|���V�5�� ��I{���4�_���y#�a9�\8}�CC�����nU�Rs�Ğ%��N'�/O82�h���>�`����z�K;r���<��owu�v���Y�߻ƥ,i��9��wҒ]2�#0�bN�
��_�fFS�N�{%~Ah)��jW��f*���Q����BK�>Ӻ�Z����_��)$���"ȋ&���@�X}�o��88��lg��Ǐ�VT��iHTZ�J<͖Y-]��a�Q��-�Ɂ�H�D�KW%�[2��埳��b���imB�a��B@�X��h���?�v��n;���J/"�@&Mz>`SyJ0*7B"��N&��2�3�}�&������?�	 �B�>���`ga��k�Q��`���Լr�"p3�1�YM�#��� ��<>x�pK�����L�s��� ᵡ�.aRi��^X{h�NnR
�^|DRQ�q!�s�i���RWZ�t`M:.W��m�.ݦ#����)e	�7䙅����|�5-c��H"K��ϸ��F��5V�̚���60�J����"#�=nH�.,^��v��(Ś���2v�V5�a�[�8�r H�ޥI-�Q�C��#��_"C��3U<Z���в���L�+]Խ�a ����:h����\��?�	��&�%�nd���)��y���^s�/9j� �Y��p�`"O���w>�o@^���'/2Yza�����]�9PÇq��#d�7�����>I�6�|�);�Q��`M*�ٗ}�gJ������]fM��7	*�?���W��K{}\&C�$\�R��S'~H�^�H+�J(��Aew
n$���ME �)���S)���]�3;;d�:t|����o�0wc����\{^��d�$�\pc�՝��}RB%�3x��&��➋��(``��,O���O<a;��۵�͕F`�1y1�kAO���C�.���C�N�=�ߊɈ�r��e��,��������݂ �����W	��I�-�؃�S��
�9�4cV��
��KG�h�s�x:��t7�ln �B9���Q�iM��J��A6�K7�%��A^$��}f��J�oZwL���q�R�Z�/w��JzCǄ~��wbO����]��\_������J ӧ}�>���hHCV��&��6j���@l�~[���+4+6����8L����yM�1TW�8�]��pS��h��&�~Ѫ���d�x�u��5�({��؉8� �b���b��A��K9��T
Ӟ�x$�mAkTbv�j�Q�b��h��Etj���;o�ۦ�5��d|K2�s��	X�	����z�d�8R�pT�kG�\An��S��$�e��A�=3n�IXb^�cJ���zFS�x�I��ַ����+Q�ɝW�~&5�|"x�(	����E�Hg�rZ�c��4i7<�^���L;1����k[� |<��_��(c�����s����X"ݬ�%վ�HI ���|�|��f̃k��)�{)
����bo��ig�n��83��5���DիE$[0�R�?F3�bQ�*N�t�?�؟ �����0�|4&�0X##Z=��7 n(���r��x� b��}��~���b�cU����1C��e��_p�2c,n��S�+�H���:gao9�4)����p�~��s��Y�C��[<�S�(Y�i�W-���w�`��L��*2U�������2����֠r@���7��������٘�)6��/e�zjE�/߈7LQ-��Q<R��J��v0���uó�&U��PS�XB�=\Hun�M���AI�-�-�*��N�>vͷ��������S���)��<���o��	����rx43F����f�e�y���!P�b_tX+���'����!A�Cڷ���@���$��]�v��"���؃�~T~�y#�'K�h������ƌ��zľ6t$�J�P[{rm�v'�j�	,�?����਋�(��G�~x�Z����\�=m��'�S����+y0�W�Fђ��j����]��b4<���T?����>���%
_�5<+bZ[�](f�I��+Uyb�`����L�X �v�&DkP WqI&�7��*΁n�w�f�J�����x���x�X
��@2{�����SU���@ۿ1{�.�\�
��.qJ`���J�V��Ag����#�����kp�$��[���}��!�K[��]_o#_R�j�V���n�(ޞ�������I�+��w�#���Z���h�oY^���崾|L�ؤĴ�2ID]ӽ�K����*�>�]V�j^��)�f�:f���އ^%徊�g��u���	�-4lG>���4�e{���n�:#&�,��L�]�gZa3�߸�W�-�ecy���$��I��2�/�FS溊Z�T[�"q�wq+�ˬs��6Q�{y����7��F�8m5H�V
�'�=P��<�@�NI��������N�.�u{v3�~�����ʸ(
,�M�����b��L�����k�L��y�a����_52Q�i��R�!#�u���]pt��ە)2��,*��MY`=jn�W�_R��eAxu�1�ҾG�� �ҫ�������v� +�9���Hv-��-�@u�G�uqc`�%�fe����x?��;�;\�ˎ>�և�<ѶK�^fy҄P�����≵ߜ���H�WZȥ�r��k�V���[�!]�,e-*�K`P��&({�E�����|�3g���\��V\�f7����xnx}���B���	u�;m�"�s�i��p�WSy���;��`��I�$u�q�O�;{����'�"pV�V}36P&��BՁk`%�)��C\`_!�.��*K8�=��Ap���*%@a���AL� /t"������q#5$��
W�#����s��y�5��9�x�G�R�&N��𼆡4m��d&���y��;\���<��BQ��7p�N��і��N��^	��م���$}6�6�n��cH�us�`�L�=۷������ͻc�TH�M�p^�S߿�[T�H)�3�q���Ҝ�Ky(�{j1d��"�re+�Ə:�h��ڵ���}М�����4�\��uW�Q{1Qd�l�;(�0�9�G"I/��X��∭p���F �+CA(��~�G�u<���^ ��:a��G�IY삳�.}!u�k��z��WE��wU�r��)�,�� �5�V�.����aB�G���+�<r+�� _�ΏZ���<�{p�l��=����.1���|����]ϟN~��3j�(���3���z{����Է�m��+n��A��FL��_��i��l��&}�:�x��>��b6,z̀2ݵ6~>Ar.7����N]p���뺱��G�&;��9t���v�b�o'�5!_{�.�)A逐��l�-�������A��:�$���&��D��m:��2d����M���k�i���VV�Oo��D٘�
�`7�rUs\���%/Eݻ������kD����W�� S�X���_j�uw䅝��^O0����#��J�R�K�h�҉/�*�@�+�=��9��Q߾u��7O`T�T���v�*͓��/��3�I+,���^x�iH6�P\�w�v9S�zv���#���Ss�֊�{������0�4�8Z��0�:��hTRK@7��I��3�o|��f��U�˂��&�v�3�,��I*vUd�Dm�CuS[�)��
��{�,��&!����ֳs㫙=q��E����&���܉�n�|����(�/�����+%�X�]|%�W��ݬw#4��'��,W�+�vt�j`�h��p�n���ռ���ac���W�#�q�5�y�|M��'쑜&/�\q�3�D�K�6p,��^�"���%D.�R�hE��� !��Gڛ�(
LZ�!ω��@��ի^տ�Q��(KEt�Zt�OT�x�^ZEڳb7�f]gBK.	&,d�"�4?�mh�=_�y��A}�h�%+�0�7��' �o�Qc���2Lhr�_��8g����C�y�����a~�������*���%m�!�ۀ�x0�E���KZTN%��Nҽ+�G�Fq�DX�xp�t j�^����'WZ�qe���'sE��::�[�O���P�Pb��r�fb� X!���~�>��M�,�)��&�5b�t����z>W�#!|���B=��`e�P�C9������Wjn���9�����2�]j���e悯�P���N��dJv�LOf�\Jp����B�����f�i7���Y�>�j�t�� ��Ͼ� ��O�ºh��'��Z���R*q~S��>=ٜz-i~�Z����Lf��"I}t�.�����}��AN;�Z?���J
{�aD��+'�xE��$tQNw��F��|~���84�#|��A�ˢ�y�vN����8�$lK!��HNҼ 0��Q4M�[r��4�u�Ō��*��R�'�*b�]�Ң�=g�ٻo==M�k�R�>z�H�ٹN'��֝�R,I�6�	u/1#��7�fu��K�~�R��>���v��08�
r$���B�M��u����$B������8#��2?�t7�ѐ]�q�2�,�sh5��e:�����&�Pm�����] 6$-n�$M�@>�ٱ�Rb��W��l����P.�U-��с_ł#yQ6w0݇k� m��O9�!��@IF4�Lg~�k�9�^z�i(����<��Thw��b���K4̌-�G����#�+�/��v�I����n$s}"t%��7��u�]t/�0?�j�0�&�('�'�!���_�|�l�1éB�rn�A֞���4x��D����������H��y\V�l�9ȿ#�KLS#U�ۜ�å�fa�yJB	;R���,�
��Ŋj�,K��q�̧�a�{�"�;��f(��+m���UX�Nv��L�Cp`e2�����z��V��`�İ<M����\4���lc���m�wmh�C�ʏh\���4ZZ�"{ӎ�R�Os;
5�:⿊���6��+z�"��MWR�HP�>C�X)��ʐ�U�8��4`Y�Z$ȹm!�U��"'����Y65�v��T�n͐y�Q&Ҿ%���!���e�{S�h�g�^����ɾ�~t�V�d���9჻���Hܝ��ߡuw��7[G��M�n���"��(/ Q2�F���k닏������ysxD�%Z$jY�
��V�_�`� �KHs?E� �{�����q+�L&5+p��7�ۇ���	�O��s�g��Qc���+k;d������u��k�n�.T���ߦ���ڒ��l���А�����R�����]��찁��='0n�lA����,�]��5[�|w�5--[(Z-C���M���\m+ &l�dQ!�zJK}
�T8}0b�@�s
�����m����{W�'OvDD�����"���	 X���M�o��R<u4��w~��mJh���`��Q�8�Z&���4�ӷ}��/�/̆������,$�k��質��<%x���
� .,w8�������Em���G�檹���&�"	���!�X�W��a��{�01�x7�*ͽy�|x��^>mD]�@`c��^�"�8ь�����,��N/�Ƀ����$~_���G�ٕ�_MR��qܩ\R@us7��߁ʀUsc��$��F-���pC*	��bk���A<S�P��d����ˬ24o�SR��B�[%�h��N�~\��ٹ���2r7���!�V���5<�H�z��=?Q	��o�����*d�9n�Z�lI�1�=Q���Xa�ϑ͇ǆޞ��A��-1�ifj�����&;��h�xm �9�T�Ie�!�A��5�Ƀ�a~���ӭS��0�Xd��D] ��jox�L���"��`K<G�BjB���ˑ��T�e��҄MDL%�s8K��8�"���-�	���[�+P�+	�{�,�l.zs���܍Fi(����)c8�����Z�>������~��&T��q~UV���
�t(�fWF��C2�d�����1�ŷ��|�C�����q|�ʁIz�/@�J��r21��)�H�c�
O�a`w�Ro���N,��r@��` R� &��\|}��p��^J���S����tZ��U��]�yuo��±���~�"��]�˶��P?K;���C��^�vtp]���\����R~C*Ժ؞���2~�d{�B1�ۖ��@7!S��4r���������E/5u7Q&
 j��`����
�ޞ�h6%-*:%x�HN�+���
u�IȲ�|�fx����O��`��KS�c��)r���30���"V� �*%�Cr��y���:L��e}-?�)ײ����cy�Y���������ĪƉ���:v|��n�TƇ�� ��U0p"�!0�	�7�ɥ������+g�b��`����z���4�F_!���d �g��Z�jr0�ML!i��эP��x �!lP�����f��:�;�o��9�s��_���om.%r�ܯ���s@��C!Z�3���:�F��Y �#95u�o�� nY^��5�{<���L}^��������J���$��x˛���tOg��	(H6�@��T7��;�����>�����4`C�����HH�咔n�V��zx�Z����*����xn�F�d B/H������o�����~��6yD�<����g��>�(ԙ�E�2�!e�}��O��+�䜣t���md�_��1a峈\��q��Җ�2����cJP6�6ǋux��%9�8s�+����M��wB&�H�N��li8F�MP'׀�6�L�{MܽGh�����7`�6I�&9�����2��(��u���ԇ��7�f\ԍ�qV��]2��R�$��a:��!�I��������ܩ��x�8�������^X'��xN�7��O?��z%3}�(��c��3@��L��A�Z������M��@En���L�ta��wl�	0�T��T'D]�ϖ���^��7єҧ玬��P3CXz+g�P����>�WQ�~6�ǀ���Gi߂:�Z.��]a�Pd�X<%� ��c1.��tdP��s壆s�$DRp;J�o��U "|,���5�WeM�* �D&\�vt�����Ñ�K�{O��Pß�v�����YEh �-p��oTP:�����ZEY9㫟��^ռ��|�R�IO+�R�nuF 1?�"wѾ����S V�=V��bz>���t̆�������ݦ���n3w��C<ԣpwe*ȬC�,(��5M��E�H��4�9�@�N���Q)���j��j��U}��[r�����C�v�D �c"i��Z�ŏ��JV�����.�\Ҍ1�N��-q�D|�x=���kZ��we*$��
1@G����|�b傪!�<89�ʊ��V��J�_Qd�v��X^9��D�L�������>A$��
C<ܛ�! 3$�HN�϶G@�����n
�a��_΄Ϫ;#�oGL�=�c�Z�r�eNlFD�&l�I�D,�1"ʹ�-pom:i��Ò����OlƲ�vV�-����4��s2�'��򘞒�i�3p(س���k!U �����sv��n�Q�">}3턪���)�-9%��?h���26Ο�%�z��_�qp=:��lwz)>��o�Æ�DE%SK�Y7���M�x�c1[��o��h#w�2ɤg�`#��@�y[ܻʨH\�!�k<g��AS�1`��}qT����2���D��R��QW�[��ϲ~�S����p��/�z��B5RB�[�^#�0�*m�,+O�r��;��݂�}J2#ǵI�NZm� �x��Zא�煋0�k��w�Hivt#A�u��(yfp��:Ë0�WE>�]E����D�J��N�a�%�ŀI����aڴ�cޕO�gc�jU�Ɲ��_-�b$j�S'�b�KInҁd'֔���|���q�ԃ�z����~B��*3N�7����Ӌ�2[�$�/��^.�"����I��o�k1p�Uc��{�[�-Ǯ6�S)�T$L�5m���E3܆X�*,�B����^D�z|��B�X���S��X����NcW�q9�zʽ=�2�uR��pW;|Y>�5XP&��^��yG�y{O_ի
 �5BW��Q�?��p='ʓ� ���)��Ev�����F:�鋙5J�y�f�*s�ͨ� �(��|���M�"�>�y��`	�����[�d>
e�ςt�?��DI�	����*�;��ZE�j�����Cl�;��[�%Z���)��9�'�����s��jpE�����<���a��O�|�w�$���W��g�����MS����v�sK��$�LT�����;<G&��!ڞ\�$۴��Pa6�3%�0�i.X�����v�"�T�f�>8����'�F�V"(��Ka�&�H�~'�����������0�Cm�]㖻�kN�r^Àf�*b�/@� �O]J%X�@Y<�9;Pe�'9g4W���A�S��2�kwpn��� -��k�)��O[�Ӣ�W5k�h8�䤷��d�{8��,'���S��;���,���."O�h�Y�yF��]�;����ό�F�kP��
,�kvV��nB;�[bP�8�Bh�T�\�� J���*�Ê �^u��A��������=����%���^�dD���̰�O����P�ko����ȩ�*u��{�BQ�2䷲|���p��|&�7�xK��/��9��s����P�t��q��8Ֆ�����Γ�ѐEGM?;�U�p]�{�o�^�TS�z�P�����y������ڡ[���������A�pYow@����w��:v5�,̍(���K�z�/i�C$�<�γX5�L�V�2s7���`�ENc�'���X1u{Ѝ�p��3�1ֆ�?A��)��-����>�Mjt��d(��K���V��n���$y2�N���N.}��x�D��H�(g�������+�����[�R}>q����MV����B����c�5��C�fH�����{�Aw>��>�(����0=�K�y�]s#�Ժ>V9C(|��C�*�:�0�)}띈�a)�c/U� ��.�򏴧��,�z����r�:�ݪ��v�8}���#5�
�`*�hu0�y,qM`��mB�o�e��q�;*�nw�,m��&w���r���L"�=�ʑ�r;�7��#Ӗ�^!�C1�&�.��k���AG9D��I����5[p���.':�p�����X���ZX\���a�Y`�R��7�ٮ���H`�lq���߼a��{�vjk;�S��څc�k�O��x��Z�A�ԁe�����g�,@E�o����s�@p�	�T밇ͻń�,��ğCh���������?��u�����5���S����l��[���)Fd*2�GB@���ֽ����OJ�x=��F��n��Te\6�}��^M��o�gW�^H��[A���̌kߎH��%����o�X�/�^�j����,����s�v���(�V�>;�.t}���KZ�X�oB^��%�q
����1��A=��#��u��k��uEd �Y�'� ~��O	�j����^�	PՒl0� ��T� ��4fR>hf%����V�h��l���2�92M�pk������:_B�_^=�*t��`sϛ��o�{S��	�L�.�6ʕ����]�@��c�k�>�&p���rV�C~�#�m\NG�|!�X�����An������G�f'-�|H�YJ�0�%&Ց���O�Fp듔c�Y}]_v��5�K}�p�tE�{��
�9�ha��@��O����kMHތ���Ǌ��Ғi)J��X2brW��ԣ��}%q���@��r�&��ԕ��0��)�WSЃ:t͎�!�~��P�ih�e ����\�ٶʯ���$S|�T�yRE-t0t&�-��v�jMX	|e�/@�e<�Iu۩F<T�JbD�Z�L���yε�z�{qs�E��"�DCo�)��z�Ԗ�|s��~��������	�a�K��yV|`tA�I(-f|�r6����8,�`��Y�,��`�ɓ�R�r��_�^%����9��?����R��Q2�	Su�6�>Q����ud�V�����)�`�s�\R<cVۖ�J�O)%�k=+%�A9K#�\:Qroؗqح+:jyy�ꊚ�M���_���[ؽm�*����5<��"_�,���;T"�o�KH�5�%�1d���}���Ĥ*qmVQd¦/��Z	�W��}�%�Z�7*<�FL��璜 �G����霕�c���[��ƙ���b��雯! �ΰP͋*�I3���5foY<�̚=+�`5d����!jLI]�$DT6�����o�J�!��wo�³Q`d�������H��*J�N粴��^���M ��m�]M�y�"��}���U#���7����9IG�4>��<d��<�?��7�3N}|��+A׋X�"�aVc�i���r�j/��g�&��� �ӆ�2̡3Uە�Y�'\�p�Y~���lx@�g wT�w�r�u�Y '�-�~D��$p�H�)��ܛ���v 2Ι}/�������Lw��,7��Э�S)����f�sG��0I�h�C�uD�wБ�����y�h��u~`@�eO����p��ӂ=��|a�)(c a 0��;��[��J�4忡�˺K
�����[��A�Rʜ�n���+AYK(D�������t�q���@;���rd�̪]4�ˋ6��O�r��12Ѡ�44��d jc���^2�I5�5�4l	�_8��W��ڜqG��>���=����Pul1��(j�BPP~qjN��Ҵ��S�JJ>�0|J��.$j���m���g�!5��.ȑ��|O��3P0�Q
������d�SJ�Y�]}��E�]�p	[3r(]n�GHA%�%�슳���Z��J��l�������y�,�����t��~��7�|R����l�D\��as�}�� �R�����4��d`�<}�nǝ;Dᠩ�`�ڐB�q���z�#��0NE�� �a_�ɩ]��1"1�Iw�(K�t^����$qi �x�\�����/������˜_nP	�тD��(�z��_d��w@�{C0��������l_�.�g�RU����^LB�3��9(���גxj�2���دմj'�-�����f]�2��^��wj(���o
j8K�1�`07d��Ћ�̱@=�n�{Dy2���{����o�G'wH`�C�8TP�:��K��C�l�?E0�A�L� b���m���1��a�K�,������E��~�.{7��:wϟԼp�F��0<�t҅z�����k��<wx�{�� �s\���;���B�{��y�v�BПDOx�UCz����M�3QƷ�8O�RGx��h3�x �Z�n�����Q���BG�_�&������u\ΥXn:%��������ݚx�i��w	���ˡ2#m���rTO�v��B���f��r!�R���ލ
�8�0�����4"ђ