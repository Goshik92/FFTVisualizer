��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]������]�g�� }=�G�b��LU���k��݃�`w�V �L�q6������mk�zA@�%�K;�M�g��N"��Ȑ��a���R�r��:ĭ#��W�ݿdÏ��]>��S ������'���|Ti��ئ�m��Ж��f�@L���{Լ�uu�!�kn��A�s�n~�:� �_v� J)�h��1"�?�N���l��inx�Faq�}T{Kn��a�9 �H`�ї�5Y�!h\�!g��-)�"��(%��w��vR�	�T4���i��`Jb��ϼ�]��Ok����i�$ZD��y�].�pCgﶚx`����k�,dŪ��l�L�~�_�׉�x�7�I.�}����?�t�)|�A���9�J��V�y��a�ooomp�@�|eu�v���qu:���L��<�tֹ���\F=Я���Q#���aQ�D/"/X
8�-+�g�Od:�G�x�6H��J���X�u��@7��1�	���%��\Q���xol8�Q���
{"�$I�'Gxq��R�i*/{�S�����ƖZ�̝�tU/w%���O��{�?��R�X>c����+���r�z���|܀��jG��]+�j S����'+��i-]��3�����.�Wn?�m�<�kW�w����lB�eu|UϞء]5����&l���4�mcsO�jŪ-�Dj�1�zAQ��x��5L�3���n���gO&%�k�Vc$I*���'�ec<0`=&�8Vi�U�D�Chϕ�y
K[��#�U`��Ϫ���S�r+d��F��t�*?�����@��R�?
ӆ��?�/@v���mHg�'��`,yRy����$l�:I��y�k��ot6yB���An-�rd��Sj�<`�k�w�0�n�]2*�����[
´�r���-:0}3X�w����y��"��Eta�w.��P����{�i�hm5��&7�m�-��YN�8�
5����̞��?M�F@w�Y>��TК��i&8�������k�P��T�_�խ��h�!s/�&�I���ƭ7�����[3������-g`��#㐳���3�d�կ�&ٰ���v`�O/��hr�<HY�ݞ��L}6m� ��/qq suS/M�<�J���d�G$m`�1�Q�	�fQ�9��g��j2{��# ^�+D��E�~7�ލ��l.�t��w�������q��u ��j��̊���~;@=��;w�C�����j��4��śP{�(Z��ě`�Z��m�8d�*F�Vٴ���M|"e����ٌ'�\���]���a���i�	��R��9[D\>u[˲0������Q;KË���a<|����gzg�Y�;B���fQ�߶Ĉ�4#mrq�L�cNr@+�kr3ɞ(����3eLT�8��"�Q�7�H�(4�ײΘ:Q�9�B��.������Q�St�Q��JdΚ�a��mh�g,'�N����g6��<	�3��{W���j5T^���;��Q��o}��.��rd�<#�A�[�+��OG���=����SJվ��Ik�'~-%�.�~$���@e��F���}�[T}/n S?+�|���s}��l)��Ɨ5i%��e�?��p�,�",����N�p&ۜ�v��Ÿ�Q`��q�}��J�F��
���͉�ڼ��q�5����j_Rl�r��S�i�F\��k�\k1��CdN]�����d2���idgdrz�-�&y�te�Z�Z�Q�s�][������� {��Ka	$x������ct�{E���V�,>v{�JS��	t����S!�Ze�g�� 1��7���e�G����U�R'��|�2K�
�x�Iq"��U��G�hhھA3�J	l'�2���'���ܲnGu��A���_ ����Y���ӢʼݓZ��`��	�&o'x�L���OCO����E����j��8	<W^��r��B0�x,k�*zE���E~R���6΁��J��f*�~?��C��t��	;�O�Ѝ�(�BNHM�I�;����������̿����K�L���$'MYP��!Z	Ȁ�Fu� �����a�.�tƭ���D�J�+�ixvI���C������%���/U��cK�t�� %��ASh�,���a x��[�z��)�'
j�m��HN�M���a<���������Zs�i#Ya�0�t}��"�s��G��љX��
�� �T^��� ��>�����r����	��x 6�A<��>��iw��Z�z&G.�s��/�D��P�II��sEp�2�$uY)|\{n�
�����k�࠺%�K�]��>��oR�J�
��a�)�/K~�l񭵣�'��6oS��;�*�Q�L	�\A� vw⨈�����fy�'<r�<<{�M�3�Hka�JK�$��%��z{w���L���)`�L����0���#�/��
�́V�;�3��=U�����&�x�T���-�s�uM Rwn�ׂ�\�]M�Z���`��D��T�����Rnb�q�lo���c�bB#ֺ��P`I����"���#��E���Z��� ���˛Lb)h-��(=�Is�N�k�{l��kV.�k�8��o̯Oj���~�~���"�)���]�`Ά<����Yqk��?*�
"���QzW���*���Xc��)ٰl�:��yO�{�+�y�ݧUC[Hqf����������A?W��/�u��^�h�,��ӸD15�
Tl]`�]�z*���ׄ Ll	?�8X�F�_8�+u�Ȣ�o .D��d��`�,�^���E_p�UXb��M'C0�Q�e����=v�8�؆���?7���[�
�K��t�#��Be�/c�zX����P@�q�Ɖ��B�5a��n�|��l�
̨�R��C���nǯ��������GN_��j�7-)��ޥ���X�ڹB��O�2���O?����$Y���[�!T� c�=CXey�j�k����ƞ�X5�\`<�j��͢dV����L�E�u��W�.
a+o��s��<m �����'k�&��z2�v7|����,��[+Hkdҩ@���]��΁s�ݝ;";�Z_(G�,;���[�ŝ��T��٧�]���>3Gzŧ� �ęXۑ��E{P��-���a�I�#	>��b�g]����~C�����zA��B�YŘ�TE�]��I�y���N{��t#R��0�f�R�e	�I]�9te+9��kU!�6֎p�y��(��z
O��G��A�fX�6�X&���>Lw���N�~���og@ȩ�Bz�N]���bN@դ@�<���R���-���q�$C�����ߍV����ۂh��qa�cv���A��ǑOK����˪2�u��-�s��4�a�)3#5�i̘[���8n�/ET�9�G��b��y�\���׻�Da�[;��������ݴ_�?�Y|b�8"
⹱}��ĝ��a���f��S3�.�+\���2�c�`�c��n���Q[���)FD�N�?E��m��ΰ�*�3Wͺ���&�z�-���=��~��Z�����? ��8S^
��[}��]cvC���1�����VI�hZ�m���8�M�u��d�<[��������QP-�6�r5��T�z�	�]���T�8q�5֙�ܴ�@>��!�/�!��w�n{���W��V^�p��1Q��!�>P^DD���ܹK5&�z�Da�[���b;�x���-�O��/k��n"��t���;��pu4�}���#�d�M�1���.r ����}f�	,e�d��'�_R*�:ɳ.-1���A7��𰮔T�S���S� �Y����������o��U��zgKR�?�@���V��ʣ�b���x�@s��d3��oؖ�}:����~N��f��F��;�[�'}h�[Oi�N6��Oƚ#��B.[u�Z��4�|����o"�-<7�b����:X��=����Hl����vԁ�I¿*ԙ�Bz�@۬ϧ1x�Y�zG����`V�^w�f匜Nm�cg�t���6�/P�[��ջ ��'�KQ}I�6�O�&��i �V��':�@]"��$��)���>��N��Z�MK�������u�l��DN KM2����9D�إ� }�G��P���l ��li�UV[Ǽߊ,��h���\���u���@͓���1��X/W�R�@��[ڙT�8qѩ�<B����J��khAC������=�)�������@M��Ǌ�Hp����&�	�:�>\��d'D��V_(����bR5��|Ի�Ӫ|���d���o��d@w}ʡ/��o����jR\Ku����7�b����lL������0G�b��!K�.u�36,�=̚P�E����Fr���)�3q����W#<Q�Ki����u����A:�Ḁ����=�k�B�������DD��	�KM
u#b��JM�WP���w�6�g��7��|^ޮ�pﺚ-��bvD�ӿ�H�S?�|��|AD8ּn�}��GXN���@a��`�V�3_�M;*�MW�_Uݣ�]k�7��:���5�r��-�@-g3k.#c;�0���h'�??�Q����z u.��mC�A�?by�%Y�⮐,�`�К?��~7�1��^-%NX��ցno�0
�`��vaL�߃�&�P�S�@��L���Bs��`E�s|�����KE|蟳W����Ёo ���/x,`�bU0�-���V*���J���w"`k�Ĥ�:卦y�*��biA������!ӡUV�lə�U�7����0\���%���ag?"i�m���i���z)c�\`S��*,�`*�w��{��S˜p�X��IQ�}46` C��>��i���M����5������`1�6��9�Q�a����	o��8�vŐxoX�"��I-�t��t�㨥������;ky�^e&%:��6���n̆���C��o��PGB���<:loR73ڬ�W�{�#[Gi��I�]��"j9��J	�Ng}1mD���ǫBu�*����g��F���3}�(��[J�i��g(�rsѰʬȰ
s#��%h�Q��B]�eҷE�j�,�'h�;������f�00\�������9'����*-T�)��B5��l��o������enŒRa�&U�X�)�A�eNl�^޷'jD5�=(������T|�PT����r� ���V1<V�8����SDM�XRm�"���#������u��.i��� F���~�����E? Y|����z�����q]�������@�g��..�S`-�(�Q� �A�����#[48�P�~:�l�[���|rr�<����]'h`L���dF��tPF�+$(�E�=����^��;�9G���� ��u�犀��O��_�jz�>�`��r���ef-a]iXN�G��_'���:$�_\��y9 rE{�Z��&.Fx���N�!D4;.`���o��/�I���_����o��]J-S�Q�2#M�}�"�NۉsXNW�L`�K_&3$��SV��No�/�T�
 ��j�]��)]O[ݥ�1����t]�)c>�	mr�jcOf��sj ��}�Fk�\��;�8i���~Fz��s�� �]�o���Ҽn�}�s/j�>�[��*����r�d����$��|2�h��o��d`�Nl�~�HK.la���h�����3�05�/�2x]����W]F�H��J�R{��M���ΐ.iz�NX�; o��xN�P8'z�E����
����l������|��oMGI��BD�{#qVY{��"r �\�{��%�U1��^��%&�����45`��S����31�g�"�9�l8�.B�K��9����P%�F�8�y#7� t�����Ʒڻ�X�/��
s.f����s
�;����0i*���§=�N�8-n����8��;:�q��u="�dw��#y͇V�ZWɞ\d��2�-S�@#K�?�3�(�!xZ�L�F���`f�˰hC_0d3<��;F�5�g��J.&���&�p~������"l�kEVٺ�7��+=
�2�MU�}�/Y��&�v|R��hܧ��Y��]M�e�I�����z)���F���H)�� 4>z4μkyr�4C$��b��J���k��r���㡙s5�m[S��1Ad?E�?#J�?��ݧ�f!��M�X2��9
�
h�ԝ����*V}���B�oF)�D�Ǔ{{�,�z�)u����XRx�9����?����~+��#X��rʌ��z��;8gx,�w2���i��uBc�;!뻨��tQƎܹ��$�×�a���Vs4fc�:�Z�lqy���<yz��
Y�곖0V6����+Q$� 9�vkD��cj����"H%�텚er�
0���R��v��5˨�����w�?d�JV���F��&W�%�<���A����[K[�A3~�uY���(v�me����������)Y̶	�P�P��y�BC�j����9J�%�8R��{�:�~&����#n�^���b�Hߗ�>�v!��В+7V���l}y��7M���K��<���@��z�A�٨���Ʀ˔��(�A�c%7S8ZQSo���"��Sw�]QceV�Fy�Ƨ�\y�u�.�@������䥞�������G|ZdR�>��_| ��$�t��f'��k��ޙ���{�' ��v?���ZD��Γ�5*���7m}b�_�3t>g��5,�@�ʂ9���b����?��0��Q��K�ъRI�S@��\��2�xB[����%);���� !鈨���_��`�$���;�{�ܘvx� Y����k�}�=hiezq¯FE����Z4�9���zctCY?�*�_����\�q�D����64�_#%�.��Mju��>�ѓ/��<�|�T��4����+�N�c:@K�uT�,�-�3�~���|�2�dٗ�س�M�2/77�L����H')D�4oQ�<���LL���Lޝ"��J��"�-:�.���o��tk�dg���(�]sy�03���	=�Q�Y�4�����K��Ƞ��s��?�h���ߣ]�����V@�i��V3�둙�G%�Swc��Lh��C���I��af�0d�"�g���q0������\��"�d_a�!:[kUʶP�59�.}i8#eu;�;���䙄�`����2d3�/BB����<$��"\����7R��eQ�x�*'��!t&/�$� wr���-z�]v�26s�Z+�����,�(���1���J�^��p�i�B[4����iT_[��w��U� płyR'M��������k	/p��E���9zac~?I�A�r�W���)��T(����0�o�y+��=v0$����)ù1�`O�b �Q'����s���k���k����'�H�h�c�f"{(٤�eX�M2ͧ����g����BwfƓ�Tm�ǒo�!_���!���/�{�zx�a���]������W��N�"6i�{��l�(�S��P$���]�X\��C�r��8��$襡�|�jNû�*�-��Rͬ��j�"�-|S�%�E��S�z~�ڙ��A�g��9շ�#m���c�mJ�|
9�6~̵>��/���N���9��.ŨΘ����]J2§@�Y��5���I,�_�ˁ���cK���`+"K;��Ꝅ�
�=����K6�*�z_�r�K�ˑ����Z}�$o�F��Aj��Fa6i��h��T�s8i�­=ZN�ųK���[�Y�q���� X�R�Wb�(J/������g�e���,����7��������`B3�tNb�.M�;9_�PF\1�<�b
�*� ��Z�oH���ӯs
�H{�t��'��������fR]�S���1�T[p�[�n�Ю��{I���1�sV/ѻV�T\dy�Le�S�����t]&��;G���5}�exj*+�T+Y����=5����;~#~ /)��C�?�s�i@�Z�GV����d�7�il���Ѓ.*�\�R��+Q��A�|y�;���꘩A�d��tG��Z���o!���"!p�^ߪ6�8=2�1X�v:6�Uc�|
�ꏨ*�d��S��]�{Fj}�@�#��~hy��C�P�p��a�:����w+����7	xWOݦ8�Z�
5���������x��q�ϰγ�2�����N��Et���	d���Q��0p��
�C�^��x�s��_sU�WCਪ
�/�"�����gr�+�2����#U��ZH�(M��U)٭Y�~�a�p���%��$����Y$(�!dNY�_���Ψ����h�k���Ra��T�0�:��јK���������Z$᜻p�w��7ЕF��-Bg�Gs�Y��u��	���y����B���S�2����0']����! �m�[_�Y©�{������B�I��t`Lo���[��ܲX1a*���d����<@�3̫K��!vn	�7�7"�q�����>"<�z���}���5VJ-b%d�!0�4ɀ���VLbY�݃\�9�fx�c�� 
�:��q+�#K���n�="p����̆�}�k��:�����z�� �Wr_��
�uZV���4�gۋp�sȎn�VLz�}���9gF�1�a�b�DWZ'?4��R4�I82g���J=r�X:L�w􋢫-ӈh˵��t��e\�S��xN�~��� Fn_�M>�OkK�V�,�hH~Qʅ�۟���$�j)�����w�+	��T�k?�s!S