��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|�&���ڴzk^�2�.��ܗ��"Ä\�e�E{��#�B����+�8�~z����.৫I��e�SM�,���}8��	\���wJ�jp��L8f��͓*ܡ��X&�hqW1-a|��^�q' /ڻ�<fA�SG9��d4�*��;��\�2���?��cL	�,x�~��W��zm.��p~�``�wT���pVgx��OQ�J����&J��l=��e����O�����Cu-H		��M�ęF$%�o͕��$RD�Ƽ�������>_2)�Uސ9���O}��=��0	�r��,�� @8<v���Җ�=P+�ӏq�(�m��| fa�9�T��X�d��4P�ϩWh��%�ʎ��;�@���g%WS�8q�Z��ї����#�����F&�!ޣO|��J�ۏ�ǚ*��Ά���8��@II�&=���JpL�wKyw�#/1��F6B����EldK�?�����yUk��F��������8��N��bP|z��zg�$��^�'z+�I�r��G;9��2�["{�q�ZUA{���*�;�ӌ�I������^�M�iu|� ����ӿ��ְ��{N��:�"�o{�*#8;[Ü2O&��ӟ`%�:ϹtUi��~"G�e~��M�������o��x\��!��&)�%y��c��6�V�A��IR��ڰ��¿���NTfH�;��%�/0�XZ) �b�) ���Z7�����X¾�<e��Ag�f��A��q��u��R���uW}P��1�B�H���9B�G�y㐣��%���Ig
"[n�|�^��7E$�Ii��䷦�#?��8����Hh�-�0n��+� ��q}�����a<E��$�x�^��-pŕ��\8e��j0U��q�
�X��I��{`Q@�TT>'�p��K`���Xy���U��k`�4N�1��Mmj7��i��k��:C��:�)pB�=*�[��jC��TL�/�l���W�-h�vz��cl����K��bL��v�܀9�y�T~��j�CEM�cTk)��)6�Q�����q/6�+��&�C0�dIe���,����_(ʳ�X���WËj�������	C=��l�&$�x*rS�@Za�9��_�0i#3�PTD~F������Q��D�����ە�����n(C��vD4;����񻘅o#���|�%�$�zF�/N;���<�u?� @�.����pT���T����-�{]t����Xݤv�V���z��N~0P:�OI�f�}��p���r�h��pC���h�;:*9�����Qzt�ߗ�L�-���!?���(�eS�o��B� /��L����<�����g���#99����m7�}ǃ��07<�?�3?�i��=�ѹ"p��M�scS^��XOՈ��4m8_�u�o1�K9�a�#��	~�˸����7��{7��L��J$:�0�:����V�d�sm��q �#{�[��	-�R�nC9��A�iL�҈}e�q��%C�5q��6𚞾����$��+��Lba�f%dU
�n5�l�W�9�H��4o��Q���S���C��@�rc4����@�	��$��&�G��#k�g�=�F?T݋w��czͫɱ����7����Y䩋�������O���r��,��N�������*��=��\	'&��M�Yg���O�b�Y�i��~���Br��H:���<͠ �����
�H�HX��>�'��;Ѭ����Ҡ{YK�o��.�%�L��UB� )Ax�b�J�iÍ</0��`�Rr���|O�:XA=������	Z��p��(K�s#4�{���gp��9#!�H��_���:%��o@��������T�zc�ʂwfu?9���iշ�c�~B��[ �>�vf��.v���4O �_
�Y�qJ�r|�\%7A�m�h���վ-.��$(���=$&�$�s����-1�u�UE�28�=��Q��9��<��;�!�ōJ�C]ǥY�ĩ���'��g+K���7��� ���JD~�
t?�+v�7���ඔ��Я��u�� t�i@a�������M �������_
�;P4�@w���+��G�ƣ�b��]�
<�*~��(�.>�4�!�a�Ʀ��c�?���>�2F�\�6���e�_�Σ�F%�,O�
3�+;��&&}�D�Jb`��
'��g���.96㌗������Q=� Z����_5g0;�bO�s�Z�(�oϧO�� �K�2��Z���7��\B�C�F�Nz͠GU��Q����S�Ρ�?��@0�vFQ)��a���V�K�BVP��b�E�w�'>{��S�>2�ĮxX*�L����}�X�\�c��D��!��Q���M�U���~NR�++~�dAn/춣l6|�e�aX.ü�l
W@���h+���q~ݕ�ӈ�K!�y�j{(�O�B�{���v
KT���Y��z�y�ٝ�D]�J=E7���C�-�	�Q�<q��a���.L9?��ο
��r"�xYlF��9w�� �	��zQU�U�� �%�I�/v=x����臥�f��w+NuNV��Z�i|?�k^ƒ���?3��F*��.ڥ҂�Ó�+D5$��@����be���l���dQ�EgJ�vQ��X�/#���^�C�<xc	^~�ה�춍e:���/���|��!�*q&A�8�4! �:�ܹg��I��|��|G�����5C9�(���l,u0��8���,p}�ȋ@��{A�����������8�YpkH�quy?��z��zo�x�@��ڀ���-�xSr!�H�#2�'�LT ��<$�*`=$d����l�Y��;�^P%��=����&8��t����3��zΫ���i���)5��j��=����L�F������Z�!��W�7?�j���e�U�H�'Ϧ5�0}�L*�I͐�Q���N��S!��Ų����&�}��'Xf��df�C(���]�@�p��Ԫ���������)� ��]*��Ș�f�-�E����>F��Q����׎;;�)�����*ǒǗ��\���і��@��F�T>0���̴��0C�z�E��t}����1ԛ�v��%�PGy��rL.��a	��u��Wؠ�kX3^_|q�q���w[���5�,�ai/�0߾M�ҹ�hj!6��Y�,��)��di�X��(9?+�x�"�E��`�،�W�1�������Ss&R�<��iw]4@Pd���tN�ڑ[���y��<%�E��Z���0���ExA7�tT���O�77�A��6Wʂuf���꧿��~	�1c�� z����W�O��~Aw��9欒�ƹ����Y�ླྀ�H�	zB0�:�r��(|���
F��_�n9�Ķ����l3�N��v�C*`h� \��үRQ#%���,K�8@0UƯ�O)K6�<%�9��Iڝ��$�C��2���G}�m���x�F�c�~��,�bWz}�h�9C��Z4c"a%��\C=[*�nNT+�.ӂ�v��
�>�ﶆ��8�����H�y9�8x�C���-��������h/�W�p�ۏ�M��e�Z�Ô�3AGssm#�[�� �/�q�M�|�Jy9�1pɚiȾ(��Y�D����-Q[�S)h} ^'O����`��A��X�?l��Dr��P��i�|Z�$ڗֱ4�	 sz�����P����!�of�6��K���*a��>�p�E��u��&OεW5>�p�Ej��+�񷦓#XZ�:?�p�[�6����47#ޓ���}�DO�� �^X�k�2�/�U;wy�hm!G�~���S.Sl��9��tk��G��ъ�hM�$�7�ue?�����W^a�<���*�>d)QS`9��?	�F�x����qB1�a���,��)�)Hص\=��z���-(�k�[輅�ƬsX����E����b����
X=�^�A2">~G_w�Y��żr��lؽm���(b���fX7j��������q@7��sW������B%�g���C��k��Y� ��}�8y�c��
��s�����A�_��q��%vb�N���,ڡgS�f��s<�Sw&��̳��l��q�uU�7�%��Y��<�$���f42*	k���`J�J�E,�����VÅ-ak�nRK�4y��!����� ݃��0�-��{� ���;k48Bm��x!˟삠M�O+9l��?_�FWI���"t���fȗ6��!�5�2#n�b|=�H��V�;=��c�T�p1p
�b��8��´Ȏ��NI�yAnα;�Q\#5�f����]�X��!��o��ʓ�{���5}cz��i,�VL����h���[�/&�hv�Ű(s���bY���]x��j�*��Cz�B�ϱꑆNqˑK:&�x���խ0��gՖ:�uכ�b��(tL��^UV�n�x4�IDH�k�Ф�'�~���G"fϳ�P}��\b��ng�x�2�s����L뾳�H"��P��� �;6Ga�����dH-�bs�Z�&�y���9U1kL{0@�V�Zg��#э�.f���Jn�$k7D����f��U_X(�I$�����Lx��]�`O�Qkn�L/#T�_��7n��g4z�4�km��.�_t�*�j�	��م��
p�$C�:���u�ஶ2�GSS)$��������;}����޳9�gQ�]�ĿʠN��"�j�g�U	xp��J
��Tw�0i�v��<�����j��3®�����FI7>���a��8-g
������+/��"Л�N���U4���z�0]dJ�ћs�n�Q���W�xF7���zɺ�7�֡���hۡ4��ݺ��8�S�XH�g�҂U�o�	�zup��0��V��2�G{vL�H�S4�ڃ
�����{��,La��/���ϕ��gZ��Ҳ�����U~ů�P�<���(ӌ�:�3\�梧1)�Q�3�Ӳ7�� 
#l����Mv9(�9'�RLWAJ��α=�������w{�]��b���u=�ϣbe����/��a��'8p�sJ�mŉ�Q�縜�9�,>-E��NT����:�f(g�M�u�x�ok9s)I��Ha���3�������J$y�g,�A�k�N��5��Ʀ?s���b�O.j���HuOMWJ�1��V��j�=F!�%]�|�C�=�D�CU��/�C,�e9F�탡6� ������������\a�l��X�/s�/�qo�)�wX�����2�G��D�O",�k�D�E���� fo�ú����2�U(���=[���U�! @�r�yä��(�AW͛|�J�;fA�SW�����d�9��j�'1�>D�|c���#w"Е8��l��ƝP�V�?l�%~�wo����q۵KQh�X�M���E�)'�T	�ygN� ���2����<���y�|� �HD��0�ɫ�����ȗ���Y0���iw�-�XjE�� �!�R�td�NZE������C��m,DOu���J2�H�Z驤���U��e�t:Gb�h��������=�����7�����xL�������.֞z
\�/2n��y�э�)�0�n��9��%���#���` �n�O�*����+$mmVt�&��	h��Ғ��j3jÊ�a������
���ǚ��^Ĩ�(BT4�+H,tk���֫Ǧ�Ǔ��f�jӈ]�6HU_���'|�y�ޓn�E�.���7Xf��w�/ȉJ�U��2���|$R�����f���Jbč�Z^�BM��`Av*Y���:��vz؇����Ec��'K��O�Q9h'��<U;ޕ���&�Kl��T$��2f�[y����H%�W�$/�@O.�3 
���n��S�Z���ln�qm��?f�`������ 6Q`�ܧ�J�ٜ�1V��\0ѹ�e���N�z��,�������B
��??0e�3?n�`{�Ik����a�[��ta�x�K�L��w�Q��/n��R��F�a�����(BM7c��"��HfO�������J�Vg�_V�;��}M�B���&��c���*���GIi
Twn]ͷNBr@�Fj��E|a��+�.���Rcl��)~��e�p�\�Nrڔ����ms�)�K'���E�s64����ӣ�:R��H�o@�gņk�^|�Q��lc