��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|ۧ[���{_H|7�chb��kS����L��ݲ���N�ƬK}�ڷ�!�rT��Y�������{L=���j��=��!���j���8L�h5+�}�=���jE����җ�&	c�ƴIlנ���Xh�b�bh0��w�.Ǆ���.�*4�'���������`������2WF��fu3�[��NK��˖�¥��r��E�_z�<q;�8�x��8���̀ i׳��qu�T��S��$� ?E��ӗ��+<�J�F��F������K5�H���*���2��Ka?/_]�F�W`7�(^"�g���#�4��Y�U���v �#}����.4��>��+�}���l�w2|�v�=<m�I�z�e�(�&M��a��)<�5Zq+�is���r� �����3Ϲn�z�"XE��0Ӌ�������Ȍ����(}̩D�������L���f��������܃R��T\�8�t��ϧ�A�GU����&��j^.�bAڷ�$�%������r.z�Gly�M��x[�	�x���Ѐ/���bW�)����>
&PP]!���=��B�
����g��\̤�+���5�2#,�2Ys�@N�����l�Uy�VDc���л�Je=<���H���Ԑ��	�_ �۶��.�_�����J�S#�*!~�.�	H�!"��%�g�v�X殂L��\��<p���]���Vn�j��k�G�I�
G�c^
`h�����3�
�Ǝ�_���o��2�����ļ7�XDs���D
*��/0"�8[���3d�b�Fl xHDA�GPDX�ny�s�r�M����~)���D�6�v2�m������bT��33�T��#x�UX�s|K]òp���������Z�g�z���gfW��h�A��b�[:�pFm�aP9(��ȕ���qX:�	κ�ӇU!�(=�u�wz�]�C�8�'`o��rʯl|��I�e\'N��d��.7��-��Y?J����g�Ҳ8h�d5�l��Ň}l�>�!�u�Rz�{�h�#)��.f"��K?�m��A�&g+I�j���UH�	���p��R��x6]�c�=�
���(�
m������_��D}� K~�Ow�F"[�_��$��h�f�%e��=�`;��4�*l�-��'r1l�Gp&c2��c���nD�c̽��p�*�O/̲A���N�_���>�w�J�k&��k��
�D��{>��Z/��b5�M�Q�g�}�Ʈ�]N�OM��=��uI��]8>�ez���!Ri���5*D�T3�����E�W��,�ܴ�d	}�b0��|"�� k9/�^wQ���̭�d�Q����QF:G�������YT��E:�C2���x�Αf�Ў�dz��s�͈R�X/�8bT��d:ɓ�2H⒁������$�%@s֚�|���tO���.O
r�c8q�'�;�H�#\���kx�D�zg(�K�/�υ���q[��$**R��r�z�I��xp���d�C���Æ0&Y__��O�րyy�:Z��u}	��y�7�CL���b(�Lt��8ዉ�`�QZH��;`JX��KiX!k�� �i1S~�ݢ�k#8k_����܁t�DL�͵�%Z��o� )��>�������[/y����pVH�d�K�!֦0n��P3�%�����r���R�ċ4燎^
P̃0��L2��ՌW�l$R����<:���k���KY-�[ ��ˁ�g%�$�imF�Ÿ���;`/���_��M�l��\��x�?=��Ƿ7(NlZ�p�y)������#W��Sc�\
�	Ç�y�J�j�P��ra�dd�=���J6m�����>����S����|(���sƊB�~�	�b���T����@l�`���ou9���n�
�O�x����?8rc%�I��	��Ws_�V��1�p?U\�C��F�S�i����+�|���5=ф7���RJ	w����1�S��V_���)X�&�D�ӓp�Z����g�]�e1�帩B�.o.��E�֜��?B6]�"@^[�9�D�v-��E�vy|ObJ�������Fy�Ԇ�w�4W5�z�v��Z���Qw2'��;d���Z�bW6`I��̪�R�_MZ,���qU�YG{쯿_*0�Ǧ�y�Iv�[���W5pn�Op2>(B�*W�*�<�,��#����m�c�;s�p��Y|	���{i@��|�g鉜`
���B3i3�M�C;؆p���S)�9CA|�i�w�#��I5�r�N�u�Vf�P��sX�2�K�3��1\�h=�/��#�gğ5��e"p�ns�_]ā��L7��;?枖�C�c�l!;hS	��������[���n�����QQ�8�;��3�u�� �0��k�:u⭅��ez�qfտ{#�|����"�:b��b�d��ös�k�$%о֩L���05 ^��̑�e��>�1\j! ��:�[��b��,���=�;��bߟ�#ӌ3�8�G��Ȏ@�||��=��{���xE��j6�|:��Z��aB�����wt7�FUܩ2�Y�����2�l�7��Wt��k���3�G����o��S��y� �KY���:S�Z�y�\������2'��mckpw;p�F��t�\� ���,:"�)ƨψ�7[��	�n|���%bՃ���ps��D�nȻ�M
Y��e���)X�������`w��2��O[��i�j��\�ǣ����#�_�%�K��bdj����>�Tw���qb���vι�%�˿�E�d{r�u'�!#f��� ���yW�r��hq��)h:��a�ི�M���a@J�hJ����1��@5�<���G$|��@Ul�Ͳ��m�ϲ=3��<�e�,�9I��LrJ]UZ��l�ܧt]X�fnf1Ճ?`���-��7�⫘F!aLr�J����HC�&��Q!`�oXp4��!g�W��m{�e���v���)��sp7=Q;�)�)����M�R��	��B����X��I�g�9Y*�q�#%�􃉔��{��>�ZL�N�7U�&>�D�K�K�mЪD8�P�#��v��9�O�v,%�/��Rbh5�m��:0U!�����/�G$��3}�N�sR�_:ߢC�/����6��\!�Ĳ�ǟ�	Q����9���7��lhqY�����aNq�Awi�����dF��J����eS� �V5��f�%�RZ��v��,���3=�z�;���n�d
�n-e�Ie>7V��o������E�g�u��6u;%���%�(�Kf䇁�N�Vm�cA���%��k�q��_G��t���7ɐOht�i��C�L�� v�%6R�#�癬�ޟdu��r�\��%�=�Z��d<?�~Z3����P�CȌ4@}��-
�Q��,d�C9!C^�gl;c"΁��v�?�-�)�j��;$#��Yp��g�ZM�?-�s�o��+[;�w�v��Ff30�-̄�#p�E��+m��-�y6�q�~�W.�v��76���c�PG9�?�e�&�����BWFq=)� Ղ�J���ut�V�~��V6^�X�������j���M��[ _/E��BHm�˱|.f�x!}�M�'p�A���6³��o�����V�i�����K�6͎��M&��r�*
��-~�Q����2hA���;l���W�&<3�+F߭\}��ϑȮT�vՑ����$�Ɨ�U1��M~X���ԟ��/��m�@��>���+h���˜7ĕ�3&%y�9s��k�8��B�w[�d	
��1��T�]�5�n ��O���ЃMĒ�>-��k�"H$9��a�����}�g�b�$#�������˼W����w|(6�ҷ��揲�<�v+�h�ӏt��UòNM�����A�}	d3"����M�h\t��/T��b��E$���h�P.�*�H �T57���Z.ݣ�匲�9�<��6�	O^����]���I$N)}7��,1#�;F�59L%��v�x�`RW��1A���a����'GY�1����N6 ��G[o?�`���+�-�mQ{��娻	�Y��1�,�M���͘���S��O��s�\�ê%n�ӆ{� /ŵzG=��̲����+݇����O�C���3ޭ���ډ5�d��ٝtR��j��q��A�����ot_���v�?>Q������J}���f$�һ�Av��d$��^�3�T]乮 ]�^;ĸ{�lo�T$H�(S�CZ�Ԇ��j_��.���X����e0v{-��!�m�����1�����s�a�Y/(��w���S�+�TbT=e�@I"k=xZ$'�8z����ß�|�Vg-�j�����h%�x��RZ8����2�VS��MݚC��;P��8(
>��m-$0F��!��N�q!,��}Fs�'@R%�Ζ}�O�����Wl�z~���%#L�/;AB�GBW��
�V��]��`r��Jd�ߤG>>ce�7��%�LS���yw�a�٬n�MVl�x\0�g?L�0� |N�IW�h�y��v^-�E^ܥ6��ܣ��9�5P[J�+�wA�(�����X���_*	�>g��ed�l�}4+.s��k/'٣��l��ՠ���9`���$���G��|������Rw�<��e��u^},�XNV36�H�.�7x���� +�(Ǻާ�Xe�)�'(ɠ 3��\O$o��g ��Y�vfQ����a,"���7���V�NJ#Y`2���ϙnP�y����&5�Ȋ��> ���ꚸD����_|dm1�!�l��y*�`��.�Z'���EJ�b��y
���kW\�+�)����?���=���A�ǐW� �|^��v�ۼ���J�3��Is�%�W��՝EK�
~R$7H�AM�Y�A)hC�D�:�D����nY�r+.4u#b�ި��
�ES
ܺ���P�bz��W�:a�`/���'��k�?�-��h���$5PZ7<[j݌\���)t|�xso��G;%���}��,���~�"g����5=�=����3�L�u�d] �ĵ��4��fu�4܂����U���H��HfFo�5�	��|�w��1}��9���* �s|��$?�-:GYnc��D-���	����cҐ8L��PW����}w���'΂�;�$��5B�.Ͱ��~$��������_H���:s�zTR��h����ɴ��t-
p~z/���0����f��Md��~r�0���9`��Lc��}��Vki��}Q�ϱ5Dԗw��M2I���9��ׅw�N�(�W��
������ヨH��I�ؤk��*Ӻ�mq/O%燏K�!FEZ
�BB.�5a��+��<#�>�M������:�BPt��B�L���5�=qI�4��3���6l9l|,�wG����`Qh='�	�Ty~l�*;�P�C䄊�b��c�"&���I>L}�5���Q[�Yh����]k+#QE��W�;k�/�f�}l (�� �Z��u���'(~C^[ ���!D]E�O����U�G!���T['����[�8�}ʶ`��(�(��wfm ���p�v^U����>�#sq�l���ƯŸc�o%}�#��<�%��D&_��=!}�چ0E��hh� �[V'${W�d��#}���o|���.:���$��
gk�bΚ?t�%�(
)M��j��	�&���e��\`�ӻ���6Q(Hղ��yF��T�¤�?���جo��o���}@����*U�iЗu���G�bx��o���[hLU+(/5	���H��@O{���Y�pj�欩psʰ\Q���[�c�1qV(�����jb�i�Ԅ���>���R
q���/2m��JH 2x>���ʶ;�OD�� �S�����6*�XF�"G>
������m,Y"�$��HS��_���"���������6��ҘY� +����`�[�]�5Y������wt�#X�D��ۦ\�{��C��D��4��T
�2r)�"i����?4&� Y�ud��4|�eK}��N��5汲/Sk�~���:��(�*�%"{�ȁ�6�&j�[�w���5wK�l^��=��,q�������e��9.0D*_|�Q���55�ܧ�]��d��}&��YS�뎛�6����U'�Μ:�fa�uR�Q::���R"��j�s�B���kF�X��3�f��M��@���v�/��M���WW�|��P}�48���1�Fd7�#_�X�9�z��?�±��̆Hv����f�BS(��Wh��)����Q(�GD�q�iP���-�����L����9�%O��s������D)Il����*U��	���?�.�z�`��_����-&V0W�L�-�	J)�9��b�U�=d[��d|���-��3ϤF���P�����7�d�
�"��b�ۭ��喛.�S_q���̵n���Ǫ�����<�ז��{�� (%��Nx�� �eqO*Whs����	���lx�z��ւ�>0�e8vT_�p��D�%8�I^t�vX(X*::�����v�)�k*yQZ�˨��󐩍���Q��{���y+�(�"/���
ւ��x�b!z�{���'h�$l��)���G�X�r��-�=���s�xP|,N�E��	�u���!N�����f幍�j~+vԘOm�!��/4���,����=AܗS���%BU�+1OS�=�Rv�.+�d�J&Am�k([����=�JF�7Ǥ��Q3�\>@\�`�-��~7	�i� �j>��UV��:�^(xg;��(1�)й!s_�I��� �ϝ���<�!_�a��I�B�b���,�1b`��@����EU�~bwP�~�6�/�+�4�;0�
�dv�H�A�;���'�4�i'o�4&�3R P�ӯEY*�))IX�c�ީE�����2X]g�z�61;O��ׄԥ�ɽxT>��+���T�ζJ�T1^��(�����sl�n��)�������Q��J�#��P��0В�!\.�o ��t�h.���h��.9fh�Ⱥ�FN<��is�j�'��m.X��[�����a�{}�I=���ؖp������X�rW0W������)m���+�����I����+CI�����]r��Wk,�oE�D�����g��U��_z��o�	x�%-=��a;�ؠ�\�&��QA係�
|�%�|[8xh��<U�yn�(8��u��?���,>��Ra�R��-��$��O�<�[�����3[�W�D3�;��Ū�n�$2�E��>Ac��G<�\n�o�i�_"5if�m�l��K�����KCž�\b ��yb�&>O}���e�$|!��a��k�˿����,��4�ߍ[�(�NF;�9����ʪ��t?6J^�������-�p�����~�(�K���ZO�_�[ݧ�U�˪���'Ǎ��y"��{,�n���q5ah3�N7�C|�4: ʶ�o�ae�JWRW���c��t�O�O���M�- ���}�A	ǆ�n�ۏ�=��z��ƣC��ux%-/��x)�W�[vs&1$�y��X�6��̟9�0��-%�(Y�h�uR���ws���GU��xkE�/2� {q�"����7k������x42���]��g�=A��e"k�;H�k�x$���k��̇'��*� ��t����Y쒗�\���%(�Z|1�r��Hi�<��`��z��(���!���?�;�9P�4o�Us5�,5�&R>J��E_1�`�$�I�X��z=�b׉����f}�N-�'��^�)�ύ�����ԛ�K��"��Z�ņ��Cn�F�ۯեCt�~G�z1,�'E\�U�m2\{4����ټn��z��#	�
�/Q��a���o��b��RE�����zf������p�l��:�#���#�����+$y{�|�J���FՐ��B0�?%�Ξ�D���v�N烪8�s�xg(�=T�J�5��>C_��*�bKGW�Z"�c.a~�hZ�T{��ΗdB���&��࿎J�\>IZjo�y]�G�ѹCG]^/�� �xm�g$qN�T�*Ȟ�k��<�Qs@�#��Zz�`d����L��<�}�4v���_��iTl�<��q�WJW�+IR+<�}�n��}6~�V�޹b�h������mW)t�Uh�"iLN�u�O��f�>��E����쇐Zl|��x?�.0Ys�%�MO�x��l���ҫ��~�na0ǖU�Y����3}@iy6G�r+E�ߚ�Bo̪���4��M���\9Хt%&%CI^اq�)��<��#m�"�6��=�if�Xz��ڤr%���0B��.�b����ϟe8�)���^J��݅J�=r-�˿���?j;IKׄ00Vڬ�R7Bt
?�7@"в�ZT�H���m��VԂ�W����>�9��[�e�F��(E��´II�B�Jj��aC�oW�%��M}��n��H���уʋ��(8�Tkn"_+�#5���DcHH��*�o�r��cs���H�� L� Qm*���>����Q�vS��D����E��A����n�N�T��Ɂ�M���Nz�=i�%͜	��֍�0�m�&�N��ھ��"�r?>{�b$DV�/ -
�qwv��i��>��!MVy�J;/i�\�&bN������;BS9�x[�a�����l���ɭ~��g
�gJ]@F���$�����0�.�<h�YzC>#����жy��C<���u�0�� 1MT�8U���$��JŶd��8�@쒬+�C�]�ߓ�mzM���d�?��<S=�ݤR�^��hl���f�l�-`�H��c�A�mU�?�Eě�u���Ж%dfn3 ��#�9�X��G����L�����q����T2X*.,�u;ɧ�?�ٲ����ج�5Z�����4q5[�q��:���O��i�� 2J�'�ޙ�%E�G b}%�O4�|��V�I�:R���˛�Pʬ�Aώ���N�\���ˉ�Yn1���d�,v���{~��C��n�)���D�	v S�t�[;�9�q<YJ)6"'���E�� )L�������Nd�q�FPG!�v*��m.�gG芨��p1�a���s��$��A����izRL�p&�����JV�I{8v��A˕���Ox,Y���|�M6�s�>)�� �YX��������!������A��!�_s�A�@r���H�R����,�;\��s�}�h��I���i$(��*��x�@l�[ 7U���v�ȩk�s�__���!�q����m~y,N��?g ������o�˘��WU�=�I�6�q��g�~�@�K2/��6��d6 ���흙j�[�k]j�9=�/����L��b5C��]�U�e�k�M�j*���^IjV*�+�wO�O/�<�%�wx��kZ�,l�Ô>瞅/wT��q����$Q0@�+����j�L�ı��z�O�v�H=�Ď.��9���������hȑ^;_VrJ&���6B�ӌ6��6D�����([�HΉ�]���m>��p��x�H�Ȱ�u[(=Isd�'kl��|z޿�G�M(�p$3��!Ǡ�rO���ͼ���)+��V�%�|���0��:tLz��}	��b�O�UrmS�ۃ ���^��I9+̆��~1cu���?Ϣ��������I�Y�1(��΀`A�#��g�؀?�ą�i��~��< F߄��@���62C���ISdx�\�2D���k�7b�֎$�e�h[���e�p�5�/�ӛ呱�Ϝ2Q������/��I���FN.w/��)+�{W�l7̥0MRro���o~y?z}خ�R���>�#����^AX";�
�*�5��s��^i"�6kiG��n({zc���0��HS��4&^@��]��+?a���˓����2:�o���v�o�����I����ӑ&]첢Fs��8�x{��{2p�_f��W�D?�P���L�������Ƹo{�NG��N��4Yc��5P�F���idm�A���M�݂��C��`��J�ǂz
<��"����ݥ���7ն諲Ha�'&@n,��7m�@�.ٲ
���yվ
3�ޙ�&�=4�毠`I�y���:Xl�l�B���[���A��i>ׇ���Of�-�N������=��̙r��Fv\ ���h�����w@ ۙ.��2�c��#�J:�� �\�E����GWMR����r�໢~=���8�;X�av�/�+�V���ߴ(����}��+,
Q�Ȣy��u�Tn�@Q'�CO��|( �vg$������H�m</��C*O��.�p�Ph�����c?�����F��O�ŵZJ�$��̷��C^�O�C��Ҩ�A<��(Y���;?B�\Y���B��	uY����L�YPV�h~6��6�O��� ����� ��1��� ����4t�
�`"zm�>��_0�U�Z�����C?J�{ Kw��Fn!u?4Y#��H��a���"7n�G|K24�yU�x��̢�����s��V��m�o䷅������Q9�:�0��R�o5u���)9a�e��~q���X�4?5��x�[�4���Zۆ��֣����q4>*�z��:Dwέ�Fh�i�<ŝ�p߁�D���v�Ű	�KAN4ﾽ� �l��}�پ$}�)]8#��'�`�����y</�`R�	���Õ�ډwz�츧yT�=�kx#����e�$|҈1S
W<G��g���v�j|�%~]��K	C��Î��Q"� �Լ�ÆAt)������9x�)�_�a̩6-&�ނ.&�4���Ѧ����l����v�5(u9�ߕ�_;V��|��Dfl+�<��2�@NqoQ	fϵ9��+���뤽��7����0�=?n�Rj����Sf��j� 5�����XSԳ���]�����G1+p��J2�`ّ�dTu������@��la�L�KX�V�45�YM?���yV�2Pj�W�1��Vj��$c1����({3�z����įJ��Q�d�Q�3��;��)��yH�=��^F�@",w��l���c�8�j��IÜ�����r)��������x���s��\o
�6� }�����jX�)fv~�RsW&L��x #u�f��� X�p��h($O)5�q?=��0z�K���E�8����?�vq�9$�@��BN�WΘ#έ<U�/�k��l�،�r�	vf�y"��z9n�{�<�[��q��1)�\���x����3���}��~����>�(��C�ņ}�}%02���d�ݪ��pr+x2�tJ6X�g��|��/��2d�@X�9���'�T��QI�rm=ʴШ�bE|��>��dDUߊ���(��e2g���
Ŋ��D�`�Y CO�@��'�A���D'}B��ӣ�)wW�O,&�^K�6�E:�M�:����qù�I�͙87Q�Q�HQ�*-y�i��S^xe��Z��3f���vbt)K��д��m���Qk�E���wU���{y�(_+�#�T�v^ؑЀc�.G�b�
� �0�������,?8�;����r�`�.=��mi]z�6�!7�<:d��Ǧh��b)}�T#4()I�gO�HΈ늜�
T��̟G�������E�d�#��>D~����9�x�/�s�q"�R��I0���c��z��1v�A7�
���'[gi�F��C��5VE�;6��
^���2��60/Z�йR��)�X�_�Ě�Y�]��n�K�P������tqɨ���DI��D��5��ov0�?�/�G}�F�PP5x|�>�uň���+&��g���=2rA_��f�w���jR�V���k6��n��-H��>�9�_*�2�NnX�Y����u�T�BXwz��sM"�I�ڀ���c�?C���͡�>�`��(^���W()��jzJ'y��� �r���m/+n�5��w*}Df��T8ig�z���'VW��Z�0ē�X��$ ��L��;F)CU�N�����	�A�U^}�"uJkm�
�ӳ��7Y�:����{����|#��r���ST�ŋ탭�:���c����<@�<\U�N6��

�Z�J�@��i��[G��v� %�d	�Z��*�VU,��gE�O�<�!�������������E������Cxj��s���C�G�gj��7��C	%��Y��@���[SU�&�V����b��u�$J�`����ѷG�/��v#h�Q��H��AC�)*��ڄ]g�T;"�2��o��	X{�>5�R�y�gk����@����		�}Yh��@C���>��~�kj� OF{<$�m�U��fӘ��nj3+�k/u�����L��e+�P��?�#��h���.�R����L����L
LM�%�FU{l��=R��0�{K�:�q�6�H�����L��-��H��|0Y��*c��+@?R���5��9ku� �HˀM�_#$�u?�%��#�c�C���5�DP��]AWw[7l�cՏe�9N���'���_�V���2z�%���VS��`�&��<-y�V�pPD��]�H`r�G��!�@8��1^0uY�@�~_�P��J�露��W
HDַ�A!�b���oa����RΤ�D�(����J��q���~�:.z�Ib�`9w6d�~�Z�7m=����LƗ�A�@;�h�B��0(�h,/�ݲ��ƸnDX���W�jb��^=���~_��K�$����u�q;M��_� ���[�bZ�#��(�)�)�`�ڒǽd�� ���W�a�o);�"����jXU ����y����gU!/����_��t�\k k(��b�6BԢ�#?i��x�Yk%���?5G��R���|0n�Uh�5T�E%D�&|�J���ܢ�g�	�8��k��k�@SJ�AF�U�!�F�9 ���_l=��U(t
#PL^�7����Ӵ�~η��:��\�����7W�MD@ׅ/���롚t�
G�0����=x������+S�:���O뙮�%��1���@�YꞼ���i��ܠ��2��$}}g��6�i�_�q�1dh`���;�0��˩�6�������E��h<��ޏ�Ò�7��X. xr�8�'G"f�~o:Ba�n�x���[Ɨ�p�(��ԞL��*8��]n��Q9�(�@�댒z�íMo�X\�1����ՠfO*^g��3(�>𣏕����g91'���~�>�h������=���WY���)�lԲyr�͘�].�\V�i�f�����Y�
P��oa ��<����������M��&��pE*�<�V���JMq�K���̺^�9͔�r�'�8�V�F�#dc�@��fȷHg�[q:cD����w##���Hi�R���dt�n!�x��&B�(>���2O
37k$8vL{]�,�s�b��c��YJ=�稞v�~Ϣ�V��8 �>՗����P����wp6n2�%�u�1+�I�U~G�һ�)Z8'�J��+�=��,0�<%���E����H���d�s$���%��'47�Ni�i�����	�FO�ͮ�z|*�Lo��]���Z��(�R��P��+�,�K��"�%.�R �/4X�e��j?pe�Eܖh��ZĘ7-��e\�-�H�����-�����}��g��F�8�n7��#؉���	�>®��؊n߂3�c���j��<o7��EpӚ���'�&f�IJs�?O6���B�{k��n��9�z�Q�0������(���:B����������|�D�u=i����q���c�X�3�M�r��.Nγg(�Z�AR�H����Qz]�c�x�eJ�"�fK���lM�HiV�X���2�S<�̮L���M����˝��JL0�'�d|���=,5�d���c��`��������6G|��y5M�ܻ�OOa�I��z{b]�f��k��{��p��Rn�Ai\f�$�g�n)$�ϋ��m�jOMI��!���m�)�n#�l���'���w,��_mM�T�P���~�ul�f�*ħ��ǳ�5�7���je�V�"	{#)A�w'�.<�iUp�3G�wfy0H�#����ԫ+I���ad��	�W)!Li�Q����G5�W>%+����/����s6_�`�1e���h��-����D��m��m`�FW�?}�i���60�5V�"|�t?Z��d�j�o�x���G4��7coӮ�������*�Ra�g=%��,�)%>W����@Ǐ��}�)-��GG��e6���	��߷ᳯ�&��}����)�)��^L��X.X��i+����".3 �aOM���+���N�0�}����V�Ƀ}��]X�6��<��o��Z�~؅'@!u�����C{ו�r�/g��e_X�Q
Pq2E�F}\<;3LRO+�Uy۹!�9n=i��14��iYkHJ�*�h�
- �� ���Fo��tj�
���Y4M��]�<9��,27�kd\'(���
��QG&��%������S��:,��E�ƌ��(�}����k1c��Z:��� /��n��K��b��K�v�_9��Y^�"�Y���+eR��2wNu��x�Eﮝ�^��7�t(i̸{K6b���s���u�6�lt��`{����Q��ϗ/	GXv�'Q�\�,�M
8N�<�hކ��]#���$#"XNs�tr�"�c��]w�u�ţ��V4�8�J����)��hInΩ��6�|�XA^�#�R/g��>�|Ӭx�0Y�^פ�6��A�
cI Y��{�޿�=aRG>F�eJ�&�ĩό��Q�bKr�h�����q�et�DoM�^m~[��k��^�W9Ĩ��lF��_��"�'M�����
:�� �j�W��Д�C��:18E4�
s�K�g_�)ǥ�������bA��s��b����ċ���_����}$^ʊ���#�� �3���<d���Ql�N�qyv��Ë����� �����+��k�Y�H����6fG�1K�á㧶nD���O�	xſ_Dj�)�i�&_��g�6���fۖ��"�N�O��X��]��b�ҽ�hn{㢉���&H�C�������W�_v,�������>(.f�v�
^����b������!Fh�fJx�ĭ�f\U�9��8�1���F�VuBa2T���c�k/�r���u�b��Y��im�i ���n�T/���8��r
�E����w�! ��O�������� ���Մ�ε��S�Z^2c�����ɘ!M�L���m�2������5hvc�6';�̣:�{�{g�6F>Gf�|l��M�3����]Y�㴝���Y�9E�n��3�f��u�x��[����5"x�Zo�f����C��w=[��`����/��`L>7}���>Oy{�2�	A�ٻq��E����rx�ݸ�.t�?�!��q�=_ ���[��B).����-��Vؔ\�w��g�!+r�z�rB21�:�����X]�`���FE8''�s<���s�_�Uh�4ߝ�>�?!֎l�m�!n03��$P�,�6�)�!+C�6+w��O~t����Pte�v��-u��v/�՝.����,t >�<���~P�D��F���g.
}{�k("x��[v3��|3�'��5gAw��hk��(Q@��p'1|�3"_��$�4G�ʞu���Z�Rb��U��ym_]���v~��Q5j�zC��21��8Ą�S��y�%�G8T�U*9EkX~P��)�K��Z�Ȼ��\�J���]}
B�&� m��3�Cu��vi[q�G�G��wH�Y�+'�Q�.����U�e� �r�5�^����Ľ�xy;���i��L��7>�L�_�%����/L�;��p"1q��Ҭ���qJ��7����2�3S�kY�Q� �]��4�I�E�c�9�M3QOt����H4�����?�ǱxrYAr_�E���j@O6x����A��}�����6������oμ�������p���ȸ�"*�)>��*��D87%f�"PV�+cG�X��l-r��R�>C���0K6��q�@!�������s�p*�h�ws1��!��K���Œ�"�Vi��H�wO㵾�<TY��ќF�]00N=,�	�>6S)8����'`�CF^?X��Us`���A� X���P�]�6c$|��b���:�V\��F(N�)荨����M(�#/x��@� M��D�LW�9cO������ׯ�����oWtz�@/��Xۼx�=s���6
z��8qρJ;ߊ:=ǹ�c�,�,HM���A�\���k��u�%�Dx�Dq!�ͤ��ȶ���T{�ƚ�wP��0�[G�JO#�K�?;�mn����F�w���/t�������^=�zƜ���
�#=_t������9ɱ���$�� w�p�U]~���В�XrD��q�q@��r��
Yk�s��p��	�P���^D(�����\�JE��S���hLw�Pw76cy�ퟜ�����uT�ۇ[�xioU� ɶg�3��es�[�O(S�~Y��#c)雩�<����h��F�|�+��*f@tgi���fO�E�S�����|d�h�qV*m��5^o���=��ā�pg�X3�*jD�K)��}��jR�ēv�[���c�s�F ��qX�OBǩ1{w�e;t^G�xp����5��eɨ�9�?�?��������V�cb��h�j\�!&Ʀ&���^�"24��{q�?�H���tk;xb�1y��?%	~�q�țٟ>��r�Q{��G��;�KLs��xZ�\�t,,��HD�ѳ{;À��h�]�`(o�䐼�<f��!$E2�|�J�vR��R-��'�!���rS�V�u움� l:�����o`h)s��kIoȝ� ����x�65~)�^���ȧm�p��i9ND�������ϦՖ��/C�ri-_���˜����x'�B`L�+�����`f�!$����d���j�*U����F�o>A8�b��8ɥs�)��Z�ec9=}���z��z� 6��%㺖pv�	�S���A�R+�Z�7�e
��+s$���H+1^+R:/�ġI �����Q(۸�ї���������EW�,�@��#� ��}���<~b��2H6>!:v�T�J��Xm=��d����KSs�J����j�'L�k򑱳%�&�`�7C�4�r���A
a!bv@���q�����j�a~+R�QO�~k��ℬ>�ӚL��j�MK�e�rCK޲��`�'�H����C_+`n���t+�5 ^��'�R��Fe�"�������s�,�i��#x��_!�.������-���mZ+wUV�n:�e=�:��z�=�����v�]8��S��'�(��+�M��[/�����|��5�Kzr�1����1��`"v�{F��o~���=g�&�;���s^��,P����ѩvf�S����,'P_�9툊����n:�����N�8E��~�_a�R�#���C�f�G��3�@-�]$/{N��M��uu�ߍpq�Aa,Vڍ[S $�^�m��ؤ뗐��R�ֳ�=��ׄ�?6][�U�*��+��C=����݇�լeD�!HW�
���Ò�75)�.e�E[��SD�+WؗS 芛A�����X��K�fGY�ʻ�o�3To�Ҍ��	A��ְ�̑!�l.֋Ap�n�O�E�F�$��R@S�n��m��1n��v��A��6��=�i"��?�M|����zl"�G��Fз��Y�5�f���]��(9�F����;V��&#(lDd�"D{np �lP�$Nۘ��#�krމ	w'��X�E���V"	�~� �˸rAF�� |)<�PN���qR<��w{�� 8z%@�5�>�K�<燖P��M��vr�Ȗ�~�FLc�G^Cʗ報��3��R��X�`
���u6�G�s��p�j�{S�Y;�t��0�qb���&�W}ly_�ܙo6�M�L�jX^��B���B	��Z�V���7}�e�Rř��kV�p��r���/ �@�㈀��������S�_I�G�@����V�Ҋ�P��4�Y��(�;D+����k�
0&�ɶ٤��/� ���	מ�
�m�k�<�)�6QmX�3A�b�=Cی��a�*e� 6^3��ī��f�ڤ0������o>^=�w{,����=rk��3�p�*�7̆`�A�,Yx�̨Jk��^����쬤g�Z՟�C���yKi�,�N9|� {�3j�<�̬ �dڷ6������� �ъ�_�Ԫ���	c�K<�j�Er�ag�@a��:pu�hh3�Q0na�篗a���*_{7�%�1/����xU���7��&�A�9kJ>�����+�$����%������p��F���ؤ�!+��\��s�$�g���b%AٕV(ho�D1�C}��ޮG�ꧩ�7(dD8�hQ	+-�SO�����,�2"-dos^Fl@F#n�o'�S��a0�~���Qbo�#��3)d#ԇ�5�uXK���'	bu�7��)�"����H��d��<�	���J7��gޞ��  ���{\�� ��檲C����3KJ+�!��n�W�8-����]��x9ߐl��}��l��D�I8����pQ�h��@�	4(1�Y�� �	�����}��2�:��m�ezxĂ��?�P�/�7n�^a�J�kD�k9z���C��t��3�H�::}��z������8�"������0����j��G�n��Á{ʥ�QmNlB��c�A6X=����+��Vd}������SH71J7l&T�Ǜ��2Dv���D1u+����c��e;lhk\��Rԩ�Ãc��*=��l�K�j�����~�~��s!	��|e������������r�8g�T��-��l��I����{��1�[���wɧ�M�������0��Z�`x#�_���!����4d��ς`T>ZY|�70Ш̙�P�e�|f��}l�2l��q����&|ol��� ���>r<r��A6�ln�U�	��RK�C�Y�\���������h������GD�CZ^�Y�\���OM�s}\�1�,B_���Ω?��G�-���P�����}j_�5��y{.6�j�ض�O�$�{Mr9?Մ����Ӊ�fb��Q,d��0��_��5�f~Y���\�V����c��x\
�=W���P������-�G���uW`�eUҾ �\BX�D#Σ��=l�O^�~w%�]cW �>on�kN�m낀\��H=�_]��Ö�#�n"�gK�j������| �e��u8rP���kI�Tv~U�C:�/�.:����̉�0�J�o ��[pN��$H;��'_k��d��m�d�<��*���DY�%N]{n��F#��ke-b�%���JA�z!w���y#��g9g���!/���П��~#�����$I�n�?�z�W&j��� �ޓ�����5˟�6�6���t�U''w2��:��eTw�t�b�� L����c�xI��V�ׄ�$4�?_U�4��k8���"qE�=aAk��{m|�(���&�v1�a��cVc�Bk�����R` 8�`f0��2o4���e�2��r����-"ǻ2d��>��ҍV~�T����f?���P��%���.�N�r��aB"z��+M`I��z{��'�F�"����ߍKQ?�P��Tr��2£��f��V�ޒJK>ͪ������*r��)jK?aL��y����nȼ�3��E^"������<ڶif��sP�o��x`
���Ϡ������iM��Bvx�}k2v�H��k'�c"4�i�$i��$�ȜZ�I6�2��Z���y�J0�����sLHH�U�ŧݩ�%��J,�Y��Cr�9�i.��ȄSǒ�s���a�C�f+��C�Q,�j��r?V�j�������V�wfL�7�[��%Vg�	�Xʆd���=���D?��&x��ҧwaS>�Q�!��������:���3�D�JQ��ڹ��iڝ6-�\��'��^�&��r��"n����������$���"�J�J��*����ݤZL�@�e9,�U�9���u��� ,�\ˍ����a�ci���1-iO����9k©{ҿC�$�� d�(sz��`N�oZ��Y�EZ�~o�o�O ���;�>`ck�[������/s16���d�E
�"8Z~�g�\��;�N6h��/��<-l,�Z����[\*�o��xpu�����[w�3����j6@d~Z����x'<uֺkN͙�!�۴���T�7�ͅwI�NnD�u�������u��|���e`��u�k�c�c���<��D�޹�s�(F`tN+������#'�(��)�8��P*�������Y��*���� x����v�\L�P��vn��B�re1����X9ǡfA����*�|k�A.��$G�tsFu �s�73-T����l�Ŵ&��bCy@���&#T�<��M4�@3����E@x�x�xQ�?:9��rj�&C���v��tŘ�kWGD]IЎ�l�ˉ;5�,
x�*L�i���	��.�M�(��F�`�Dk�rr0��O��h�^��+���� s+?Ј-��M���U�7<��]����or��Әa�:���Z"sA�RU����y��]6�U��}UZ�gy�LO8�)��,��4?�O��o��RwГJ\a�\���AK+H����ǝ`(���60s��IS�3w�F|������[�uⲖ3���U�@U��py�]��J��V�c3Y	���[L���c�nw��un1�v`#�m1�b����^��0��1�'O����
F��X|�!߀ok�b�1�� �ځRs�����y\����C�}�@����:�DZ��B������0^�۶E���V����:�����;�1�ӱ¥�)�H�!U} }���7�N�g�m���;[��<�ڲ8G�
b;8h�y:��c��� 4e�}>g��,~�KX
�JI^���v�V�xL��!D�:����� z�#�f����Q"eg�ANEh���~�K�V���}Ҹ1*v����6�ǜ���N�a��MW���"���|9u �S~��V���f��nL��{��}`�o�8m8Vr���)����r���A1������.�tGHȓ�x@)�N/�*����^B�ts�s���QH�f�]p����5<���'Ӿ���}�=镻��=�Ʈ����C"���|@�U�3�S��DlG�� ����zм=��
-���yr)�,�!46ʂ�G��	Te�)��if�m	sG+�����������q�=�5 `R��4p���	oN�����l!�n/�����*������T1�i���8-`��{n�x�ؾ�ي�h	3S��9
�?2��.��R�:��T�Rz�]u"I7t�9}[|� ;���ë������mK/���[���"_�%(1���s��{ �6K=�2������t,40o����=*��д����=�u�}��nD#`8�������Foz���.���~��P�I2!��J�VV��;9W���E���*�U1gE�Fǩ~<�a<�W�z�E ���&Qq�nQ9ju��_N&U��X��\��K��;��R�4�HM�����ߋ�  y<�yx��ki��k���_��`�{�zt�P���҉J�@I�6�������7��)z�O���}��z��ax���(q��&D䮲�vZn��`�U�%\(��q���]���7��h��V�8��U 5�J�b��(�.dn{�08*[gGJT�͗�0���H����+Ձ�3��l��v�m�UH����!�f�}N��a�z�'(s��N�^����=q&��06�P���CQبc�S���6U�(�L?Jd�-G\��m��x �W��� ]]�ˠP;�^��Z��䉛-��V%��B����Ѫ-x�Vڳ�/�9,8�l�.+�K2�F�̙F�v�8�р7LJ2�B�4 r�n�����M�����k&��4���f������蔷;Q�x��wJM�Yf���<0o 1�AvQ^c��%-�(�T�.�^w]�:\ƌs���2��Gy�/,�X�Dt9� ���9���e�vƕt߰�a�tb���XյX��|�]|���
k*3O�/[lQ��DH��7F2@�����X*��X)�T<��V��"i�KU�w�5xH��kP�c��͛�SE{N�A��fXed������zc��i��X�<8I�T|��*g�8����
p�mᨣœN����3�T��R��>Q<7~�kw����q��ٻbp�SeE�fS\H��M��2栏���� ��/1�}&�?M(��������Ǽ��gk�i�����Ob��W%l[}����"4P��w(k6�\m���9��>�tE���,�@j/A�޴�x�*��G�Fثn$���*,���=��D0��4�.`��(#��N�Hb�m�Bl���۫�����3�����J�R�S�A"`K�)��Q�u��__��YuC�Ǌ�s� ���1�x�<аצ�+y�F�
����J�*W���(��F;��%���DQ>��EP���Ӿ�?:��{�ï�#��D����=��y�?<�#ݩ���_|M��{̜��:>!�Y�L��L��!-�,�O����w:ӜQ�Dzd���RCM��x�c��!3i&�N��ed$�ױ�á�oU���vt��i&Dt���+��9_��j�QA&hk?�[B?�X�ۍ���M�!9 �����H
!�F{:��w�WC����j�]�գb����|�D��hB���FQ�RH��� ��;���_%�sG��I^�F �k��lW��:U ���* �z1���5�Y�&�_��П!f���d~TtBr;3�����Ik�i3�D������> ����`�tU�1u�6o�>u�&����ג���̈���B9��IA���h�ð�O�M3rAo��Fg��h�0�Ka�u0w������)5����OaTC�&�?d�qΰ�7�	g�ӑ��/JC����[�n,%؟oqE�xq��>�RS=���׻�#�|KUVz��9q��KԵo��Cf]hд����k��'7�L�>/e�Ehd�C��{���V��`����.�Y��,j�2�"us��U�@ݚ�܇}㪁���ӂ��� ��{����I����� ���)�����s���j_kO�"�!k����;����l��~�V��kY�u0�&o�m��S��1���~q�ep�b��B��5r��@�NE0�ޠ�K�(��ң�+���?�u3+E��N�p���Ʒ�'�gd��R�Ճ�y7��-q����7ca��������>��c��vJ�W��g��|}Ig9�����y��<���gS|��=����и���u��	���!�;j)�$+���M�%�jϽ6���E�͋������#�Ibr�F4�I���D�v  C��7`�R��3��=�x���jtߒ���?�DÖ i=�s���eh�a��r΃K��TV
 D=<h"d������$��b��yL��­:��˓���zʕ��Y���� �Y���fkԅ[�a�ګ�t�b���%��nl��5���@��U?g0�>g0�Z�(>C��wB�
�7b����PF�/����;G�>!hy/{7:�W��/sʟ:�
����b�-9�3��z,̩ݔ����5� #���w?���8�u^�2�w3'0�(��ا:p�y��p��5�uܭ[�B��c� U���T���A�,��ht#Ԕ���P7�tmB�wQI��`.K2J���%��O�e�寃y�\y��v)�Z�ž!w]�=}aVZ��d/�&��m69O��Uw�5�I���)�%J��y ��M�~<�;�M�e�C�I^"��$y�v�>���I��t�h �b���O�l�[NAYH[s �`�G�j���	�0~���yV�A���#'jmjZ�]1I�d��{�)�@�5;A��6��AMDw���#���\Ę\�Dd�(oV�sHy'LN?-O"�nd���sL��r��Hٟ�'J���Z��0��
AWQ5 ā��#b�Qe��fީ��O�+P��ib�W&��ào�39�S�S+۰����iǍEW���fҸ�s��7�o�H�;�<�q�~��� 70�,
��%��.[늏��P}t�D��8���^Vo��ܥ�e�o-�DT��P��j���b:�j�")pa�G��ڔ��&��/48����͢g�[A��<���j�GI�D�\H�~*Z9�m=���J�'d���$\��ʠ
唃$����>Q��@��{6�^��ۻ7�f�k�i�_�	%)��w�K���x�Fě\�`X�{L�7����J�W�|�W�/G�� `�jE�e���]����	�x����hB�"�`v8u�lj*�x0PTP�V�B󯫰hS���Zzi�̇����|��E�p����k1��.L�nju�T�耺�6 ���� �����$�O��m1Y�\�T��i��J���_0R5=L1o�Y��A�ڈ�҃�8�=A2����Q���Ch%�jT�W���s�����N,�G+㼻¿cP�H���Z��%�� #/�=\�q�#o)�k#�[���i�(rH�{�~�
�2�6�~VQ�#��-���Q-u�����^J�4����l�g:)�k5�YޥnC���=fQ��/Xm2�%C���*On�l�����f̄Zxy�qF���q�`���@�R�-0@��x��\��Q�f�:M֭4%w1��K����)�{�W.��H�����y�/� �Q*+�RG=<�'][���9�B�(;�q��3�>��q<�
��r}�_	"P�h��`��ꍵ��l�����U��zȏ�x���1�Rt�ֽ����OU,0���1�7a�/3K�6��6yU헒t�1�0o��60���I3����hqbA�~�'7P �#����b��w6��-�V��h�*�$f�"��JV��d/Kkڜ^Jw�S�m�a[�%�ӫT�r��O��?6�d��I2�}S�9,d3+�o�(˲���KƯg����8�M(
ek������� f(���1�_-:��?��ÝW۳����Q~@�]6��pH��L,&_|]�8�,��F�@J�g�ܴO��Ea1IW��˂AJ,~o��q��1�`��[�{�蓁n`=X�fx��|@feM]غY>@�KZ�Ȅ5^Ԑ����`y�j�OX'�>鄢�
�Hۃ�=���T��A͔��Z�_��K���B�¾\��	���w�X���\|�VO��5����H�+�,�N���ATywz(��g(<�����q�5+Z/]�"ִ��� {	��;�3�[�v���E���wݪe݅� 0.	��ʋ��>�t�����w8r�Z%�}1bZ�ӼIƠV��m->>�l��V4���3�᱗x�2��W�U�"�#1��1ݫd�wޢƖ��f��S�K�g'�z1�������pȭQ�QD҅�w�Q2%������"-~_A]u��KãsY�8T�Bk��)]��-&��4\觞��F�
`�V/=�aOl���@K����("�ļT�IC �׻(�	�J�3�Hvŵ|房T��o �3�����	5��7��Y⫄l��H�F^�P���Ϭ9��|��cz����*Hx_�?Z�g)>� )��R�3��:��;m��֤N7[]e/�old�Z�o����!�����4�R&��Y��I	 1�Yr�0w��e@�*8���m/�j��2�r]w���Un�,8�f�i���w�	��/
l�5P.�m��C2C�t$�0f��ӡ�ʊn�w^n���^�� ��^�]�K�}&+������n�5^�6���Ty���cB�w^;osq'd>�߯�HLp�-`��a
���"�/i�>�0�.�ۥ�?���Q:ј���j���!N��#Z-O.c��\��>�
�֎��m��	Dt"��"׹��r9 �D�ڐ'w���P9��+g�Ƣ��ע���PhC�֨7&��V��m`��ڦt�燛��L�TGt�F,��=i�e0�E���{��b��B�7gUBJ����I
��U���:�m |6�Ai>���߅�`@���W$�x{RgF���[BO2�Iָg{����ے�W��v�ٕ��5�+&�JK�
ǜ$�&�7�o���3U���[~x΁]�P��y�<�P�-ъ]�Ey��Z90����O�x����fYU����G���J��m��,�'K�:F)뙩�(�k���.?��=��)Pڢ}�b����\�)���b�.��	�Ap(�ٷ��
��'j��l������K�{��m�a'��`g��Iˋ�s#�=�����%�D2[з��̇<m�Įb��N��|p�N������pYÉs"ӅK�g@D*c21�=L_"��{��u]���_g���=�P_WG`d- �I�<����<�}�nhDV�V'���O"�tk����&�Ai�pZ|7i3�"X������)�.�cv�<_��1�>X���%NY@���Tf���a޳0{� ��x��#ivÂ��w��H�d�QU�'q�v7@�v	e����eC.�#��J.��~Ac��wwlNoO����P��W}r�d�4�� b���*���z��3m�8�����r���� �v"P��u�ܲ����&�j�C��\L�ANjF�z�Hc��d��C2%,U�I�Q������7E<�3�n��.4�R%v���V՗��l�\u�x�7[�N�A�#��E0#Ynj�t��~�k�C&V � �v��,��!�Uޠp��;�e6�>��u�@�Y#�&�\,F{$�V��:�v�9���ݪ!��;�*\J��|�x�O!+���59 1Ѐ�e�њ��vnO���mܦ�7��s5z��K�Y�_T��~���:G1X(��{�� ��H��JE��\P+��2�5����bu���XbnO�+��B~���3�Tz���h�p&�����lV���Wcn���cM7��g������E�������6�{Ш4A��0'�r�^�8Ku���?��hz�C�9NZ�#��Fbĵ�h����.��KM@jw����>&�)�Mp �\�x�d%NPe�ޔ�����X�@���K��tz�B�.�L���	Ka�
ZL ��Ck�E�鈷�NO�3;m�{6�}߼�9�=	@Z
�����CrRF:,S9���ҿ!Cn�E�S���+�^MD&���o�j�@�ū�_�h]@��Cv�YZɭ�J��P4�O�ڛ]*�wE�=�~&�D�d�JV�������K�@1(���haYk��W[G�pk�=��RG'^��^����b ��E���C�. T�5�F�M�n��\1�'2�j90���B��@�|�������Pm�$w�~3�L3o�0���p�gc�4/t�Ē-f�6Ɇg[��
�����Z>T�B@re����I$%��I��ʑe�\�N��C�&�ճ&Oe�n�T��E&�����P<��Ƃ�l�P��(�h�X썿�@.P?��6���[B�*˛�X2����e�}8�wH��bP��^ ^
�0�dH�M_��m+���t���
Hw����7å~��S������m%�%,F\��޶ͯ�w����E��޶��~��G�Xk4w U��E�+�U�\�(�L�\qg�aإHJ �,r8w}�^��'�1L���ӹ�A$����Sc�� y�����N;5���k�Q>����� ��Pl�1�a�J��YDd��w�s3QWd!v�fï��2r��GYi2���u�`��;��N�ǔ?�lP�Г�y���'���t݀se��h{W�����Bп������)�}i���#vr��Xw�P��읋�9O�o��_��FQ
�/��'��$���j#����Y�
t��p�E;�p��u����͒�ڒDU�F1�YN�=/@Gy��X�!�.��~a��M�T	IǄD��OB�`�Ȯ3Z����`JZ���ܪ���/6$_ $܂��Q���-��i�aѩ�p����閥���S����8O0�E�/E���@��B:�:G�Y�Q�+"��EF��u�5>�5ij�r��kTr�� c��}�5���>��K=�4�ck�.��x����G@-'kA
�V��?�_c�1����9lJ�m�"F��{��t�?\��zT�*����Py�!F�Ϫ���3��,�~��Hc+�����M��5�0�|Ǿ����:I�&/�\@÷{�[.��7\ΐN�c�z��M�n�FŽ+�db��� ��C�+�F�B	ڪ�����o&�8�	��J�w�e���5�mN2��qɆ�^^�R����r]�x�,�}����`x�?�����r��|S?iUoP*�S����Nf.�Ǐ��/�������$y��P>�&8�>�Y��;0��L��ܬ���c"}!jz}~
�5�w�[`�Q�= ��I&�����D�,�݋�BYK]��v�A�w�@��;�"h�cHĈ6�`7�\��7��ۣ�O˞YGT�����`�ٹ�OIf����c�5w���sg�#�Gp	�U�����R��{�[h֓�,l�m���uTۉ$�(�t81-��� |m���롞�5�o�BYk�%+|Iˉ��ƪU�Y�������NM�+P��*��5���{~4&T��	X�#(OL		��5���HD��Ǭ�K)���Y�8�lv"Jn�@j �'x�|���L�jP:�zĮb�n�s]��B@�e��Ш���:��9����x���h�n`��	�{��ɧhS�O$�r��DD�g:��A~I��6C��F������e�Z[�?î��N=����N���l�K�Nr�uG�i���cLW�].����Y�9��j�I���t�i� #bK��K�� ���:�����Qr�����v^�ֳH+=,\�I����Y���������&O�岇���t���-5A(X�ǻ�o@���uV��	��}����Z��ٙ���9�%+�")|�QZ���z��I͍�Ck/0����$[��qZě�Qek�j��h�F��(�X��0n�)�'�p2�~�ܓ����,��զ驟jO.�bi�Y�ZX#���[0���EһW���j+�_��L�T���︯�i�:����IץN��`x�W�����,=����ؕC��	 Įles�u��5Q)��]���a'� ,"�4;�E��7��d���j�F+��]�:�D`�t�@:x����!�wm��d��h�m��,�O� 	�Q��W<�zwH����i��){B���:Ԡ���4�1�e^�~T[�	=��T���Eg�rJ�ndh\~yܡ�7��U���x��6t/c!Y�4@=��}��6��F������脱F�xV�%�O�[/|M0OƐLf�����RYK��^�"��w�Y�F�v^�g�Yc��������M�W�N�
1	�Z5�.���Ů���4�w������~f���ͺ@���W��H�x�Eeѫ�#���my�>���ǁ �������B��2�'%H��q�����Y5����&�XM&J�I�P��|�V���*4�ɝ�_��Z�Ç�s��t�ݦl�'�ֳ�i�V�|�\���zr���1rio�d�U��Io�L
�u����6�?Ie܋��#gPF�U��C���Kߨ%��'���~i駂����_Ԍ��w�OO�
�.����,?c�I\A8���)�}���3
Ω�z0�8�Xõ�.��za�{^o��@�rHr�Vn?�U��a�����]�8��>£����k�Y+�%t��&ا�ǚO��ad�L��!��$�=�6B���8��Ow�� vY�[ƃɞژ�e;Z�Ҫrr�f�C��^I\������E�~G���v�<
�f*ͦU��8�fw�x�=���[�眧����8��9,��U$_���p*�Ǝ$3U0ϤB��#�S�M��#ٺ9h����'*�?\9`;ll����N�yTJ����!Կ o��J[�t��0��~[������w�����~����`�g�eN�T#�د�m0��E�
&Tνu�s����������Qw������w_=��h��  ;Ҏ�^@@�7���QjwJ�����������!-W�$hж�G/"�[����Ș�������Z���]�6�x�=�u��(=1��'�pѥ�`QҊ�~���mӧ!XޘVRG9��T��%����<�'ta���nu9lˤX=�ԑ�viS���(tU� 	��g���VmVy<3R�8�3�Ha�S0on�-e��[��D��!M���������m����"��E�#)K�>�GД0��
�j���W��{�C��B�mH� �T�d/$��R�������z��֤�O�I�t��!=��� kI����`^��Oe���={+�	z���q.҂�p����c'���gyXi(�[g8M�A��R��	�
�f��p��7{ȘǸ�%�|���Q�]T ��(y�`�&+����Zy�,�?�^�CfFą(K�*������ަ&��rz,�:+/^���{!���`�6�	���"�)ѷ����m�Z5�0ݔ����Gۊw�Z����@
N��q����x�"��r��±p��)�_W��Dt8��`���kUA��e���!e/SN�2��O1�Y}f|��0=Cd�g=R=����ߜ�C��� �|��,S����������{Np�p"ރ������
i0�=��2�6���L��IX1_�s�L�Y�X�J���㮵�>�$�)^�D~�h��U�%qXo�p��o��|Ԭ�A����Hq2	I��32h��9e�+sѾ����#]tb���/�f6<�{<?U�d������G��1�����K�ӥ%�UTVM��\�ZY-n�/ۆ�k�ȑ�3�w�) ����+bI���ֺ��I��XO�l#M��f����<VSć�>\n+I��5�6��R�	`$����j:���������+�C�rٿ��Sk"�@��N�w�q��_,R>�-G&�+�A��#�߄nٱ�E{'��
�PblO08���c *Y�ɪeV)h�w�ڒ�M�c�x;vN���X`�,�~%�w-�����ir�.j�������Y���ڭ��$��֫B�����y�9�ӵj�"&�μ����YOe��	����Ux�Wt���[�
@���^�72������VZs/~���M��2��=��\o��ìߔNCY���P��loI��G;����<\/�'3����5<�h�����"��H{ϫi۴i@�9I�������^�i.�W�~�F#y�9-$ ��sH
h��*�_�9��|z=��){y����IҎ�BVb6yt�ǌ�"�}1����VƷ�%�i�K=����vq�8��B���ܥ7:Z1�\���<�D�Ҫ#`��=����r÷��E����@˹�^=��fm�[F��P�ʿ����0Đ&�	ѹ���@ݹ���V���� �V��yHŃ�� ���6V�M.�X8(rC �Y�כ�@���eV�Q�8��b��n	��g ���`Eό�����Lm�l!����y�ݧN#BM}��S�{�G���}�E�[���=L�n�i�Nu~�X��7���7�E�����ؾ�:`����һ���'������O_���œ	�y��8"�5\��Hۅ2&7� ��� ��^�P�7UD�zX)eI��1�,U��|i3�0ۥA��+��v�q͡���^��4��c���S�j�`C���4/�]��E����@h��Vw��E��d��("��o�C�Q��B#�gP�� &}������q��G��4	�8|ƽ��s����:�^���4T����8�0X�	�b9[�K6��"Yj�S+�J��'��9�䟗�b�z�O��t1�LYI��0�B,%j"�-e�HI�g��U���%��u>⋽Թ�*���p'#@��T�O�|�F��؞]�_��;J����1�z]C��,��7�5��VC����.uP����=�����Б;Yܢ����鰱g}�~�]�BY�v}ba6X|u�.���VE��&���ط�?� �k�����Ԏ��H|���DU����q�/���Q�#��i�h>�lQJί���iOm�'��m��Z�t��p��Gze�H���&�z�Ѥl��;&ѕ��wf �99����B����e��9ɘ��t����s5e����ae�Xt�
�� ��(���Y���W�U����^��7^l~�C	:��c��Hk����@O8�a2�m,7�?�b���r�H��(7x���O�r��V�T9N�1�������{��6��m���sP������v<�@%��137�����M�Uw�\5h���Nτ�"~���egA�� ���NԋG��!�ܲ >sx
�F�Ew�8R��{�� �0S7��i��� �	��G�2*�p�tY���p��p催3���3��|q
�˙������ŋ�y{�����w�}�`��i���h���E��wqe	�����>te.x>ݬVZ�&���uU0��_4m��njRܛ��B���V����}������!1+�ɑ��p����Ew��R g�����84Q��3�JJ%����3�ۘ]̀��ʛ��Ҧ���9������\����j�t�Z�Bu���,�̍��5��1���4a$����Ȇ��c+�f��&�}�r�hj�������v��e�A^g�/��-k�-3�3	�� ����i� .R�P��D�'9�:��h�u�:5h I�����XH���)��
�'��I��ɳp:���lm�?l\��f��2vz�%h$c+{_��d� ;2(��ZWr�TV�Te��}���c�$Ҋn�a�0	R_WR@��������"l
W���L�2������ܨ���:�dv��y�8*��nU/%*b��"��/Z]�"o��"���3�N��y�%eu@#8���&�3����zؗ۠yT�!��P�[HR�>u�3�\q�$��I�ʛ�3�'�(^)発�7W�<-<���2���[��r����Sa��+��̖�s�xT
���m�E��t���QL4!����FHap�c�+�g�j�*��9rD�aGЅ��+��:_\*��y[��9}L���CM����y�iɃ�x�;,���?�����&,�_��K��_��"�u��zz��W������18ב�	�)����_Tw�,@�49d!e�rOX��2�����^�B�����0CMru��O�R�i$3Xl��%�q�	p��m���c{a�b�����V)d?շ9�L�#�`r&�~ڈ�"�!��������.+h�ɴ����V����Ɉ}6�����CQ�jg�P*���=;{*�Ke
'�7�Iѫ~�{���j�4��O���k��L�K4���%%RƯ�4X+�H-w_P�s�9��½=_�mn5�����	�����g�g���YW��q��g��Ӥ-.2�[�����xSaDt�]���G��A����_��*�b�Z���7 ���ї�Փ�5��Φ�>���a���fb��毟J���J��aw���E���s羔9,;��a�6�'LB7��_F��c߯I��<�]�>9jzpך�w�<~�(�ANH|3�z�vY��z��:�W���4��h�])b�-������)L]xn�F�&l��I��rU3)�L��V���q1�f>��qN�*Vg�K(&���$Oa���ͽ[�)�i;�0��}� B;	�:�Q�6�^fD  ���Z�
X,�D����{֞2� ����z�5ǏY��,QZ�X�!&ؚmi~m����Z�hS�����
]>�f9Y����[dJ�X�`��u���r����}�=_���AbHy�،��`<fG�w[��lx��g�[ŖE�+9�&� k�l vad_!���'��
������ŧ�<��S�ON>E$�6W' h�.��=ݐ�Я
M�(���i�������{��J�:���6��iv�#�����U=�k���8��B�)#�7�oSY�L�D1�$v��P���{���著^|	������%�[��o���#��
T�5���A���6�Y��� �v�Z��*yQ���Y-f/OQ�wٵǁiv�+sGG�x*��a�2�KVA��K�&TeX�(��m�s��榢/���l�}�0�:(C�@{��̟��D�T�?晾�=
����^Ӿz
����[��!��@8�7x9�� �C:?���4L`��iE��������~S������?��'�3\L�v\!w�t�����@ zxy>��TP��K�P�=�5�3�G�Q}�Ӧ�	'�H�uZ@�O]�0����������j���/h�H�`����/���w�*h��n��ra�C �r�Z~���@%VT�^L�}_�Jܯ�+��nД���{��%`�?l���9Pq��t�3�^פ�m{��w������dKUډ��o���>�bf�C���-�c�
���C�(ݏn��3�����F(��L��U.���s՜��w�����z���(]l�����i��kA<0t.�&����Rە�������y}&N>a��`�[�D�r|*�{���<�_B��a�:�6��e�}#U��}w3t�`W�O}z�D޼��F(�nQ~P�әN�x;9�o�Cl�~U�%�	�T��[��v��V��2�u5�|Y��t�.���K�4�!�T�sI����S��59���O�h� ���PY���}��p��$��f~W����$B�_M�A&�*i@���Hm����}IlZ��T��7�yA�#?mgQK�+�Y[��*$B��� '��e�[�1ݸ���z�X;��ݭT<�]��g��4ڳ}(u[DĄ}��o@pD�̟x*�3��K�V֋B-�/ʩ�����j��l�KB�.�>�>�4<:���O��V�r��*! 3��qf�5��x5�[��JI���
�I����b��pR���lU��A��Y/.�&������c��W��izj�9�*/p�MUe����|��:���%�����K)�aQ ZB�`� �7�������+������=���2q���l��WJ�!��⼸���v�����fc�#P�_�?B�����i��j
Z��e�kIV�7�@G|��:E
]�^g��eK���dT��9o�S�x�st�'O-ܠ��b��2(�r ټ����A�4�gJ8�	�?�Y�É�H���4��5�o B>�9��?mԼ����8M?�HuY3�`�������/�o��Qj��J~)���/�����1�G��wI�M�c��T�>�Y�� ���Z�|%�t���WG�~�Jdꉧ�	��c�j,h2
l[�7��&l������ىuր�=�/�S]�1
�`4_��y:(�}�q�:��h����	�X����P0ħցt;��u+\q�Ѩ5kR;m����ae<h�;؞8~vy����4����Q;�ϼŅ�U��8��m�˰� ��`���!�,�۪c䘀x��Ƣ+��B�+lJ+�*�c��gɠ� ��e$�n�G�^u����HU;xlQ�D`���p��<`��L�㏶��_,����x��>�9�#e}�댄 ��uui�֝m�7@�C���n��VM\;��۪���bi��P�lyA�\x���K??�P����Db�l�J����H�;�.�O����꘮q�^� A־E��	N�3%	�W�\L�g����k��C�8ø��w��e_�i���g����=��w�^mxz��ŋ��_���1䊅Fk�{E��;V��8��>���lZI7��$���p�t���Y�;6���3���ߙ�oY�d�����3ϴ%a!&��3ԇx<_-P�R7.kVc�G���q�'������Jfa⼕	��Z{1��^èsL�5��?X]+�sA=m���������}mi��
�����$����?�SsA[9��p%0>��o�^�f���?R�
�Y`w�'�ظb���
����̢MH.�W1�4D�K�Q (%�#�B�#%�����n���e�7S/@����;Y9׎{��Cx���(�}�|������>���.ް�Eϡӳ�HL�A��5bщ����˩飴6Т�o�$ԯ)˘P�8����- 5��1��|�[tq���+�K�)�ZJ��u�y��H0
�w����0��t��IO֮��_�`%F��+���Ƹ�B�Z��e(5�����ר�����s:���"\����u��=�cu�l�i���$��O��^��"ŮA�8� #�Fj�M���Unj���ڳ��^���1o���I}e�{H`޷ �]}ҏ�;�����!��Q����cdZ�]��}����G�)��zQ�|)���{�r�k�!��ٗ����{��t&P��6��[i�P����t�E`��BY�3Q�Di���M�Cv��41�\���ex �f�����Z?TU�=�~�[��3M��$��([S�W�,�FB�h	J�ȭ�����s
7��;�@WWq�F��k~@FG�Q����v����PA|�s0oo6��ZwZ��l=���y�ӳ��#��q��ytLo�����_,�� ��UI��V�4PP���n���6k=br��v��&G#%���]�֖��zx� �Mμ<S%@������M'"]����B�N,x�B����Ck�)�'�X�A�+�u����;���U=U}a�vm�K���t�=����o��_�E��4�A�xQz�%�� ���A�.�\�<I�����V��3��k�+�	���v������G�@QȸS(�>x$�x�C�X,tΜ��4�8����+��k�K�ٺ�����^=d=u���ik�I�Y��6@l��m�H��d���s:C����[�o��C�;�Ԑ�6�:�����V^Vӟ��
ݾ(��QȒ���0�X�ݼxg���H)��}�L�V�=v̨��H؉q����#����~�O�O1���ɤ�'���%�e��^�or��7 ���>�Cl�'�9��4\*9��+��h�dO}]{u>����>�oS�D�&&����!?7�UklL:#\<��|K�@+ � ���u-�4<�I3#0���1��������Pp�}�A�G2�0̳���a�?14R%-���z�,<t�8�I���@��<EnY�U���P#@ӻ��.�p�`���1YܔM2���[!Ӳ'�zKL��Sr�Or�!����/�[3;YVs|�x�+�K^�"3�:4˩x"���We���)�?B����2�����yg�Ođj�(@~�F�P�X��r};8C�xY'6-\�X���v&Pm_�Վ�0�ȶ@踨�S�y!�l�0��n^Ӓ�ՠ�:�/�u��!2G�;H���ך~��t��K̎�Ǎbt,9�UlH'2y�Hs\��`�����=wi���ߊ�Qh�vbF�"�1�����j-�4�trBtx���Q%������[$��}d�X��4�,�O�LB�6E�ٵ�0�ٔ�;84%~Ɩv�g�r��
�y�z���}��FZ�C Ε�����rc�
+�&�X��,�yV���S)�3�kj���&�t�d[�@�}���M����5����!��`��<_��'����]u�#�8�Ff�F�x�Z��6	�j�P`�G�Bj�9TT�1IN���I�,�M�X.��K�?�`�o�����\&����C�:�[��&W����tA��!d�2�C팲E� i�4P���
��䋆.<Jy)`Vj�.X�1@s(���Q�E�(��޵�,CK��m��#�,P��>��CR��d���9�����9ۄi�T���k�����8��K?W�n(����+���$~+}�E��83?�ּu��(�2���<��`{(z���ud�ɶ؍�P�Je�_Rw(M��ք�Ѓ�<�Y����w��M+�k*�V!��;@u�E�2�}o,���zLO��ss�P�r�~��n�u(��Ι�D���D2����ޑ
�k�k��E�k��\��ݓ\"j&�M]�L���
Ͼ*��(�Q:�Y��X����)��fL�2�@��e��r�eE�Ǡ湎�u�����!��C��)î��_��b��	�j��Mr�f���H�?�i�q�V�<����W'!�����)��P�I���L�2=T�I���ʃ��dDo���������{�t�D4�?:����Ύz�i)G�/y���U�������58��N�LtDxGq]t(˜"� JS�[7�,�mN���	�Tb �����{�	@�97^X4]o�]j�ԗ:�B��
s�OdJZ��lMHǶ�����xqx[gϴg�����b��Y�^�N�3�k!�H/�P���T�k"Ft�]��~ee{"釺2�ԙ��J��0}��Pi�l�u��m���J��9t?o�be�\<��G�� d�1����7k��kE���1??�3�B2c�y�2�=O�@"�P~�Jh=�� ��ph 2��J���Ow7X�����,ƈ��MT<����9!9���V\M5v;"#D'�딷��ǯJ��RZ��!%{��Лb��e��	)�?�b���^^SwF�M���r��u�;RI�UzlP�W�C҈�p	%���xe�����T�9Zx�3�\��-� ����Zjb�
�Ho��"�{�6b�Nar�\��(o���-!�"�9���$�R���暘hH4�#��D��)��j�;r�w��w���-}T}{c�3[�I5|P�H���������}�C��p*L�������S��Ǟ�$]p�	鰇Y�A���Y#U�\�/�_6�������D�8Ɂ��N������2O�':�)l�EQ��T� S'�Pb��!���ҍs��^N����U��s��SS��y�_�Zx"p�S���h^���K*�G�Qл(�P���
qrv�,�f��6��C�$�,L��W@�o���MW9l�)�����N�-�w����lyh��%����:���s[cZS�T HE����ƌ���l|\��;�7:�n[7*k��@�6ҢJz��Y�@P5L�3�֮���ϾN��ejH�d~$ξ_����f�0<���ӫ.�5�b�/LX�^D��1�b���[��GWe7�޻J�L���$EF��w9:##����̳rg���Y鹌Uع��ǰ�O��x8�IV��)������^ƉcF�#�;���n�t)�wYFLx��?�ۚߴ�Y�ńGAN0ʊ8F�B;�U��J]} ��)B~��X� O��E^��.m.����т����NѬ%?6�qx�d��#0�Teq|wA��8u���6���-=�9��������~{�����R�h�e�L����Z_�-6��,�o���Qm�w��6��kE�g��E�9����h.���R��g)N	D��|l;T��Gԟ�*�g6��w��cw�`Q8+|H[ޢA���ѳĒ��6��pg�q�c�9Z�h����^f(�ldG��e�
';��>8�����Tux%��r�~ġf����%c�Tx���{��@��"?�Fav���r��f&�aY�h�*���Kg�nsNn�zr_�?uh�g���nY����ғ��~\٨�z�p�5'�!���Ɲ��wE�]B30�QH�N��L�Q�S$��!�[�(=z�y�Fh�F�~�q����-��ݛW熬�5&���;L����F9��};C�􀹕�ތ,�p}��%G��0�zSy?-��~:��jj��{�h���7�
������{��Y�\����ԁ�Qg~-`ttf����5��M��c�
u���
�H�~�!�Y��;��dZ!�3G�~�H�t齂��	T@�eN����E���fFj�FW�������۞P
��ceZ8�LUT{���`/n�S��B�����Vq`�a%�E�S}̨J~���e�����4ة!PM^�����������Wg78�2�ꑪ���p�����ݢIdܳ����[9���^��ֳ�ݦ#���g�6:[��Uߤ��i�H��Pl:��"�*
�c]ޞ����
�Y?��j:G�"7��L�� ���)}Ŭ��ȹ����.�̳J�-�tĞ����!`�M��*�
��7E�{Uњ�vՒN5�n���&T��*yX����q��P8��nIS�����TI���t�=#�/��_�D�?y������"��տ�\�؅�����0�qQ��;q_���Вڏ?��l�q�L��$h�Q��Ru��ߝ�G��EN J\��i|��X�������3���7g�B�i}�E$���h���H� �MŚN#��J}�+#�q�@3��Z\��TB ���⎾�)��8Be���6�/8ٙ���W��^�8$��3�j�a�`�G|�������u�z%H��W"˵�k�&��e�����<l�c��>��������#['z\�?�n:LY��x>︥��{2�����n����zm�h�y5AݶB|2!s�SQ�C�Es�&�&�Ϟ�o�{���r��ڑ=�c��s�qjC����K��w�����uZ��1���쌂,#�� ӛU�n�x��G����7	?
���"��4k��S������0��8�}z�xmhg#UqC�=A@<�v*�\���j����j�{ �g�L�4�F����e���`sq�Y!�Jb!^{���6�>"I�VBg�D �P�U���?���u-����MKi��6���%Ƨ��h���$  �� [`#�H������u����Al�)9�Fn�n˾-r��`�u'kC�� ��nj'�[��~�2����h��G�Ѕ�r1+rO�Ǖ)qʵ�'��	O��PV�cUр�m�Q�_��9~�����+��fR���(����'Q��Kר�"6��c�#�@#����l�\ѭ �	�3U�oc�w�@�L����"Co�S���?�2����H����9j*X-|z9r�`�EH�M���t
����T��)�a��Stz�;<���)ow+L���c&�j����b&���ş�F�m[)��!�x]���K��5�"KhO�&d�{'X/T���(�^lB�3n=X�KC�y�k����?aN(��PL�{�c��h����O�v&DX�k�}j^�������G��Z��3f@H��z�����<�n����P���>���)ڰ�V���Q�������?')��KN�T��jׅ�y�њ�C�L���I��,?n����s��ҍh�k��._��nlľ@�9����Y��5hd�`i.$J�����
tV5�_.�{/+���nB�P-��M:>�����5D�_�|=���iV�'�ϼ��7��"ٺ���
=j�?���� �W���)��zA��H�
�}�E�ˠA=�_�������$�����3OI���rj����
&/���JZJ�Lk���sc<��/����Pߞ�3c�>�Y6��^�G��?\��=�U����ݹsw��CY<� �:�Y��C1���2T�	<\u�w[
薼���eOI���~� ��;�Q����A���r�ڬ/�+WHCE��|�JI�	�e��P�#�;!0�1�]���y����ٱ��y7<Ī��˵�����|q��:%�.���q1fm+�O2�h��JZw ;D0��zA��L>q,�,�@[&�ۄ��4�Wsr��Q����y��y�2�7E�@�Z�Bc��w�I�����E�ڒֿ� �IɎ���)Ba͘�Q�g�3X|�]f&��8G�^[��Z�(q��wZ�p�1�#�	ScH�.�������9ݑ";����t.���i�9����5-��X���"������3��OC�^|��	 &�t��^��QCޭ婋f���%�#HHCDh�K���&�F�3�a�v�B���O)LJ����G���v�)w��ʔ!�V���l��W�V��~�$MI���Rp���@s�c*u�u��qN���g`eS��w�$�o��يU����>(��)��pn=�`o�?Y�Jq�f^|����*;�9��t�5c��k7����='��*�N%���<*�&��zl��9|�c�~��m�	��1ͩ���&��w���JC��nG�q�J�9�>�0&��:�\�ܣ6c<[��WSۨW�OO�~����U���6�׋-_m�6
d
KPo���n�6s۵�:�"�G�W�l}8�;d�h3�Γ���Z������>$c�xn�b��@�����7A�m��=��� b�w*@G�Xҵ���H�W�\�)'�m/�fԭ���(
�}�G�+�p�C����HAjK�dSiT�(�� �474g��7p8A}c���aO3��y�i���GF��ҸѠ�nQ^|�`��$�f�G��g���N́�3b[2�����X{�����D�Aq�C���9yR�[�^ҽAͤ��t��a��_�n���x?�)j�m�ҟD��(�+��$�{���oQb4��	q�A �u���F�� �Szas�W���p���E��A���V2y���W�^pU\�
�l�鑂��=_j�/	���`�ASpk����ǳ����&����J�UE�D�=��C��-\��sO���!toP0��4B��Q�	�>ן����1c�c�ȷq=:��ēw =X�$��D��B?V�4�u'�����qB2�[� �����[j��Y
�%'eۆg �泑:��ɀJ�����b�NOK�V����!��U�ڎ�L��(%^����#w�F:�5V�'�f&%�Yw�caqS�=d���V�y8F/�v>��2���~O����*��b��]��F,ޖ���Sf���0v�r�M���P���
��xV�E�Xp�ءo�p���FT�}u��#e�#Zx�]�<k(uA���u���$}B��$#��fM��o��h���o}Q�B?��33��8ݤ��|c&���#�S(�l�}�D�'¨��	�������O� &im����d�F�� ��!b�S�Ȳ~�*,���^)
�Q1���������o����Z�iJi�h<?��)�GW�}T�[2�)x��h��i�������v����g��#�+��~6���?�`�8�5?���٬ME�߮zq)�f��T+�8��c����({������6&��M>1ԡ�R���ĳ^=�:�@Ĵ*[F��4(4n��57؏C%��� ָ�2>�	::@�P���Om��O�%Ă((Q�����-F$���0Y����+�6ɉOݢ�9����0�I�tC
h�A�&���_�z��}T2��ݔ@���x����d.Q�U�M� B¿��_�E��N�;o\pg�@�.[r�w�6UZ�b�Z���)ϕ-����A�X����v�n���,��SX$�I�X�<�2�K��$o�7'l��fϾբ��L��	[!ʗ`�'������!)�qxv�P�cy����;�e;��U]]w���
~�e����b�-�Pd��UlL�f��l�g(�.��4#�{@䅣�4~`ﳂ����C;a1�uz�[��� v�JK�H#g�������BE15��]�`�{�`�I��6�������̂�9��ys���T��k��}ס�Ǻ�]1���Ҽf�����8�[Ss �^���Š��>k��<q����$�w��%��>z���������9��ye�p���p���L\i���T�z�xY(����������*^I����3�����X���e�.m�͖���Z��y&� ~���<���t�v�6t��v&_w��4���E�}�0n������팟-ۡ7 ��xտ�����e��bC��)��lM�Qf�.������k��ZE3+�T�K��v�/z?�v�b�^<"h��1��#k�=�����4U��$$>d@t@��&>`�Ֆ��l=sa��ܒ�� �o�˯ߎ8�.�xD%x�43����� a��̬.i~ �Bԕ�ݾaTR��Jv{ ^"iK�}�����P횯����c9������Z9'��\l�V��fκe��+O��0���NZ��[E
��2���@�L��׶I��Bx�ZvQ=��_iDq�Fd��G�ZI�R~9+���.E3ڍ��i���e#��i�8��q��B�d�,bM��<y��uk���ٓ���H���<������E�O�u95�����\dkaBCT�܃�@�25��f�.�ҟ(�%0��4lG=�{$��B7�����,��}k��~Æ�Gl?H{�{����1Am$�j��������O픖lity��>��l{!��J�hӮO!5��i58��纷O���kG��Ǵ�K_���/ !-:��ڠ�g� P�G`����?k�_k$I��Ğ,�0s'���šB����4ގ_�m��8���ɛj�Y���K���^���qY��/��(0c��u9�'S3��]_+^�<baZ���þ����p���{�j�(����oh�? �3^Tٜ��K����?+����e� �y�f��Z*�B�	}\����ק]��>��F�Y��f��g��=u?��t��8<��q��Vs5<ZH=�(̺�La3)��X$+�1���uN��ֻ��*���'؁}�O�k֫�v��3�1M�bR�t�`��B���lP�5d!K�O��aX����"��<��<(�a���Ɲh-�/�uO��6�!#���{�r@Mȫ�GL�Ga&�vR� V����\'mwH7�h��/�;u��g[�4�iȸW�8�J2a>�� �(ź1l�A(?�m�$eC��/z"���G���꾇�5D���(vY/`w�	t)6-v<.M[<��"E�2'����GM&>���%9v���^�&,�ڳ��Lg������qs����t��U7���-,S�~�ܵ2���'aO����r�<�t��k/vQ6����f��ֻ���lx�@��O��k-`�+
T�l�'�4���{��{���*�E8�Q!<�~�| �kN[��a�-&��_�ݨ{��S��7��
�� ��E��{�H"����v�DNҚ�qBZ�]��>��HX�<m����i�j��n�"�/R�u���������F/�l؝ �	>&���2������0�w�ιÂ�g:��=!Ś��q/I�Y_� �W�Z�pB�o3��������c IedѵWnE��,pa�w���0��*�<�ި�
�[Fǌf.r����j�u���S#t�W{I���Y���b8�w���<M���v`L�i�>��~���vJQ��-�e��� rbg�m�RLf=��(����u|ɞ�_��6!򙀱�	��ʬS��N��)�^���gs6B�s�M�0P�;Ə��M`�f�"Xo�,�|a��,�_��Ad�?w,��Y�v0��k�?L۰�6��Z��c<ȀܹS>s,DB\Ϛ�����㻛ʛ�C)�n��S3�S���D���i��M�.�h9
�_zK�'č��ˍ׼Pk�;6�L8ٯ���J��4>d��0y�Ƴ��;2}-�hځ�BH���{�C]ęV%W���;������{.����7���q֘�ߕ�W���a2D���{����?="�������-z��c�2N��������p:EA�9�4x�13��o'��rɇ����H@GYj�f3ѱ��/�R�H��O+%��a1��H,&*%�m��
��t^�p�D�ޥ�@Jq���jIFc�[�F�e��a�!L��g��]C���V�V/�Y�u��G����I�!
�QM�����r��ƍ�V��C�y�,�Q5q�V-�ӂ�:[aIij�mo�AR$�>jhbL��wQ0#��@�y�3�'zF0�:7��ڱȠ��a
(M	5U$Y��.s��)�a�F��s'�`���!�*g(b2W[���0`j1 ���wZ'RJ��P������OF�'�bIO�0�T�%J�r��.��<[y���L/� K��-އ�rHeg93GK�B����m���2%+ȫL�����y{��2���༃�o�����֜��(+rQ���6�4�ɓ�h7�ֲ'�I	��͛���p��Jf|2`�C8mO�/�hk�ƣ'��(��I}��Hڡ��3�rÊPc���c�mH7u
e�{��~�0�*]E)�!� �ɔ&��O/˽>�'N�جe�6QE��~���Sw8�C��K!��V�W̑��8�f��g�nv�ulxgԘP-y,�����gHދ\S������؈�� ���__�[���$!��?�\���@��'�M&u'V�MA:wŶMt��[;�DR^��O�y3����>�l�ː5����=9�U+Zr�9���*#ozHs}���V ��õ̫�0���D!�sǉD�x�[fײq�r]?1��:( �����Cʴp�R���N���?�)Eӆa�T'&�A��&�~���9ѷ�K�P���;,�~(���&Y��j��ć��qilD�A��������j��̿/�	�ʚ�)[84NoʗL�
Fx3�'ZC?0Z@Pcg���Gu1�H,��HW$�Ql��5O������4�C���]���Sl�hw����|�I���-
�;A-AP�@Ģ�7��QhoS]��5��FA0���~�辖mN������7A"Ԗi�F��I6�~�띠1|=!�*x�Ѽ�i�3�?K�r9wHj�H�-��%Հ��L�͹<G2a�|�)6��
����Z`�͘�Ôs��:p�9�o$UMu����8'��AtJTs�ؚ�3��ͧ�W#�x�y�T�b��&��{��G��-.�Es�6FiIWs�q��醫�R=J��#+���� ���&�؟��Mvh�%`E�>Ef�'	�[^�N��	�;\?�6M�"�X��$wN��(�C��Q�����c��V�z�����h��՛�/�ۅ��,seA$���E�� k�H��+ �U��fWV�����Pt�Gpf����v�v���1�"��$Ѵ�N���e����d�^q�Y��>o�1���]1N��q ��O�zL��D�����[G����0Dbmr�g��͋SD�*���{[
q@dqSy�(]�iB��� ,�}%������)�Z��u���$�Ru����7��}]��^�%�Wg��.�"	����"�%� 4w��ӯ.zC���C�(�b����|a��}@UK�R��u���T��h��ͣH��-d��=L�?�Q���)�B��ސ&�8C���J�l��3�>,�
b�����sLR!�{v�[Ŵ�V�L'�H]��K �[�}}�5-�yDEf�MV�ֺ�	�P�ET��:&�j����X��¿"Sg�(C��}��@�7�_{�Z��VV���/�����r*���K֫n���!�Z���	���]{�5���h���.�aOfV�BW��q�<�(L��W�p]���DAu"WE�ĵޫDߢ�dOBɗ�^/����.�zb G��q�*n&YIjF����N�}�).Qnja�%��y���>��Y{�"��X���%�C
<w�F����*4ӥ�7uWĪE�0�Mַ	M7s�X�[}\u������jceb>�y�pR�;�	$�6Q��}߳]&�������5������̄�`<����������EJ�
s�_'�Q��T�׽��T�oz�e��A�пN+m�ꤺ7YB`��&ڶ�uљ��/7�_�N�	����H�����H<�'%�J�S�j��u�=�d2,�?��'���h Mj	��$W�qV��#�V��ͥ>��gO�~� �Y�JV�1�9)���ׯh�:�s/G]
�wT9�7�M�y�7!+
�����!g�Ngp��(A��CSMK0�l�����;d�ɹ��A*�A�E䃽�>.a[��xQ�u��`��M�x����b�lWrE�4�V�ROʳru���tN�Q�����Y ��\e�<�o���쌱C;I� ����r�vƈ�}�R�N�7���C�=�+)8��^��Y��G�W�������z�<��TEA����J� i��i
b"׿x3O4h5�ʨ2P��ʏg��~�~��W�딬�q|b���KX�b�u�:ZğZh�1�|k���A��U�9�!���0���GVi�{��?ݾ����֍2�ۯ���R��k����P����?��D���h��䪟����P����>�GG&Ӻ}�%�����ȅ�٫����4���ڭ��d�bM ���4�c������i�c`�49�w@qhқ�6������aBmi���i�
U�_�ӥ�T�g�`#�E�g�mߐ1�Ф ��E߱Ph�b��y�.*(�Ը�+�U�L��(�@�x��fv�Y�4��{¦�g��#��G%C����uȚ���]�<o���!���'���'��tE��8�gMez�L��h��Kk�)�MK�6.x�rwx_�P(J�f��2�����Q/ю�~ڃ�\Ɉ��RzH�m���M�g'�O�)k�
ό ��8-�T4{��{���Ȍ
Q|�-��5��X)%�mڨ�<��-����X�z�4N����^�9�e����fK@�"�֭��S�a�~)TpęS�����Jb-�>�fnm]�[JM�!�]S#�س���S'<��Bm?�<+u��/���φG%��^�L�B�@;�rܩ���������g�
�@ѤjL�n\�"�wh����'��y�s��Y��o���ɪ�m���B(S�G-J,/�q)������@��.�%H�0J�������S��T�(����bJ�!��Gu.g]��=9N�9�-���G��ӡ��"��¯���|��c�n��t䭩�h�ǡ�8�Ͱ�q�ĞC7E�Ŗ�t�&��O�
�e*�CS0 �O�������q����8��`U�N4���C�>����A>+�Y�f5a��R9�6��1x{L$u�|<��ca�@�CiU�����{��]�ޕ��{�Q�_A7��j�{}�(�5y�pe�Փ���+��`�eFa��I0����2�-��^���#	O�EU@X5Q�����+��sW�!<��b��+֙��3�\Toи���&q1?��ƃ��Bƅr��}hQE+Iıv�z��Z�H��A}�oGg3-\x��4�3n�A�sPA@�T�@Ծ$$eї;�A
Y�@tkC6��h�Ї�S��x3�1O���TE9$1i
�&og C~�eϞ�����l�*T�N��7�;;���S0�F" )s�����JT@.��и��|{=�2a׼��A�W��Ə����ں.Rk=�=����^�(Վ%�n	���k��H9�l͎3V�x�!��-��ʢ!Y<���yO��	j��f�$S�Na:��mf5�p�z?�w�8ѝ����Ӓ��%��U��ƋTt݀!� ��>�B�\�*< ��:��a��Eb��cBU�_����g���;ฮr�ҁ#P�'�#�4a�Ywɣ�8�@��;�x5a�fD߱��G���)ԧ��Ѻ�{���G*C���������S�5Aŭ����,���k����l|DR P.d!c�GN\���t~�)�do^,žx��ۑͧ"�_�Β��ң�n�b�H��h>=ܞ ��:N$��h����cS;#8J0�K�j�����{)I�Y+�f�0/�Ь�-V4
8/���+�f�2����w#�(D;�|�U«w�P�[Y� �kt��� �y�8�41�/�o�tU�;�$*��ùU��ALi�@v[�gcH���y�6�ёtDÈ��$j߱cY�榙�X��R�33�m�%���SD�Š�|a�w���n�V>��pg������F`?�_r��PI���	�G� ��C7��o7�@�?��Sc<z��/.#7
[�:vz��0��t��uU �������aVɸQ�~ �h�DXJ�,Ǆ{XKa�I�5�"F#��'i��F��D[�GޗN� c����Ы��&�\���fK��Nxyb�c���"}e	���~�`�E"��� ��^��>9�d�'��DOی�p�Bb���!Q���G�/|���BY�p� �[���`��"��9124"0/�C��Y��?/t��'�P�ɸ�N�����0��!�O���]FeDݨ>�OG�M��4�����y�X���?C�
�ࣿ�813'��4�f�:�6RT����UHA	�/,��`�j�n;����y)_0�*�y�t��1-֑�d5k�<k�Ue�=Hެ�欑1_�xK�":"mw[|���4t��bVP�t;�R�|9�H#5��V@4ih�z��Ҽs�sc�P��"�Zv�Ȋj��w噗O��Ɏ�V��vM��D�t͈�
�,��j��Iδ���-R�vJ������W72�h@�f��b��y/��|B��`0�%���@7�`
&�o@1�:ߩ�&��������:��a� A�)�}�f��/4���({�߳�i]�,|@����8��(w�6�_�c�q�D��?M�է��O��&��&,��t���	��<������%jpPR�J�7�p=,�+]t�[���S.O��x7���mP�TOi>GHw���-��
�#�0��!��,�~�Z�Om^�I�(��ݢ����,��\�ܥ@\�~���:���Gѱ2?VEDe ���S������<r��$.��F�/� �ϝ��_<����P��⽰�j$0����`�R�kX��ƈ���hݍ �Ev���l�@fo�@�P"�+��$|+�z��!R����3c�Zr���Y(E[k�H�}�F(��X	�Q��p�:�B�P�c�_V������h6+�b^vm���A��w!τ�x�0�����O��ᖕ���cZN�B��:��{b�����;�~
��Hv�N4���6f���4;GH�sK/e%��=-b!�s3����Ї�l��$��脪�y��ٍ�i\�]6���B-L��G�DI8����#F��|<ge�>��Y/�>�ʈ�����mC�~:J��{*z�4
q�F�(i����窧���`��9�+
Xs2{��3��D6.%�x0�R��n�
A����*��O�Њ�q%����������)jv�~a���
�g-�Ã� I���-N��ΫG�|g���W�/��]�
�%�����������Q\<�:`��b�Q���=o�z�M�IA�(��!H�^�.�U��-C"��)�y������LyH%�	���qr��3��JK)"=:K�#��I�X{hF���z/����;po&���rr����Hz�I��(93��0����"ȶn���b�N�#F*�U4��?u�<�e��|H1�"�x���)۱�0�8ܪ9#���R/1k�v
t��z�6�b�ć9(=S���fD���=��Ȭ��@��e�N��D�6w�_%�bo�X����\�*��r m�8'�����C��t�X���a`���ĳB�<2�[0���,��!�A��PyC@�!�b�,�[�x����$N��]�<ζd>���!������8y)Dr�گr��,	�c)�| /�,� 7��~�ې]f֌����j������Y��>$̰�L��K(��&�Z�H�^�������q�^��V����P��~�R����:%���wn��?k%��xU2Z$����f����4�(%���E��ѧ��pRF�ɦY��57	�ɑK)4�e3����H4����-�)���&��!�	�߆�1ճ$G�5��C�����;¦2λ�oV����Vc�>��E4�Q��n�5��<�	�����ZN�J�P?d����ko6Mu��(VYC��5��V{(��V�.MY`hk<��GV�ku��TPpJK��p#����"P�Բ7�5�}��\�L.ݶ;Գ|�]f�6�Ye��C����@��b�O��^�M$;��
���c!k"R��<�ߔ�;�U6�N:���8�,��N���F�&���J�ek��q�����̃�.��4�͍HEМ�:@�gC����kMGX�`��uu��\��8���P~i$Lz[V2��k[Z�7�ؓ�t(PQ�).�Ru��	�Ŏz�����n�r=o,�U�W�-�K�͢�|�3Wi0k�/��"� ���ӹ9s��l�,�3�~^ȥ��w� 'T}��I]9�o�o37%P�;�墑$~�I)��`�P�a5ET꼫֋�.�F������>cD�_�����l�Ą/q�6�<�������0��e�0BE���M7Bs՗�;}�DΠ���~lFg��G�-xŌ�'�]$o���b�s/7ɗ0��x'�>f��K�����E���햬�5_�7�b:��e����ԃ}�ʤ�V�MN}���D����Bvb��`?+��'�h]q8� '��U�˙���J�ԩ,G�7������n)�ӄct=)N����B��]��P��q_,��;j���t(�qsj�j�r@ԅ�����Y�E�ظ<�;��cT�O;cO&�v鞏~бU��[Ag8X
F�4����J2� _� �w!��H�A���J���ܙ������+q�l�v��ʚ~�}��η��Gv�CL�C!�;�Y/|�t>SX6Q?��$�.[��*�2�G�tq4"�;�2P��`��ң��[|��A�^��$��Gcx13�`��.���g�ϭL���W���)��޸��B�!�м=VY���앐�eh���㽆��B�����:�'?�����x�yh�)en�Ŕ�Ѻ�i�� i� �c��o�)6�Q�VJ��:��9Mk�I�$�@�:��K�-Pa2��]���fk��o7:'�.)���m��L[����r�+0,gr�gĶ��?�*>������y��{b���D���:��o�x�_B���eP}����]b�,�@��D�,Q�AU��:�x��e	�L�ݓù5B/#J{ ��n���Wc��z*:����Ύ�?*f�ޓ�������n,ߥ��Ԑ�'v�_�h�����
���sTuJI��&FzN ���-W�&�d=Dze[��J�y��$�v�=
�2N�)u��GLůkk�_0x5�?��Yy�;)�<�`�?�p��i��Ht�xJ��UؿIΛŊ��֩��"���C���F��MY��T�%�UO��[&*<��?�{'ik㯊��Z�GI*)V1~�8v�@��-��pj����P�����-WB���i�mD�Y����E�S�j$�8�1.	h�Q�a�����[���M�e�Ю%�3�� f��%h��P!_81/є��_(�;��8��e�Ri@\�1�F�g?g�?����H���ک�t*��Z��l8~���k�i۶��F�`�0�*!�v�1�+#�ĝ��c�����Tk������ego�=h<Q��c��L)�X�WM-T?���5ve¹�k���>��1�Z�b'�q�!p�mk�vg������>mۑ�HK���`B�4�w���8_���J��^aҊ"�����ALǗ=m|�ur��.6�S �s4d�v�m:(٬'8�z� ��E!�
2Ey�L�߄[�� �nۮ�a	���,69�yUc���B��7]JF��j;�UWh;Y�Rt�)���jZ#:����������z����'�ײ��Ik�7�!�`�H	��i;Ls�P��Ǥ���*M|x?q����-\�|΀&�D����ZXV�r�ފ��E�a�@�����ӻ�����ʇ�:��� 萜X!I-0�8k����\>�D�� T���ЂC��{�,�V�B;�\9Vñb���� ���F�we&���Cq�D|K�!^nȇ��S0�]�D�ɠ%.��g�pC�����v�ϽSU��x���x��C+�imY��}.�w
(�D*$�X��Ս�NLu�U�+c%��sT(A:/���E����}���m檌�����RI���b�U����͑2��v����:dfan�wW$υ<�p�{�J `I΃;Z��k�*��krIӰz��N����o��}��\�ד��6�j�:N$�y�A�{�w�Q�9�;����6-�7k����.��(�u�Tb��	�O���M|8]q=��2�))��)�}�9�M�	���̣Ks&+�"H8x�}�Q�r|{� ެ�D9TC/.���EIK��<�!�������&��.�s�����^Lq�g��X������T��5������L����F��'�("��@�P��>�ߓ��L�\��'�{�^TqwC�Y�h�P 	K��0��d~Z�Ay��k�*c��4��ʲh�hgݺ���?,�]�I3?R�'��i��3����c7�����,���ƨXh���X,,��6lw��z�?�U���{g��l�M����f=�;�:��jK������+\)���&�rb�J�����@��|�^H 6p`��4�����µS_6v{����Ǣ.�l�gR_�a�6`�����tY�E�ذ�QgF}��ˍ؉���+��<_	��*�)RN�=x�Ǵ�l�_�����B�^�S^M��3�|,�H���ζ7P���3]��b�+$8�0��^���7ZH��͘�Z�4ft���kN�m�J̈��l�G�BWO��0i��r�(�Q`p��Q�
93{��9�B���O�'��z4�N;�.�����u�G�pʁ��{����L�*2�_C�Ϊ��$��!�U6Xz�{A����s�ʛ�&z����Z���㮚�N����T�p#���w�
��F�r<;OL�>Сb<�C"�	pNMH^-9�:�S�x���ħOIE�a�t�3��r0�$D��y�{ ��>�LKAw����m��s�j�����������K�+�A�	�iݢ�n�>�w���o��ku�p]�#^�]{y%-�_<� �_�q��Tމ�T�Q���nN�2�B�Ӄ}(��D1����?P,� ��:/�	�#)J&H��z�*cR��P9TH�P��a�X�0�a����Z�;2~�SPJ�-���N�7f9̷�����P3�uBN��@?vB���h�u�����:{1;/X�����#&�W���A����T �p�~��@��aH�cW󴯻�J-��b�ȗ[ �Qރ8q̤����	[�_�>	�}�N�T�cTm���~��!U7��t�K��<I�_�=�3M��_�|K�&�Z�+4��F�wF��	��U��cj�e��\��}�d���sƕ�S������*�G����f���Z6���:r�?�y�\�-5� ����-����|� �^wJ��
3B���3~�������f�̶ՓI��8�m'�ⴎ>���Qn̶��saY=�Gֵ�=^���<�'H���;��@@���\�9�mQ�E��,n�)`67�&��X���������ZJfC��f�_���ʫ���݉ؖ�k�֋/{���w��a��c�Sѡ��$��u�ѫ�cGM.<�\�G[�c�l۽�U*$��!��G5�z��`u��l.Bh[5ir�L�Z�`��F<#�M{��a����w����Z�f]Da�2�y�>#���C>.��t�|���z�����4C�Ȼ}�9�j�����]܎s�OS��3�������L_��\�%�*΢tQ�i�n**���p��x6��ي�v�B\���6n�����B�)\;�D�p���z3ǫA�& ��]��U3��}��dl��!�UP���Ԋ=�v��HqsUUC���D�� �_4����D�;�Oo�,AX	�U	��L�H��E?�6��P/�8>��ƌ\N�m��O�6�ql���Ap�zCz�,+�"'`:R'O�� �����2�ٗ� {�J��������ѕ3Z-~����S_���c2�H��3;��@���`�@GZ�D����������3w>!�9Ɨ�/~��jRA]�	v���,3�zP82Lu��#;k�l��'k}{~��%Z,D�h�5V�q3�O���iԕu��#a�?�Δ�.�{�[���<�7���[>�k�ǿ��e�z�J6�$��r��8܊����IHȐ#5w��ֱ5���g=�%$<��x8~����#XR�x���F1�Ż���d�z�5v�c@D1��69�B/�k��jx���������i%��p�Ǥd��Tp�������%h|���<�m���	`ъro�5�	�����뚽�QJ΁�$q���=q=&b$c埛�2�I$@��K��y�_�ۡ�<�t��+&���O���=u�f�/\�5�=��W������I��O�'+�d��j�}j�G:��\��G�Փ��Z�R����iiD��������^�}NP\����6#�@l�T��?f��$7���tt�n��Xd��j�؏���"猋�[�B,e�#ψf֦��E��]������q��-h���v3�>�����n�<�ڸ:Rb�G��X[������sQ+W,�2S��H7����?�Y�i���B�=�5���݃��'p�����L��x�1s�\ZQL;	`I�}�-W�O;9pi&$������$��ā�3�H��3�����XՀp��:������%��}�5�%���t)A/�3������q��We���cd�0�%�#L�C0��b�I�~T������A����GG�De������*#݆,U'�L�< �Q�D�3��)�����
�.z���D����4��ܣ�h�/hؿexb3�h3���r���4�8��S-�{�_��D켷3�/M��p�]BK�v��Ɛ��-Yj��^]N�T���4���>���}J���R�;�2���TOۋ`6�o
gjH�:�xJ��s�cّ��=�X:���"�D���E�B0y���~��tq:����L�L��tܞ65����W���`X�"C�K�K�ZҠz����5Z�0���x�j���7��� ���۾V�Lw2j����ў��	�1�.��e�@,6�}ʓ��2<92��nU�aa���_7��ߺ��p`5 �t�r�G��i���"L�U�ը�\����	��� ����P�.�JbI���k�	�Gj����ޔ7�h�i�,Y�ؖL�{Q+wt!H��z�\�ɼ��8�Iix5�j2��N�?[�����%���̊|v�c���w��^�|Th��uy�e}s.
�A�8���/��CZo��
��9�Wtc�B^���gN�R���H%AC]�.p�VD��>"�{������M�{�qq�N�B�H�'x����f=@"���C�Ñ{�T�XA��Y��,J!���M8x���!
�{�)���R����Ta��y0b�i����2����q@n�2�y��ւ�C<��A���*�d�l}�`b6������W䍠�rH��#�a��:�>=)��ʾ��Պۈ�}��S#�j�}�6�)�C�A�3�G��Sص��G�
�U�_x�� 8L|�M�과�'�zÍ����R��e�>�s�˖�^.�|6+ge9�z�dA�3~�	�&��j�]A�h(�������������(ֆ��3�u>&�9w��F%�0��D��V�\���|E�!{�_DJ�k���63MY��4S�s�)��Y����\H"�1݄xJF�����~9���� �%`�g���� �HG��H$��1[R��
�`���X��Yq��NLb������f��+�]u"*���nP/�'��k�je�vurgc�Jox)>�fq� ��L����i�L�鍗E�	��	���K�4�dz�V�U�|s��X4�J��o�[�T]RoY	G�ŅtG�����]�u���55/��1M�����%�M�g�H�4��p�9����t<R�)j�Z�?y:�o���V3Ę"���=�O���L<-���y��g��U?���pzTI�Mj<)�N�wX�36b��Q����JP[S��^t����~��:���<Jbm���aV~}��K4hA��g��qX��?$UW��ِ~0��N�҂a.T~��L;H�T���1��f%��_Ā�Mz�I`�u�ߛ�M䶵{�4	����"V9����=����F.�	�\����7U_�Y�}�`vY��S,#�T���wY��� �>�8t
��Fr=/�R���!N&���1��b�4�ʢ�K�/E	�Z����v.� Q_��4@�}�����"��I�ꥥlb�ނ�dq��R�˙=�6�]-w�CP��-;����ìvk�n4��L9�[�\�9�L]�d6<�^7�|�5$�����
�ǯm[��<�� � �*3��7!{�e�.��PgL�����qlŠ"��e�8����O�dZ9)	9T~����(��l�L+dǣ�v���2+���dP�
%^����1�^IZ���#>�}�����ƺ��ߜ!
�+�����t�\�UPOa��̶.�����Z�|�=0s��,�s%�0��3��^��3=�+`:#�����
4���5��Éw|�	 m��
�-���Ù`��P������%\#�XP�{��qe���|�. �{�6�I&*���X̱�gL4�5l�cj���K�v����%}:L�mi�Hڄd7y>&�ڜs%Q&�Zpq��^���r&B��sn�O��5b`�]pfՔ��M�Փ�c�َ�#xEp��$e�[D�ݻ�8�l@t �9�)�
��z�8&�\�WM�"�@͓4/�<����v�S�BSe�J[��+!�~�Qu�4�^�#�䝭z��>�5Қ� �`��3h4��	��%���[�����:�^r~}��Je���g��gd?��eWXX�M�uwĦڋ�[K4X)��$�F�s;y�]�Igb��L�r�'`k	�g�j[��̛���X��E���o�a������狷��R�֕،��N�Ջ������u�D�.�A�� �'�c��o�E�_�tN	H��R0L;K5N�^ߤ)(���[m�+��̩W���'�&�N��Bsal���C^�Ѡ�R��n~�����[V@^@A4U�BEM��	���A���	x���.�)"s����������f3V�;�xC4f��������<��zq;9 ���{Id��~���m�AJF����z�@*�*��̖P{��)��>\�{��/OӓE&�Ք����i���6:��e15U�(g7�DS�N�	�'���j'�HH�����k��Z��wQ3�x��_׌�3� �G˃�
��F�)��$"�E��5��6��ʉσ~������
X��S�yS��J������
�])���aa]��LAi��dU�Xąݚ���2+�Ѐ�"�$�c̫|B5 l��ʦ�pK1�EKz�w���┫v�9|�hm'��3�����6=@\���mu�����5�T+�����莰����K���6t��W	�칎�M����q�N�QȈ�r�GȤ�Ct�{��M8�z%�{~;uW�#t����D�Y�N��[��z^ӷ�h��p-����=͕��Z>���1b�;�X��?3۳
^-�P��s�X|mq�t�
�|6�-u�D�sWbm�����pU�e��!��+�X���7$~��ص)��,�R�L�v�(���x�t7Èf�����ADPRwY�d�H%��_��;�2�O�8B���ijۘ/�l�
L�>�]Ѣ8
�t���Z��{g���(0uN�ɷ�W���;�X_(�W���n8d�I����K�0��}��kM��DG�<� *��՝�ս�6�b������i�[{(DyDxsД q�*��wC��1�q%b�%�+\F?��	�4>u&�j�CL��)����:l��}��ya��Z�!�I�_����+AwK�a������_,���G��3'AsD})N;��E�(�[�ȋ�����J�?2Wbrࡐ�`��Z�W�^俬��f�l~6���벹6��l�򯅦*	IM'��_}T�/[�sk󾫧�ό�%���O_�JW=���u�*y���P�݋?�Q�9]f��?(���6��A��BO�B�����
��z�@ޣ��0�i$���|�i���ͱrful�^�n�-ɲ���xQk��RDW���o2!��f�=�`L�,��9�Z�ŝ�L�%��{=�Yx��wy�h��PW\)���6���6.��ʒ@�����)�4����b
gx1]3���6J~4�w�г��d��h��Э�������*+�?G�&G�Rb�"7�:)�+��^����֋���A�,;��o:)3���zP��c&m�4|��G�)Eκȕ��P+g�T�E��Q�K�f֙�dqz%�w�%Ǭ�` �̺��/��}�a��L�8"�O�C�^x�����g���cZ�övBHNT�����b��ԁ�����N�yW�Qs��,L����\�����E26=q�Ѣ�^+���O~e�+6�s���R��%U+�f�ۯ�+a_���NB(�a�r�<�S7c�:��x�����#Xԉ.�TL�bM8@���|�%���뇄
$�D
�l�^��!��1V��)G�Ua�Y�)�^��V�R WO��[/	MN�gT|:��_��	N���I�
h�򅀐w��i��V:�G	Q�:�'iBK�͟�(Z���I't��R���t�G��yH��B�����c� �a6k?ƀ3!����y1;��`��ͯ�� ����`J ��G�^��ҟ�����#��XH[{o�T����m(�$Ϛ�<�D�F�ky�  ����� x����s�?�o4	�N\�IPO�U�����6�������o9DR�ؗ]���+~n<�/����ILY@F�˺�;��p��|���`y��=�T�;Ɂ�:�g��cPf��A77�AP��5`���@(�=�d��-��Y��T95wco�J� \~*�B��N���SH�y*b &c�EC��T�L�'�(X�@�кF�c����2{a��s*�����u����]�W�i������<� ������2��#�5�4�����ܭ�7<VJ��ìǤ?_>��N�p�o��*^��I��g���}�� 4�ƌ����
Y��Ty���HV����K���W,��$4Of��d�})�i���AK�*\}̇2�@���b`.�0o��"H���:��Ty:4A,�A"wa���o�\�݆����QZV.H(�(�O�MLYh� F�W1QՅԆ!?�&M+TA�_��O t�
=_L��
P8L�=���o���֮v3z:
�R��X; ��є�q�s�3�1'��AF��������kUm�"��_ �<��"�4�uqF�&�h��_Z�N�pYK����I�0�3٥�qq�H�,��CP�j�;�H���y2�xu"\[�I�����1�#�x�&?���O�7�{ܧZ�ⴭ���Fp����:�H�^�@���^ 'ĳ,(�)bDQ����A�fԽ��p���O�>��>B3!�\�~N���>qu�p�1�5{m�忄%U'�.��?` >Z�c��b�� �·�G�,�L��=[`���
�Ax���5b��@��4~|K&�1]���g���E�7zx�U4�Lo����-݅K�.�u�WC�$Z!6G�G�Yb8��q����9���@� LxI��z�ԦM��Ny�~RpN���sz$��Y�������.,#�l��}���i+�WN+�
�Eg�.H�r���z�︍�.@���28%��F�O�
:��W"?�$Fw�`��;����a1����u��Ȅ+��[�r����c����YP�����=���kҳO����@M��@�ɫ�"9
a��ܜ.e�N�U%�S���*��DH��l?��ֹ��7Fd<���o	O'�ߤY��I,@W�#�Dr�cc�e.e����w�v]�@U����ϰ'x�q.�G���һ�����C����}�[H�Q����B��3`��In�x��S��80��'|�a^��g�n�#�M{̄T��L(d�,��	��$r��3j�7a�˃���Du]�]�0���+�洞��C��r]�i�V2��iS)w��[�Y���Hj���w��OPC�hȉ,����u�VgՑ��%�wO#-���Xx/�F]S�+�I���~�
�� ��p��qi�QL�j��k�L�uqͣR˧<�Z���8�s�!����q�BԶc��]�xE2�Gs�;E��s�"��W!��Mϧ�C>�Ǽ-)��p+&w�%n����!�o07t$�感�&�%��}HH%�I�{���'9~^�1�Q]H^]���l���QJJ\,�J5�I�� 0��FMm���͉�\'e鮷�^c��7���N���=? ����8�~=X< #q0H�\���$��e���r����B�DI{��"�{:C���*)����N�����"a�ūK.#�:�+�QwM<A�{��2��j��w�(�Q���7/��m�)4C]��x�k{��rp |D��=�E�O*Ί�95L�$	a�Z��$�^�n t�FD־LO�7yR(���Tx	d�:���w��ȏ_�n���Đ���ΰ����LóDВ[o�[��BѰG-�2�]1*j���|�������Ȇ*�����W<t�M6�����EJ�zZ�I��lm�ޤ����?�d|?�I�-�]�m0�}�/�JU���e�r�HP��W�j滴C�v�n��zⳊeG���2,xb����5`nI����>EHM	Ѭq�K�b.��mK�g��!�E�X@Qp�©����<���Mڹ�c���c�a�b&j��8� �����KG�J	�;���)�~��F�R--q��1�!.����/>��^"FΘpA��&N�<̌p0L
�#�l�6�˖]��0i
P|ޠ.bꪴ��x%XXς�kV���{�Xj<q��N�`�qBk�@��������<���'��9� S?��KǺ�fR3�����ғ%�݋��:E&��N�6��#s���#�4�ǆYb�O��E����A���cXE%��J��;W%���p�.і�O@�)��B$z[���,��7�9���=�5k��
�gŊ�|�Ɣ(	b�}5Q�]���;���4�0N!�lׂ���,p�Xh�,�aݼ@�^�Y���τ#�)]]��\ �ᘽ�{X�1F5��
0�	Y�l�s���KܷK����Ң�ࣴ�9nj��4n�� �r�a�҈���rjV���Ӫ�`�T$��f�~G�}�&������ls� ʒ�tɑ*�|����h#٬c[�����Ϧ��)�$��k�����;p������A�����:[�ݕ9Td_���f