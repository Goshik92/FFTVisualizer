��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
|)t�]з;�Y7�^���y��Z��(&�ς��%2�����1X���N��x}_�Rd�`/�-����"�'�S't�+"mRUp�J����9M��}n�a���`����*F�	���w�4�bu�lw�6.0p9Cb��q�\�T?�/���෰�=�0�lcy{{/M�	:[D���ua��yyѼL�B\�n%�o��Fj���_eOfXY��7dB�r0��o1�2� �1#�g�,�w��|6�x���~���) }���*�0}E�C������z�/�P�#t��[�In�+A���g1�뚍u��dԹAT���W:4��ټ�e�Yӥq�h�+��<V��<aQ\������:\ㅎ���.~�<*����.���Fs��2�i���6z���KQ%��B��&c�!�D����:M�O!�"х�G�ظ,x���	�F̈́�tV�vS���]�������65Z����˟Y ��&(���rLo����X��FK�M���n���+�(�����#������{ρy
���Q���+Qr1V`����{�\~�^�d�c�b���9r�°"���b��*i����% ����0l�h��.l+�S��AjkF��O�m'c��.6@z�"�L���G����d�`u�e	n[�`J����.�z��"k�6cG��+^;~�n܄�r?�gT�F�Z�H����i�����1Ð9uY���{���Z��?���t����ѥ��p�&��u)��C��J�]�z��ۈQ���|V�@K�b��h�HR���hW�K�:��A����%��kC��=�~����\B���Z�{�j��vJ��W�1�e�I�I�����4���c�����O{�T���e�@�e�^��Ї
�/R�w�`���JV��i��	�]�ۥ�W'�@���!k�Y�o�s�v!���f���Z���`G�5��H��vD0kDkʛ�D=F��\�B��d�q��6��������U�{�����:�Β�8��؀Q��ttr�P;�辰eW8�����������bS�Ѣ��*�����"����6��
�y,���n���9��n�}��O���醰gT��v�!b�n��v�k�S�B����Yt�]X\��A��P��� ɷ�H�/TU~��
Qi*m&�g1N��:�&RR��=�U��������d�ܣ��z���y���t��J��y�[}#A|L��"6�R��R�1��uC_
�V3i^u�=Q��Hs��t�$�B"Y��Bݩ5�����Xb
���Ơ��K�zB�l[$Nvi�!G�	�h!h��B�皙�L�ν��^�؎"�����M$["�סD�	�E�LF�j�7�jx�}Ŀ�m�KE�%�J
�	ů�yVL2	dn�-$�����9d�5խ�|)��2���aN���_Ni����k��E9I�&"t�I ��~��f��=qk�;�_tƀ�sr�	���B����u�|�E��h�}a[�y�;����|�ͱ��W|�9�fj.8�d�������ko�
�Z$]�%���Z�O }��ަ �˅|�%��L��"�O�ѯlE�"
c-���.��kB?)�_�\�����ؐ@��{[��v� d�( �"�/t��v�-�t,7��<DAŇ+b1l	���q.��#��V� ��w�U?����X��X0�',}O+c��*��5�[@���N j�h(�a&�5[
)�8%f�D�J�P%�O�����U�GA�&O��'2����$�D�ciO���ļk�~o;[��t�&Vؒ8���vxȨu�|��mf�R���Cx|�@t��̹��O�n	.-e�[d�L���Q����������?ɜ�/Me�T��*��3+�9:�"�t�/��a�-�\VZw�#�0��;��(�|��$�y�³Ue| J��'nhJ�#"�fȸ�&�(�_�1����IP��_F��7�\���8x�ׅK��̽�Q��]FP����j6~"��@����Au�|r~��ϱD�)���E��|a��={��:g�-�z��̷���i��w�S%+��¡j�l1�%��U��¸[��;���Ц�(����12���n���:�/�07�&�g�0mSГ��选���*��eĆ��Lbx1�������f=�e}��Sp7k�1�0��֣G���`:ܧc��i���Wl�>sBq
�솉�-�A�Z
w}���]`�3?,I?8h�ut����2����Mz�U����ƾ0����Z4>�8�]��B� ���f���n,�^��3�0r)���)��()<O+�g˥�b��0E����vێ�C1�2:�U��f�YX=0<���a|HLPl'����S�4�E�����`8Ʀ�0(-�䯔�Q�#��&7q7uƟ���K�[3�Q�$�<�	��a;K�4���vr�cZ?9/�����E%��{7���b<������'o�	)�p&%�|���-��
���i���޺����.�<&k�������"]�ۤ5�R�Nn}����ʅ��R��:?WZ�N�eu瀄�j,��]�4M�M�9��Ra�y�ܔ��������D��������68b�ϑ�����.��_l!rj���_��dx�K+��3� ��W����(\v����ol<�Nڊ��.B��:�O�q�J3�7�����(����D��m��Ӯ�ܚ���z*�quDdnNd[�����w�Z$���ͽ[a�;ϼT���t~1�-q������H���B�ʟit5z�יD��:�ԫ�s<|��(u9̕�)]�e*��=`sZ�vb)�`���ѷ���OWwP����Ҹ�ה�^�"ց��k���[�*{pn��O�����E��8|"h��F���6�e�\lm���C��q���KF�7��	�H0���>3��86�'̦�Ҙ1<�Z�����=咥�J.����"�|iaY�t��T�������k���v)����� P��naK_�|��⋯�E��`�"�	~r/���>0J7�!B�vZe�}�4�����m,E��Y|�!��%���a���lf$���X%� ��l{*���n\Ş%�"�֊5L;yz�L6�q��!��y������2�\nu�lGb��f��J�BX������5�2a �$EI5Iu�7AK36��.0	��?���(�F�d`?��_�2=o��@���m�}񤻲�O	�$}��^��>�s%�>@é�V���Z�X�i�)A)]���t���?(#��j��ڶ���QBA<���\)��dZF��\n���� ab'Z ��@�(	1�hzB�>���|V)��v��=c�0�ړsڏE�:QEq)�N��]6:<�j�|�}͈=��,){��,�z��=����#��^(�Gڪ�6@���������������C���;N���X��O���?�(Z	p72�o7�Ĕ�2�x#Cg@��ݼ�:+���B���~6��
M�$1������lPw\w����U���'L^	�� KJm�q^H�~�l'3BT�EA�"�B�D�y���U��P�{���k~:@9�K�D�A���L��l���_d���{�:��O�p[��,�~.���g�e�E�[��@����w��]'������]l�	Ņ�ɘ���e�!W����F��$hɯ��̍�m�7Z�6�gz����w�PN�,u���: sGv4�R��P5Dy�H��>=�*i��o���Ż���G�dg)e?)p�ʆ�7v\2s�I@EF�땚��|��U4ԁ��(�*�I~K ���E������P+�L�+���`��Y�G���R-�����Eo��g&H8
3+�pK �zL~��y�:-0\�W���ٳ �n��j�!N5��c�&�o��CV�A�s�^�@�o�m�Z�o�5�����ʠ��ү��d�rmb��MެyZb��Q=EU-�9I� �P#���	��yBaswnC��@��}��3]6G��}����U�W_�2S�ɲW��������X�GLiie-��CJ��]ƨ�=S��Ӟ�R�o��8��Vg�ooR�!���!ؤ�gV��P���Զ��QԼ�mm ~���	���(���#�L9��a	��Y}5kz�����MID���\�Heg���;��e5�+��;��4����h�8G��~�5��"#`a� A�o����Ub^�wp":9z
�s���R����v�����]����>�ۼB���|u�����(����t ��b�D�r咞S�%��׶�y�$;b/-���0l"b��S�K����A6qE/�.���� �{��{�-�m���q�������u����>�I¥m8�;
<����3���T�E� 	w��ڻ�U�����.�"j=�]��j�/J�u�hg��f�j��a>>&��.�����~|�K�dN� �b�쥁��=��UR-(�w�{�!��H-��ֵ�V�o��W�<A�4�-)��?$b���{zO+\\*(C��TS`DR�S4rN��o� /�W)gʽ;��%��5��(xd`j��9J���V��+����,�ّ�����H|����9��G���ߺ���\��w׀��(�k �O��>�'^���g�6�0���Ҁ����
B��G9�~T���h�B��j���f�Xc�~���
�+IՂ�O.b�Z+��6�l�{>���;P)g���Pf%?G�^��h�]�����JF4��Êa��Tg�A��S	��vxݡ弰��>"�[��K�)IzU]�:H�|�{�X�~��E0CA�u���Jq�=��:���B��{�Q�95������?�w�9�͞7?��~!w�������uR#I����k�o�ΔX����N;���s�n!J�H����6ߒw)){��RX��Ɖ��1f�㝯���Ƿ-ym��Z�`+�_� S��wQH1����@���Xk���mH��p �哅v53fv����R�ט^��*d�'*-k��|������5��z'2#z�($��yC��A�Z��nuo�k`@ M��1Y~D�y����D�{��4Hq�Ϛ��0�����{�n�v�X�J��f�0�Y:���!sr`m{�4H�#�O��`R,��1?<\��:���]WH�d�I v�Ar����q�G�{�����Z�ŋ�]�E�q�.� ��3~E���_M�)�)�>]]���.]� 3уG^����,N*j�c���X�J���8����*"(�+��,�M�L�����wD4�9����8��]$�
nh�ΌtލZ�~zo����K˪����c��	�R��[���6#�%��`I��,���#� �m�Z���L��A�Ͷ�9��y�0.���(Ղ�CCכ�������AØ(m6�%ú�58� �q�4|h���$)&}�NT�P\_�Y����z�t�:6��%fʍɂ}��zIɌ��HHh�Z��m.d��*�Q|��c��e�v�g�r�_I�0�<�ȸ�{`-Y��
S��o>�1ۼ�d�<w+���\����Ɠ��XhVE-T���(g2�'��V�v`sM�.�	�Ꮠ�!��U�n�0��htf����$�W�9�v�R8�n���g��- q5��(�����d9�9\?�SH��@��>�vx>Ǻ�s� I�bv%FL��(֛�#��]��s�@�+����XQ���_k��c{� LM'�k��+>A���g��4��H�!|�z`�B�1�E�$<5���D���e�r��V����\vФ��{&p]w�$>�GϪW�ǈb<�j�Y�)�~�`��T�|�" �xQ�"����@&���f~�qD>eo咽��`є�v5u��> ��ݓ02��2lN��t6�ce� �7m[�J�r���`OA�޲���⵩A`u�ςVj�~GUx�0��9Ƿٱ_6A�ՈQ`Z��ۧ����{���� ���di~b_�dp��M)���ȈetDӹ2m��9�yQSz0�!��gڂ/��dG���N��o���PR��g�W���J�t�H�l�^9*�˚CwJ�>�؂	�_yY^��n��9�z�ot�tno��YF��p �;��M��!Nߗ*�5+�2�~�sL�
kFJ���m��W1�I�:,��N��s
�ǖ��+���0�/C[�`�:g�6ő=Й_-E"��c�bb����P�'$5OE?��S������јx����d]�QՌ��6yͰ1�,��+�ҋ{�va�\�~�������Èx�3{З���Ms��%+w 5h��:�ܔM�X����ZJ
��|9�vR�[�K�ČI@��(>h`u��N����k�.��B߄ttg"Q>�{�E�~o�zř�ꅰ�f9��D�o��ࢀ���q���A��.�G�'�TPG;�Z&�7Z��GgT�E��� �ڌ�L�ˍ'��h~?~�����\�nĂ�LyL�x�f��qp��*��` ��.z��;�/v��|����E��^�:�+k��k�d�J�M�𳮳�A:�M�m�i�`X�e�ӿ%� )Yv���r���
d�dRgsCxԅ8����:����q�{�-���������-&N}}�X���=�ó�n`�X��T�C&��Ԃ�����2Ǵ`����� �u@!���y%Χ�c)w����i_��\�^��
y��y�LI���mq��8(�m�FS� *_���7O@ 濹�H
�k����&�z՗+6���OB�eش��'��/Uw�_¡2�Be���f��Y}��x��:y\E�yJ��Y���_x�c�E�#Ŷei�1��,��"
x,��Q<���gl����(R^�N�O_%+�����В.
��‱x!zS��i���^�V)�K�F~�E�R�Eь/C^�б�Dt�;�//��w�L�l`�-�Ao'K���E<A��4v�B��]P((Ya��rk8ź�PT�֗�������I%��,
V[4�ʾ��m�V���*�f�/'��[簲(��������P��Ze=�Z��5w�U&�s������=��j��ui5�,�,��}Vs�u�����Y��>�*f�gF̻�����y��Z�C��㯂ι�p����Ek�/ �ٱ����ى���Y-N�!u�xk�lk���bZ�5�]��Hm&CA���=�z<�`ҤJ"���|s�¸���U&[�/�M����198�f6�vC�8͚F�x/��X����t�8w����>d�"�/�=�`���C�i4��ޛ=mY��N�4���)5_$���c��rub��R��rD��?A�b3��TA��~�g���֖lᵤ+3d���}@_��>��%g'zQ��1�w������?��V:����[�x���4w��?��bˑENڒ���i|bu 6QG۬N�F�<� W�=����YS���fd��L	�7�$H�3z?���q*�1q f��K ���7A^s�r
�m�T�K蜸�l��R��rr���r!q"��*WR�aJ�ݤ�8�������2y���}䆘�4oO��ؤT��]f�k�z���ث�cY��bs���:#ǯ���Y�B�W�m?��ѹ0�~[�wڬ�-^k�-~e���NՏ(��`(7�����x��ޛ��u�#�qyϊ��!#�z��ѷV��*n^�է�?��G�+�\��̑&�|������?w�tB]�K���n�-�~�\X
c�-�[m�@w���!��b.|<�"�9:">�q�L'��!�w��J��d��Ԕ$���Q�"���vP�'}/����g���_;cX�j���휅�7ѤD��Fol�@�&�9�9$]u W���S�h�H��{��	Y,k��@��+���O�.�o�8����Ed,�S|U
�z0���0C�K(�i�BB�yl�Va'�W��M7G%Y��L*�5d�L�8A+�{��{(���h?W��+y|]���&�f�)5�	��Y�G�c��΢����X���v�Wy��@gL=��"��C�xW�< {�&��4"p�I�G�÷�~R�m+gȩuD�录p�+������F����y�4�O��t�)}�\��?�WY����|�Tz�}I���؈]x�]��Ɵ/����ޢ��y\I���Q���䯲\|F�����e$�����ʯ��fΪ�$���|�6�:��QdW눀����[#��S���Ŋ?����	E�*��K��#�
�7Jz��,?u�>D�����j��W��'�K�P�:#���Yg�R�`��eV�_.I����٤��h�����%�.fXΤ(r�y��0�F����I�������R�媦���	�H8r��w��u� �d9[��JG��d�0����/����5ī�8�¢��ձ1#�
��)B�x�/�_X��_!;#}K�FX!</�Ut�)���u�Wܭ���b�׭y�׵Fd��^/�j\���ET`+�����s�iJ�r�e�O�4��C{k���л����Rm�:�9�
&'X/���A2`ѴOo�d�3��@���N��c�_�����v���->ģ�]�V]��g�{�69d���Ȕk�=��y����LKR�'{�>����ߑ�|CD�N�,F᝾� �Q�����9U��m@	�P�>�'h��,N�B����m�0��RQ-�Q4r!�=����d?s4�ǲ���?Fq����xe�ŗ%ȶ�@�Át��U��:J���]��.�0\����[0;"9"])���;��x)T�@�֍�d��B��6d �Me���돆>���k�C5��(�����ؑ1(�EmKTl�_�Y�f������3:�����*O{�p�����s�cU���s���1�%_���K@���Zխ3��Z�ZC:h@ߝ�ߛ\ɔ�*N=:����e$щIT+z��[dި��z�5� +y�F�zV��TX�r-�&�0N�}Ւ��3�8#�p�����Eľ�	 _PYݯb66���,�a;�Q�c0�h[�r�����Z�e�h�<Kd�5Z*��e�`����{1������u�)@&��]�sTA�^���L�8�{�d#�d�l0�µ�=�����曚��S��g�0
��U���Y�:��":�M_?��<^
����u�_��2)��a�ȯ��V��*�ˌ�J9�hzN������ޅ:���·��B��-��sh^�%c�C�����ɿ��!��R�g-��.��4+���N�ؐ������\�/VV����7#�Rc-��z♾���Z������Zn��]����Zc�x�d�W5	Pf�,֒p��������z�,k�zD� ML.Fj:%k2�O8�И̞,�Z�5��M�{�縷")�yJ�?�IN�$�A|�՘��}���v��m��.t����Ɯ�N; ap���r=��d$k���,�f��~O��k��mf!?ψ�Z0�#Ed�+�A3���{&3����2�t���� v��Jd�>�n��p ����[�#W�E9�;�6�/X�_��	�X����9Ļ���yغm�~Ƕ�*e�[/׉��Vf�����A8T��z����i�a<QK��@tPb�P�d��5���{��8%ΐ{�o����i�\�|�`0�ܷ��b�z��R��1���г�,�f=2������G��B��8F�5�~0�dN��3�Kq��3����jUJ�����w���.(��i��s�duj�rKR=%�����{�rS��~�--��۲��62Q�}Q��B�Հ�W@.[��3؝Q�D9��X"���;�=HIT�s��v���V��|�|���N�]�������NT�	x��SZ%��3Cb��̗\0Ҷy���le�E���t�'��^��9渚n*fO-����y�w�gD�����ۙ׭]噵U�f�5�"�)&uǦ�N����	񝠀��r�ǐ�F���q������(.�E�bfC�lN�4G��?cLQ1�`�Ad]�t�c��UZ�6������>�X�+��.4pY�ⵧ�Ѭ�ɚ�JDi�d]r�����M��7�bt_˯Are�yP�7�}v�n�-�uL��+���{Z�o� iQ ������
�/���K��/���Ю�k����Ep�X���?(���� �VE�>���~�g��31^����A����)Ȑ��^|����"x��ܧ��@M�nXh���u=d�u���V����&���C���ৱ�ry��![��u��T�}%лfE7�ҭΗ�Ǽ����:���Τ�{�M��#w�����!c���?T�&��L��uU�w��*j����B�!m��Y�F*�����B����,�<p�`��?,�H���zm\_t]B��'�y����Ěb��zm/a�`�=�e;-�}�ˠ#���KL+O�q
�T�/UP7�A����O��i�xA�OO}6����U0�M&ha��q>M��t�k���R�zj��b������UY�R�'��+xmV���k�aG��KD�/aHш$�,�s�X�.����Cė%��KZ>��9�	�X��/;R������~|��WԷ�ߙQ����6>;�v�Ȟ;e��5x5���voyN��B$��4؟�q���\���>�|j(�(���0�ػ-ſ4w<�1�*�Y6�Fsc;)c,�'���� ��\�*C���:2�~��:�M�~<wj�N��CW��N���G��]�0��:�%/�I6�gՠ�T󛧫�b Ș�?o/�2��s#q�,@[A-r��\�1�ݍ���<M���v�nj��!D�L�o�J��S���~���W���iA.�@����?����Q�����@Y��֍�ɪ+�E_6�|DHY���ts�I�I�+���6�k
Ç�k`)��W���5n+[��̜�(�����Um�2�<�ڱ��a�; ����4Ɂ����J\���ӡ�*��F�|;>m�|�X��B�Vv��k&xݳBr�4�1��k������Q�9��=U#S�A׀|��;]���������
]L�PE�ɡ-��O�qGAc��Ņ���<b���vSZ��"��ÝD�r�7T�t� j�K�����t��T[�P��p\��.[݄+��)�Y+�Ux<j���_�T�O�sq���1=��E�Ã����h�p^QR�^��=�W�? �D�I��~�1�7yC%��(�n^��� }0��H]0��X��1V���e�m�w�zٕ�B�g�� ��KZv�+���{�
�̓Y��
���?/Х%ZE /�~x(�2��vf�t ��"�>ۀ��������TI����
�q���v�Ϛ����&@����Ek�"`�]%���Q2ђ��7�����?7gzKug$؍��y0����P3m:A��1�Z�A�ܿ�!lh�R{+%�lyr�u|�w�R�f.滛}��g ިVƤ���}6�kS'�9��ļv�0%a��9ʥ�ߖ6sv���4��S�>�=�0j�$^E��Χ�jQ
o��}i1�z�%�OCՊ1����#Ǿ���I-`
y�|����KL������K�!ƭ3�r����Q�/!���,��j���ڹ�?�})�4(�i6�>�~��}F���2����3����Q�������|�X�X�:I^����e��⍄����!Q
�<�{������>=�x��0���]���Q�zZ"�B�I��dH!�ῦ
\�������/� ��O؎���������}\w�j1���%hy�J%��;]4~{V�Ƚ[����@�I�գ�~;�ޖ7kN�.��|֓��&�,��
@~d�9KG�gu]��,��~CU�h�f�Q2C��ȵ�![qG�$v�E���J�����[>�z8��~� I�xP�M�iOX���>�o-��[HQ,�@�X<&d	�R��E[�Bg0U�#HjL���p��(_R���{}Ɔ����9Ű�dխ�|u�R[���$��s���}keS����g�^t����s��s���������ÜIe����i�.��'��9�dy�=6pE-�Ԝ
p���������+����,�	�I�3A���OVRq�dK(�)�����3����T\Z���.K\#�U=�{����US������+�MW��0?SÃ���R��9�٧Ô~���|}�u4�<o�xPi��g�����,�����\N懴�Ә���)���7�䦹��k����N�2u-|=���+��5-�C����;�3�����Ȏ�j�.|�p��2ӕ��NM$p���EҺo*�`p���(�.\`0~g�/���|ۊqˊ�	�O˕��r'��_j��.�^⛝6ڊ�/Rj�Oݶ�S��a��
\'��ϫX�Lξ���'��F=jiTc�	�U�':Qu�eK���᪇eb^��؁�k����7/�2AUd}P'����i����E��2�.�ӳ�� a�n*Ui]�|3U}X�{D��$� �4���n���tS�rS�C���r�c����5�{2P�TS�Y0�ͧ���.�β�Q9z�R[�N�F����
[u�I9O'M��9��ւ8Lr,$�}�Z}�8�>�_G�Sn����H+\����̩�+����PG	�=)ՙ�\%R��J;��
V��z�%΂���>�ͤ���-Yڄ�+��y�|�������P��Z�%����f_�2��0�������<5�ZYW�7�=�o��Z�Mm :��,�s�яI��D����1�\�o&4-�܍�d����KW�-շ�����;���	ù��Ge?�yOVlW����}Ri�t^�l�֋9!���Ӫt�YT��J)c o�ۻ�IQ4j�����������!�~�5g�!�b.K6�d�4����ʌW����`�c�8���'����~Ru5es�%.�k�[����6���n�F�x���,��`���h�\�V��߯xR:��#����\�[��O���?@I���6��#o��3�}�)�����E��\JP�S}軛07�:�� �㩬�yX�"��b����#�o�g������'N}L���Zk+�������Rb:F�8 _��ҶP�(P��H�)�`qӝ��0WOsğSigz�>( q���>�[�l
#*�%��H��c���̈�ɘH��̀l����g�����^;����gZ��K��E�%ڌaN�E������p~��]C��.y�-�Ջ�4��b�_�OGtOy�V��{Y���i���-���y�%�4���V���DX.�m��Rj����"=�>���%�F�۠�g�4�[���{h[���Ѝ�_�b�-O,��=;9c��l� 1��f�zh}��c�d�H�@��b��@���]K%R���Y�T^��T�ρ� ��̯�)W�3��f��*:�چW��:�ܴ��K�Qw����$��mx���e1E[�5Oҟ+�����fE�xM��E2a~/�ZS���/�:4Z)���;ll�_ګe�����x
��U�����Ť��f��,�ʺ��O�G�*E@v�Ȫ�1�h�����$�\�����k3�8�N0��}�BE_���ǯ��R���ks�*	 �.y~��#��m<�Bd�K��5�[E;��ߍ[;,*��e�Q��0*��kd>��qK샯�h��^0��o 9ͳ���B����O��],�ցu���a*�Q�2AZU_G�;*�\�g����e���(�:��8��
�XS��z"��t �^��W���U�JZ	y"��M���"��m��t�[D���}��լ�|y�)Y�:�3!U�y@�-7���6H�Pb�:M+i�7��}յ���I"�eı�%�.�Zt��@��&.�n�%m�D�	� H��;�h�̝�w��<�`^J�&ԏ��v��?��{ ��#��d�>h��2S($�����'���
���>Sq��݇��p{��;=�����4���y��I�ӥ�P��ϲ%�]�*����34@GX ��%/Mtt�J��@,bŐu.^L8i���7=O�E�ρ�g�������4c�1Ň���D'щ�+_ɚ�Q���<��fA�fy0�����W�Kn�~; M1�Y�	~�����F�~�2��0k�=���	5	���nψ��=,J�|��oA�a�Q�3��->Zw�,��?4ٜG}l����H7�As�����̎�_,%D.��s��6�7kJ��9�!��W5m�2�*c��	��o��H��J*@�*4!��u��o*�����D;腇�Fc+�L�o/�����o#GR�Ŀ;��a���!�
���H����څ� rJF�=ؠ���%��U>=2>����BQ؞��\j��U�b���h�Yh�|��֚��{��������峾�"��?��u����j[$]�KDM}j�� s�}��Y���N݌�������������߉'��ݞ�%RP�Ɂt�t� 1�ǒϔ�4�s��U�0I3�]܏�������(���JC:��W��T���H�45o�>�,�2��f�'��9����	��`��Z�@(Y���x�T�����Q�+��Gt�0��]cD�J�|:(�
pU�;��w��=Q@�\�@�M0E�g��&����B�-�١�:����;��Q��o;}�gUg�U$�[~��i��2RϦf�7�nM*��ӧ)F`=$bp��p�ұ�T�%�n�l�yqF���<�}�L����ࡗ����iۗ�F���ĭ$u��>��8V7aa�b�_V��~�He �L��̓�4;����ó��:O_܌��1"��QK�m�u��ػCp�����4.�}�>����\��Im>9!���B����̂�<�Qjs-�p?}��ax����5��$��T0('��w�4-4��l�1?�	���Q���*���e8�����b
65/������7����O3�������_�(hOP���#�M>��"�S�N��s���xcO]�U{��2���innz�-#��sdV�� �A�r�+��ʕ�K0vJ	���H��n 	(s�%��"�L�1�!b�������֐V��Z�� ʓ���D��"�Uw�e�A��G�mOo|[�tw��O5JNϠ�)�i�mp��;�u;���0zڈ��u~%T,�=<Q"q3q/������E�S�9dϭ-zH�4���Y�.�hc��꡶d�L�JM"���e.��	�eD�������ʪC@�d'��w3�f��.ޠ��q�~e�,`?�-��/;;�8/ճ��xX~8�zW�)x�'�|���I�F��"�M`ib�n+y�/��!B�'���'U�ɢ���H�i3(T
�jn~+w!u�'v��4sSv�s��T��`{D'�@)�C"6Aeb\��Y��龽�-𲫮YY���&Ni���I��܉�v��@5n2e60�/�:�Ts��,}�q��Cs*��y+R�� Ld�kzx��:�L����3���y�=)�Fm�n��u����MR�!�
��%Rj��mM�M�Qd#�E���k߱gKLw���Ί��(�aG�&�`�}S,k{�s*����V���]S�Fx�*GҀ��~�6�V���/i��JC�<�i�� �I�Yo��������2t�g���&. J�Nt�
�;0u3��XȇC�\���i8�u}���?��ͱ���"%��':��e��Q���,�S�u3�:��3Δ�Yt 8�8���$SC������J�6�mz{y�L�05��_�pE(w&=�������q��C	IQh%�|��i�B��a�:?qB0�(&B�BS�|���pXZ�#��xHj��Jߐ���n7���Քv�� ∷ƣc`+eǷ5-���3�u��j�N�z��U;��w>�(G)����d62-��V���H�>g�LV�%���>�
�5�d STbn��� )�;u�F�ПP��uaJ��S��g�$��=�U�]CB��`����I��C�K�qï�_g�,�f7^�7Ģ ���sX��d=?8�亓�E+U�p�e��L|�x���ݾ�:ZLQ��f�DN]�۞��=�ݧOV�e��7�I���Z�(�\������ѷ�n�9�M�4�KoR�Ů�fKk��UI�f!�1���G�m�K?�)�����y q�?|0�z5�juBCy1d��h�}P����2*��&�����~i&���=5�5'����>g&ϵȓEBy%U_���ƽ�]|-ǽ�~���g5Y!��6X�x-��W�Y��58���t(~�3����z5k�8O��a@���q+�4rE����_h�Dk�bIk��\�T�ę4�S̍�۽�=��Q����-K������_�UQ(FM�JG'��1߇~$���u �8<63c���j=:�Mn��9�n1�:�%��׆m!�
�<�/Zؐ2��B|۠�2�1�S���*���� W�I!�C2���"��qu��L�l`�9'��POQP�k ����,����>b!<
����۾�8���-8fZ�;�
) ����&�;�%���`����=���i{�vl�3B�u���~� ���w�f��/c ��#1F�戗�`�/F~�u�M^.��H��M�v��H��⎦B�48�k�qM�2K��.�8���t�{��=�aL���xD��gLG�]^�k�s"X!�+i�${w�e..��ncn,�����E;��� oYg���HӬ��:8�!�S�Q�H3K�����'G���m��!P��HFO�4T� :��G�u��λ��C�F��&��ϒ��e�6�p��9o�����,,�h������Q�h}0�����?��#\�C���C�y4�қ&'A��2*7jŻoՇ;*�l�~������AQ�K�<��v�������5J(���4!g����c�����[�֚2>����W>��of���|���i1% ����ք��Z7��Jλ����{?B�u;��!C"�m��n��ً_[��p�h��� q�.�07l�#��"��VȦ��tD�} �!�t�2���nō킾:1|n]��&��H\�-���)�=���M��X)��
�$�������0���fK�])�Abg̒!\@��Yur�#�а˓��&=�G*!6m�cS/Ղ��mĽ��+����`t�
�\���k��:.	�=!�rz�ȭ-J?��a-�%|�1����&�h���]^է�xS"�\��~7�Ee5����l��N���5M�&nx���Ŝ��x��ȺT�%�H�GXi;X3����/9@�Y�a�y6�1����7f�v2VW��0hU���,�OOz��f��m�N� ��r{g;Hھp��h�	|%|�17h���Bp���KZ�Z8��$a��ή��F�7��ؖHiy s�:;p?��#QV�<O��u�pxЏ�Y�l��h*yl|;�3T%��\�*F/��HX�Ո�.�'�Q�sg��>q�phk�C
�n|gQaV&��q������`��.œ�vM�oH��#¬�@X�K�hIH���n���|��)vF���.�mJ+�t�R&X;[�.���y�_����Թ�@o���gݽ`�4`}�ga��|�I��@�I�#��|"Xi��O��^Y�:���+&b�T�x���q*$�hB����U���0{�h�F�μٞ�;��m��A8��C��V�t�1�RSH��$�C����=�SuF�d��r�L�����Q�ts��c3D�|�n�m�~I`�$Avk	R�y1A�X|��F�xw;�|A0������=[hi{+�i�����o������$T�! �Pg3���)P&����P��c-�0#����H<ʒ �YNɓK��9��A�ɞ��~&����ͼ�MD�wS����5z���m'�\�J#O����tYή]�r��wǒEĊ2g��,�{�.�;3��َ<$���������N�|j�7�D�1p��9Xl�اOd���c�dԻ��/:��K�ߢfm�ez��� /s��i��Ƃ@Liq��O�������52�Sz.��K�o׾c4�K��l,XF������#9yMra���Ju�
��I�Çv��o|܉����c��w�Gaǌ���A��wP������m��8�nT�ͱ��j�yq[�r��Mk6EO���^JTX}�U<�|cWj��~����T�1����#�	E�-K�Ux�^d���r���@�nq��Xh�	)��~��ಁ�G�D�� j��٧��e]��n'����GT��8#ʷ����q��ݓ6qٯbS$Lv'b���}q�#q��c���q+piZ}�O�\�����q�	�`Z��2B4��q����I�k!n��"-t^a.7�5A7)�1���6�^0��P+��Ծ��9*7����v�gn'y�4׻ۈ����Ǆ�]2�ҕ����NV�Ng��5�Fs�$���x����O<;-K�{؆$#=�>E�G�
?���v�k����-�����Z�ޥ7Wc_W�o����vA�(�����}�C���#s���P1���p^(r�T�gP��<�i�)��A1˹;M�p^=��6N
�Y3�a8y0v�_&�7�nw��8����>���h�ޤڗ�8���6�4g p�6.K�RW��-\�3_TM�8l�P�hc��meS�>�g���S�$�Do���=^a&�c艾rE���w��pT�����[5f�[�� cկm�>kr���Wv�����Au�bL�gJ;-���l��®>Lq�Uj!�v��2~�}Ĉ�u��q@�`f��a2�$\S�z�KL��D5ӱR�qgI�f�N�?�;)N�Th�y��lv�`T�d�o
5�J���;*'g�6�tz		�D]\i˄��7���{����A����ϻ#bUwb�y�:J�����
p�:lT��e�1��=7RڻO:|��̓�։I�g~��J̚z����`�鹼(	�!��~����sjk�� Y_p���G���� X�[�� �Z�]&.���e�G�Rh���@�W��6��u^�t�,�֒#���b�.7��>"J�O�T�p�2��s�K��9)"�n�=�A_����㟆XV�'o��y�qAg�� ��\��h�/�םM:kǲ�~K�l��r�[f׉N�e�l��u8�Aܶar���L��)	s'>��c�Ht��Db�$�׎w*&��)��,��� �>4�����3�`��k�l�1J!)������k��k�Եg�� ��w~;�(:x����Ľ��1a���UCF-��1���LVW����KSdF����e��2��*Kݠ��7�
g�2�`�ݪE<�m �X������5h5�}YE�L3ήH#b����wH�EL��a���#^q.�v�S�6�I��gr���ؗ�W���|̀��5׻%��r�ٔ{���r�߬����p��Z����l��nޚ�-�ۤ�$U�B0= i�.�9��R�%b� ʁ�Jx�9�3�����"!���B"�'�b琄+���@ T��cc�����h3=���'`*�DWI
�!~�Q:�un���_d(�1W�3˓��yS�6�J�
�J`�p�ˊ@X��($�퍎�Lc�gt	�*;�CASc'�O��x��E��R��j���OF`�l�I5�j�%�1+A�)so�Tʘ&�&w��(���=1��gLm��)�x9w��}����o�el#�@���lWŒ/*�-��P"Bg��i3S_֎zS�g��L�-��=1�rxSY��Ѓ���{���D3�jb��w,�u�9.�U�������|5��s�J _��o�Ϲb{���Ng!�pʩPH����P�l�SZ���ȉyrP���,�M)�K
�� ���e���jm F��#���j]?0Azgy:<��}\�7�����v5������Q����BX�9�~L�h���9F���)��Y0
��*�������åp�'�������M�R ��/��`Y�JSe�-y��� Ҋ���Р_�9�&��S��Z)�η�6��s���6�#�C��yK��f��f �R�A�#�Z��2}�%���7T��v8��%)GW��," �W=`���Q~fq�C��3�v5��ˌ���P�&��$��:#M
��`��}��l��n��ԍ�����L����{Ԇ�Ůn)�<s�+I��M��ٌ�K'2����f�MO��/}#%;���b����v�#|>����9]a��GB�sC�1�_�[}}վ��� >�8@�;�"HZ�$�`�?�nUaR���Rט#܅�k5+IgIc��$�}��_:��]׍�K?��'�;���J���b���C��Ew�W�<�hv׮y/�Һ�o!Al��_�-;�{j����c4��!zg�W��
;APj�j&҂)Jٿ��K���ʩ�8�C������r��.�"'|	�sT�іrmf�h0xm|7���p���qMvwl�4GĆ_
���%Z3I���I�|�^���2K<��w�i��L�h���}��S���i������"��I���Ʒb~�>F��lڱ�kң�������k2I>�y5�fii>^�x��6�V������XW�YGs�Zb֒� ��W�|�uN�ǰH�S�l��o��X�d4�B?Շ��%��� ��8f �����v�<s?�d�Pb�8L|wA�0b�p�����b!��T����+�2:w�b�Л�q���
Z���!��]d�T@M5W�ka|桷�mV9i�9����$�䆭�}Zl�@��}j��Q�����xU���X��3�Z���$W8%P>����־�(�Ƒ�T���.<V�r�t
�v�?#FU�����BTp�0r���ؘLQ���W�$���2Y��qA~�nC��3����R��hJ�7
�"���