��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�rQ��7%gN���i��v1��(���:m�>���D'Ͷ���tur)���!^���p�NW���^��I<:�E����Gd ���
��Wï�����V������a`]�e�(� ��$�z�K��w��b���L_*�Io��󨒎$�����g�-�A/��n�\�I�z�OB�\�)~������SD8?؎:�;W
�����0�Uƨ����z~��"�qB��ཀྵ��<��1c1���;>^�j���I��ɑVs\u�(�5�I	\ڷ9t� k���Ajj�����z�g�D�_�a?�K��ؕe�h�M�y�
�zo��ĺӲ�u�<����GY��?rEnZ�_	��CP�&�z�;[HC�'�F/&��hp@3/ /ح��ƈ����a��)č�
�N�F�avq[��Q1�
K�R
�翯��Gb�gEA��A[��qOH���++�X4�<Z�N	<-�x��YXQ`�"���hޏ�R�W��]&��J/ \��͊]"��u�#�K%ilQ�V{Tx���]�Jq��1�L�&����䟝��!oN��ۂ;�xUU�F(Ґ}S�x� !ej<MZ�JL/fUlB/͸!�Z�B宍 v�g�'.zw$�f���c�U���o  ���%�l�[Z��n�����)�u�c/��l�㚴3o�b���r��t?��`!�TW�H[�_l�J��hY5<QDsZ�>��v�+�K���-fvu� ��%�-dsY�.h��D�DHJ�=�`L���xE��I?,Y�,�|�M{��@	��x���Oo���vNQ�ѱ<?�6<k˅P@�l=��%ԄQ���;��PD�B3O��5�f}u���zcQ&�Ҡ?�	`/��m�|u>�yU��F�=���d%�Z�7S�},H�$�f�YhD��	�w
����z��U���bl�d$d�s��MT7�W)I~�3�sJq��^v�zUD�6#G�#DD��J���ɎC�H�śo57`ޫP�~���Zm���-Y�_�1U�l�(煍aRQ�k�T�o�Q0��x�P\�Ŋ$gU���:YJ
��uW�ǘ��;V�p�H��:U�v�x:��IjT�-U�1��{�:��8p��J�ryNk��X��l�Y�H�>�L7V�@�nG�B�w"���䓒�i�?��&��<��>����WI�+1�+ؿ�x}Pmqz�тr�p*Na�6� ��AY^v�F��P�c^��'�a&�������RH�֯�.u���hǭ
W�~k�����~$|�[� }L��{��Â�k�B=_C�l��9΁͝U�l�4.�X�ԘKG��GP�&��)�,[�f�V3�zY.��$6Z��G�%a���w��9�Ə66w��a'�����zlI+۶խ���Grի�� ��:{%�y����:��S���z�td,B>aH�ʭ`�Mݷ�����Z�A�d�M�gC��%��xρ���q&o�>���2Ry�ɛ�!�1z9ə"#��Sg�boc)��ɇ�a��Y�Ô�n�#)�k|�di����o+������
!^����Uu�y�� ����.u�pM.`Z����%�|���+)(���`0���pO1;�F�!�"ܥ��2��{ǣA>Z�	��YewQ�Z�<JC�ez𾌺�+���0�h�詎��g��K\(IM�7��v��Z?H��[�V��Q���eİ�+���ߵ���L�z2���F��v&�P��[z;�3>2�x�Κ<m}���dx��hi���J���:����d��n�ـT��� Ȫe^X9��n��UC]��\؁۳)K�f⹨{?[F\*%�)�~���ęw�N��8��Z6x�e�=,��9��i���\�%{3���<���#0.�,��t��j�?`�}�A.;�bI
Ցq;c����.]��H1D�\��(Е�Z�g=��k��f&����{�	�o�bq���(�	�@����Y����u	B4�f�i�-O������|2�|_}̞5��G���W��Oˎpe#��R���,��pˈ�G�~�f����&s�K�>Z �*�ȎtK8��v�<k4��S��J��D����{M��h���P�<>}�b �GILfeɐ�[����&h�!�����B���l�>7�n�k��
�db8ǿ�1ALi���]�ي��� Y=�?ج^��<"���q:�k��@(��zœ�3��p�k���D9|r�`#
��$���,�	��'��c���-B�h"����W�H�ք���v�K�*��5�w�����,ݡ%���8��<��<P����{H���i�[�+�T|�cUt6�{lkL�p˦w�'&dp����G$T�:XKe�ɮg���sĝX�<��<ΐNzPfkT�8��e� 9˂�;�7��azq�P HUmK��D��۰HIVIY�9cq�-�i�X'��u߷�\"�F�/X��Wf�o||Z�݉Ӷ��8ؿ� >��dT�(�L��zگ�{��eEZp�'=��0��/�Eկ�b�>+��� ؍�ƀa�
�XH�3܎�3J7;w�L�O��\x'Iri��'�*���ݛ�˩��&��Hb
�W��5��[��o�4�"� ���x"Rl=�D�����I9zb|��O�*`W�dZŞ��1�dJX6]:����N���y��g3Y!����6D��,���7}Y��C��0�}��)�����8A�>�L>*9�$����me�uk}X�%Z{�r��R��~2U�cV�3����Y��β'���|HgX���,օ���T4N�� ��͟v�s�W���h��*�w� 	,���䠩D����1n�+���������|�6[�%��a�A�����o#W�l���Ǹ%�@y�U�e��qG���5���Ar_��o�"���<�z�ѩ�f�!H)��ύ���Hx�HI���D&��B��:�?���.O���,.DI��2#�a5���b�F:�����ِ��Y�r�jR���z�:(���C'�ᄟ�`������l�V����nk��eo�F5?~O�&=c�ďp?�n}k�ޢ�Iy����(���ߴso�]�D�ԕy�O��jG����x �4���GO[����P�Z @\����\	���渪�����[�������BԷ���}���ͰC�`RT�}$'��=k"��8���э�g´.��+\��{8 uT����V�Ra��ªw�X+B�Z�������dBa|a3PE������o�_`/����U�}���[�֊A���md�kKg�O(�0�u�tlx���c<B9�,��[��o�~*.s��xu��f�J"@F���Y�ǉ���q=?� f	u|���ͼ�5$��[��4��7�0��x��Y�۬�|��R��R�0_ ?Ѐ㈛��2��#ˀ��w1ZWL�A��f�aub���i,y�@��yeu{���yQI��E�/6���P�9�<�4՘h;)�帷�_G���@��z:۽���@h5�a��%H�\7My�:v�rLM7M��[����59i�<B�q�qu��H��-'��z0�8ᰳ�t �
�G��N���J��i,�O�� ~V�T��\h�1j�������"{k>%)bI�) 
fs\+�&�Y��ʁ �{؎)c9W�&Eq���]4sh������e��[���r��͵���yz%^�]��� B[`��4�����ώ�� �W�]�b�Ӻ�?*Ab����$����r$�	s����!��y�/٧y����x޺q`�d�@xKi�ݳ�/�j8�@�D���o���ŵl���U��Z��,/�䃸<M6 P"Z����<-R1Hq�{~`�Ȩ�����ܼU7
T�#^���x$�'0�g������MCC�K@�$�s|h��,D���0=�w?���t����~"g�9K-�c&n�X���:�59�u�հc��u�3`@�7��tn��F�C��N����u� �Ju���W�w�A�b��Ԁ?�DԯV8��M�Ei��؇TT��I�z���=�^M�8�����x��Q��$D����jr�P.Z��3�����eH`�q�x/!�ȲK�д��w��)�C"��OjԷ��CgO׳"����Z0�N�������_r�VȤ��z;�9�t[�.��}'>�k���S�[jj��z��-�Ó�[X�m�#Ou��w�c�k��4@��D��M&��^����f���e��w�?+g�|i�z8J�ݏ���A8���J�{�mt1��\e7���6
Q��D�v=b���[�l����� �E7��s�༓V�K{��j�m�����cLZI[a�?H�q��c�� �d+'nd��/�>�CP��.�}��*��4"��G%O���ۗ�p<��{��M	ٙt�g�T �"�rƪ��,R�*n�`IH�Db���m�2N�*^ \���۟ �V���1e@���?��_)�� �/~��d���n����z�3��G�<���k��=(:R�й��i��0E(�ij��cJ0w��6���b��1G��6K�$	��G�ȉ,���l�b���� 7�@�Kˋb��$2��ŕ��"�p5�7j�qI�s���3{�G�bKB�4|?B
�.��R���HW�s������j��Ƅ��h�����Q���x���}�'՘��E���%�ZE�b�ն�����D��p�7�#[��+4=�OܕT_��+?��0��z�9H�#faW��K�jo�1I��?M3�{�[ |�4�(��9��̰�m�L&��b50~q�}��-��BI�0h��h��%M��||ث�$�to5-6�>����,�,��7��h{2v��J�i��b���}:�ϬA�l�0�KKо9��"����Rn��0T�aWb�ۥ�����x�P�?�q���޴k^.�ϋ���K���f��֪�9�5�"�m��<&���%4��N����Z	 r j� ��r����Ti�h���c@�hR�/ *Ͼt��"�X�Wv{�a$t҈�3�_�,Qi�g��
����&�����w\��$،)�V�;:� Z�uw1����A�(U�W=, Z���xF����K�r��[�^T댶��]a4}���,4轄�*��Eܓ��Ktg�P�,5rp�3��[h`�Ig!)��i}�u�ko+�[v�>�l����O��e��N�.�����u=�,(��Z�M���O�z��ЧP�0��/# ��;���;Yy`�
EdTĿ��yk��D���W������)!�꩙��r��)����,���j2�pd2��8K�6���*wH���qHT�%��ɝ
�����z��V<��ғn�-hS2傇��M >R1ig*�0E�5qZ'�� Q�#<�y��1h�7ģ����`˔S|�/�,���.jy���2�7�Z	�$)�#�����hH\Y���O����X��9��d.��*�%"�l)zE�fx3<�.��?�a����0���.(����k�d���βW+�L���\�K��ln@�Q�`�v\Jc�$��C�,o!�CI�t��M.�#�F�ҕ��w �Jz�����T'����Q���-2i�^߱�����xǶ��7 ���j���:���+�w��O��I�H�Ma�M0�&n�i�di�Qo-AdD
X6eﺣ���]�翵�y;U��"�Z�;:l[[�S�[��M�d�c�R��ݟ�>c��g��A�#!����RxG�j٪o���)�I�a��ς�Е��ͦ��wI���9C T�A�� ˨�w-�X;;(ouq;�ŹI������/sv4���c��:�����'?�����H���A�Yzϧ�	R���r���d�}0�_j�V�I_!Y�g���9�dC�v�^�V�73�;LVH�jMv�T�H�z��Ғ~��.%̝z��9��5ץA�%����y �4��r��#)L&�_^I~�SmsF5�*ADʢ�����~&�4�bg�H��r��z��1��i>��ݼ����l�Py�.R�7�v�"���.SJ.��R	�j����ԏ{�*��]�`y�X+:�f2�,V��	��P}�%!�%[�f���SI�t*����*(�1�k�%��M�{ia��n	���7#����~*�D"�޷vž�{�+���3��{�[�-��Zd|�l�S�(6��A_�����£�Z� �I�#}G���_u���%����"����=����*ׂ��=��Fg�����:Cڷp���}���w�b�mʃ���ud�Y�>��k+��Y��sY}�&"@���6k-S'�6Z�%����b}C�_NgE�q��� ��Z|� "��Z�]�:���{��\�)T��LX�q<6]ea�J��}�:��\�qa�3�ԧdN�JTa�o�@���)�X��i&��.�l�Z��|Z5bQq��0�5��i�V1�ux�F�tU85ONK�Mڙ��rw���v&�3x�
�u�HR��/��]<�/b=YG�����Y�K���0u���1C�X6�����z)�44@R��B6�P����Hڈ=��]CC��zd� <'�:����5wB�`�s�)�úˏoö�H�DOl�th���4T���)�*H�x�x�z�1+�9�J��%,��%�wk�?x��a�h,]ݹ�$����U����L]�;��e�f�|�D"i���D��;��+�qp$*l�KŦ�s��nh|�������P�X�{�"�������9aC�mz��y`	p����!��Q�@�6�4]i���u��jc�4��O��D��d ���	ĚFE�P����~�u��D���w�:�F~�I�$6-�IKu��ea�62���C7�̓9�ל�D_�£�w���C(&��p�z�#�-u �'�S@�::n�֊���\j�������4�Q�&�A�G� �l�M����jT�L�$3�������aݎ�ή��F	nD��;�/x�,�_@��hf�����ok�C�gOt�2�՟z��Փ�q�e�a��)e@���"��`a�P���!�����)k�C��1�q�L.*3�HP4��I`ڱ�]��� ����2�&TIG��t:n��Tr9v�W���J�)"j[tF[�!�>}i��a�fk_�a1��L���ҁ�U��Cj4�b	�J�D� �o�bQU��WJz6g^�5f�JB�o�|��.�F�"H�e]���/��+u� ԅ�`Be<9��;��!F�12p�C�9o���{/� MFޔ����9��b�����NK{�&�q�,Ȉ���c}�.�&3�2�T:R8��-�{�Jb(���Hy��lj������ё�;����*J~�3kI��#�_��D�����Ƚ7�qPƁ�OF]���OӼn���L��A*�7 =^�;��\�9����-%nXǕ�QS)�|�N��˧��?_2�r�͐.�<N��C����� ���Yr������7O]�a5�p�j��Ғ�$�H�n���P`�
�	�Gџ����4Ǭ3�P�j̋�i6�đAkb��F�Ƨ^C`���Y��p3�I^6�"��s-ߖa�KO��K�V��:�^;KK���A"�7����)(۷��/,���4�	�pJ4U�x��h��n�ꔔ^<����v� �jf�0�\C7�Oղ�ֆ��.- �٥�_��`z�R�v�o`�@/�?o�g=���@��deS�c�X~m/U�����q8�����Q��)�b|��ٍĺS��"q�Ͷ1�������N�c��q=U˱�!yF�c�,������n��ed�Jj��Үx&Z=?������i�����P���>�#�cBn���+E��BHҘ���NN���@�n����L�"�_k�WҊ�%J12j��8�����z�jV<f�}��]�<��:�{��� 1�U_�x653~�LM�fU*?(#��&X�ɸ��� _ah��CH�v^���MP'2��۴�^7uM*jGK�겹�,)�<������qwEJ-1�p�s��1�./J��⯮G?R`wl��ƔB�?�����y}�IJѶ�w��. tq>�����]��j�a
pKe�~�� ?�u�6�o��Gv|4SK��\�qѹ��#T\ԲSW�Vs�@��LLb�r���1���K�AЂ����Y�yi�����M�ȝd5�k�ۿU���������fJ����c?nH흽}e�/*iQ���%�X}�ˬ"����[ud��m���r2��?|e�"EzN���0I��Jʭ�<l��HX5)u��K��;˔L�Τ��=�=vE������o�J�� ��M��"i�L�J�W��4>y2��Ë�x��5Ѻf����t�O�*�[�6ʢw,"�(��W�n���AKk�^�|���{�P_X���(5{6����`RԶiШ��cr��<l������j�RV����!x1��D�裉�r�1��'�=QD�klZU�`��ߜ�i���� V!+]���;��t�o��m�g^G �qՅ9z�ysZ�3��P^yMV\ؑ�����Y	���U|��%��?t5�M��
>rm��]�E	\a�	Jĭ�OWf��v@<���)�'�`#<�JK��7^���{��X���Z4,�2D,��e8f�z��o������k��j!�ڍ�N@����:�����-y�v�Q�\����6��g��4SՂlu�ѵ��R@�&�e�-sD��GW(���9:ċ���@�i���c���W � ^�aPY�fi����:�}�����g��������=��V�h�(�Fɦ(�����<��+�`�kS��CR�G�+�}��ݱ��n>�������Z���&������A���wͲu���淟!#s*����Ӝ�@<��}p���t���3۰��s):+S�0�o3���P����׃�_(��9_�y��)O.r�~�y\|خa�v����p�$~�rMl��&��t"��w�ɮ^T�f����n��y��3��h����Qm�`��X��6B��1�=51I�&I��� q�V�f�ʂ��c#�YS<+��@���s<�,��ui�b��n���
���Y����mw����^�x,��&?��Ə=?�V�#��T���+>XH3�@T"uTw_I�ĥ����FȺԖ��C�l�
6F.͛ր�y�����}�Ŧ�q�'u�D�kA{TM��𒲽�p����"J ¬j��G���K��#�PC��;�'�V�X趜����Hbs�"h�	~Xf�`�#8��W�v,���%5 �<�U��q5l��v8���^�z��惻���ʣÅ�wg^|E�/�U�đ��n�.�K������D-�����ƓTpV���?OYmf�0J��|���J�0u6�J}��c`gW��,�q�COBܓe���T��S~w]bn�If�4�Kx��s?�8��%��`�VJ�� GB�z�l�[B�,ܦ�dG�7n ۾