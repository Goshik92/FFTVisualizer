��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�����mHԍ��?��͏b��r�-�R�.�Z���Zʲ�%����A�C�$b�ru���uo7���%��;�F	��ž^Su�{��[ik��e9�f��T1HA�D����6�ug�]�6��+*2�6jZ�W�G.Pj�MY���	GWk�fy��H�~��P�ө��̂+g�oG�
�t�BC$��Z���^�f p@��bN�p��V�S���VW`:�9��,�rkLp�,d���ٻΥH�����i73~���w,g��6��(+�P�	���8}O�b�t�Kt&���髪��@�ܙ��f`����%5!ÓCx�2i�?� ���Hm��D�A� BZ��n�1*H���ع*�x����Y�*�L�(2���)���P��s����(�}��C�ʊ�R^�`�wq2/��n�<�6�9u�i�_�	����r�k�υ
���7�5١H\����a��n���2�`�6(ޒ[x���^�>���=��Q��{7p�8��A����t�̱yHg>}�!����-5��cͷ�,�TD���6�j �.����%1��[OҎ/�o��'�K��M%ۓ�#��-�ڴ@�,�CrA{��*�������χ�1�a:Sqa�x��U2��������:�1@_��٢���zx(��QA֊a�ۗ���u��@d9FN��-Ԏ�9G@ �YGjk�(��A܉w�3C���]�����7��>�x�_�U�Z��<�w�F,$ÜB�����:/h�H�W��r>"I�$w�Ѣ'���Ο�ul���BP! Z`U��X��K�Zs��8��B5R���<�4f�
|�'Ưe���;�
�J'�vs����~�Xn�0د�JG����8�T.'�5�G�0Y|��v��k���|�
V��$�|}���w��̒�I����!��	�V����@ꐋW�v�C�b�2��L9�������L�Aa�Y}Q��ަ|��.�tE�>-��Y�N_����~�rOuGx��GӜ6+�-?�Z��~�xP��k�M�����T�V��er���&-�u�J����O&1�+���ٷ_�L�	���eS�;9��쯄�-��O%2d��33?Q5��?�ܬ���\q�F�\�$�G-����XR��q�|�	p�<��nV�*���@��a��3c�L�����W�}��H���������F1!�r;j�{�h�H�U��mY��0�%���9�GCP�X�&�g��������ސ[:ކ�N�ֈ�S>;.Y�y<���S����ٸM�B�y͔|x?�F�;��fa���N�d=h �5
U��_z�zf��K�D����
�����8a׆ߐ���J4�f����Ca�R~.�YPK�(jV��B�AD\u7L�#c�V%r4n�Ѭ�V��G7b����ǁ�G9z�?=���Ys�Iꌭq��y~.%�������PgZ��F�I;U��(�3���tߎ�:n�s�x�z����`Y�c8������}0�G���|��+:8W@v6��������WZ/)�f�X�K��5�܄ތq�cJ��n��jO�CM�E9]�zҴ��	�{��Gd�`�P�^���Ǔ��}d�����P�%�<��I��ՠ���Ӫ����^�$s0>��/uE	B���x�V����i��Ta����!:xw��L�=�R�K�.��ACvn��|���@6��	�k񪌡�	���I���Ⱥ���+�4)$��غ�A�E�%:�jW�Ya��W|C^E�L�w��ԸCuWf[��l�9$_�Ȋ���������/�P;��r6(.�����!��q�L�fo���T9q&o��{q�Z^c��~���[q͌B�qt�Y�|'o+@��+�=��D�z5lxu�>�u>դUz��~̓ɃN4 �RC�N\a��j�1�s�礨�g�RŖ��I���h祏B?�� �ъX\ƶQ��@=�G�@��C��H�J�h	F��T��3�|�#��>��8���ЕCQ��0F|R���A�w`���I��<�}Q�٤����@�m�fT/��~� ����l���v�h�0��-MBet���o��������ԝ�j�G���nO��0bZ�	krT�ùG]D��A����%�t݅�f�m��ͭB����ha���h{t�xKI�@�ک4�33��1q:q�βp�
%�<Q�aX���BY9�|9�J6-ԜI�5Ý���X��X=���U���^�{[���H ����^�w^�$��P|vW��o���jn��nz,��;2�T�N�ƀJ�C�%�9��~o�}!7�����h�T:�t�RXBFy���n:D��S�K����Ʀ܆��\T:��w���w��.�A�珲����͙�b�.^��|��i���X��R���@y�+�N��� R��(ѳ��J��ǅ�5�c4	J�s��.�������"�zY*��D�/��vO8�����=ґ���7���K��vslx��u�[�����\�Ƚ�oX"7�^\Z
�����}�bs�O-`X׳s���P�|y�:���P����$��p�wVւϯ��-�x|�#�ˏ��X��8����PH��X;�'_���g�V���-�$I�؇|ɗ\}����{/����*�C���!���ž*q�'Pz��7x��@�����M��30TIe�DgY��ds����ĐX�@�O��
�	&��z�s27����T����^��+�%Xw4�@��Im��5��Z7�e�-��˂��kb�g���*���=Y���yvd�$��3�A�o!����q]ϐ��o�������P'�9���1����:t�=���/����J���%�|H;�e�H�^����/O��9]&�N��8*j��c������mH=ߴ�v!��.\6n@9kw�Ɋ�)2a;Y�ڈD
i�q�$�Ŗ[��E��v]IU�֦�|�ɉ%��ݵzǯף&I��"���o���Fh�f����Hl	�D�oK��GʹHr���G�9�R�x��e�uhk��´���O���Z`RI�.$�$�Kcu)���J`��D�Vq�Adݪx+�Dt���%����q�K�р�iҶ���ٻ^�4�5 F��	�����1�,�s�s���,�[�kl6�r���5��=�6XۅO���G?�2��8�Ԫ�چ-?V/��,�O��őRm���O5�h��M���Ss���,���1�G�*�o�Z���93;��ѝ9��'��AҳdW	�\�)qN���@��������M&���NX���ӕT�@�E�¨w �
�����b4�2Ŧ����g���=;q��W�&��Du^�������@�'���wrg�՞����O��Mr���\w��������qy�-&v��v��屵p�uώ��Ҹ|/����/$"�T��D|uD����e��x��fޏ��:<G�4ZU,���e�S��6���K�[����g��A��@5l'��fUM�U4��>>��~%�O�Hk��~A-��I*����<�>&�[�H��B[,����k�T��7�m�Z�*�L�ОҜ
Ԗʋ�5�~%����8:%���_�_�>���h1�`�y
g(�"��Z"Y%��cas��VP��ŧ�×T=M�\��-� >��W�TVd���I�_E����[����w_^09w(j�ĕ�Dsu:�7�ek�0�:�i`JЉ��Q���4����G��pEE��:��FJ��zh�\ OY��؂�d^�2_�rr�t���r�/�Y�ܛ�ld/ܟ0��@4Ui-_\T�21���[A�k���C��DF��z��w�0�uF	�_5lrk��j���pk�։��գj�D����ꏟڤ�x�-�MM-dJy�u�\��s�)� ���'�0Z;�/�J�
1�W?���r��nZ	|�S����ǝn�K<(�drsI�2�a�ϻ$�S���y�;�@=��"�Iu0�f�sH���?�L/:hx�-�l"�q����t~u
S@�Y�Zu�.8W5ǽ	�|�I�Г��b��أ���ia}�|�lC�1����;�����h�I*
Eo�Ѩ���"�4�b�!���+$���#xpT�	-��v�|zф|�z��V�������fT���Y`��d��{3z{�c��MY��j����w�$��-��Ѕ�)�m��q��\���?��L�,+��ʇДh*屓�Ӯ0p�hJ���LR�l�qVa##����S��_5����qv�7�9/�X��vX��t�����dImC6� U����W�ݱ$���o1�_R��}Ր0_������#�|X%gM�'�%��{��74_�|gG���
��!��1�ha�dJ�?R�J��R��/�ٖ�q�P�ԵfnXf'��4b2��.������*�B�lE�i���K�Ǵp�?��Z�w��F\5����,y�K���꟭I"�iE���9�j/����� ��0���1�)���;�0�����c+#~���v��f��rQ��!������K���Y�4�^|�lM��Q���s�`�&��+e�$	)d����M�� F�}n��M^�5h6H���$�)@��"-��"V���F���N5V�T��(���k�s ��?�<U��ء޸��):8~D��
�f�vWA���1O���ޔ[��K�+(rE��,����O֭�Rwǖ�R��j���R�S،���_!+`S����!�y�UhM���<;���ͽ�B�{�
�zQ1_ʀ7�݇o'��5�^~�Wh�2y^�;ǌXÿ���?����Γ�>��W+n�ZF!q-�j &�IF�t�ooCg���S���e�G�����F3��(������gX���+�P__���4gӥ�V��+�δ`^��P�t8�2-�K�!�Ը�B�(��+$��hh�ż���s=����ߊ��|��T�h�)��.�1v�c��¾X���G�V�C�<b���8�nEY�1�(�&����t�R�52
W�&rǱmZ���h�
-d�n��6;�*�b���1�����S�_�1�*3"�v�����MX"��p�T��:$D�Exq�\u��9�Nu�i�MG�KX���7�z�����۞q�M��`�Cb�99d���|�;x��E8X����> b_'���N
�qD\��+�{;}Tc�%�M�*����y�C[��o�Zӽ&WW��,����TpXA��V�ؘ��T � �6�V^�_*��2��O������#H�����A S!*B����K���e�e=�ǰ�>% I��<$O�В�F���\MM-���As,�G$W�%�S\�~�(����"4e�7�dw�p�j<�.�_�S��r�@��9?C�G���Ώ��a|�;����s���h�Jؖc5J�y86q������V�gc�uǾ��d�!ck�T�U=Z�L��?��8�Mf�oH�ؑ�Υf$�5`N�Tӯi�R�H|���C�D�lm
o��k=���*D��(�l�|ϮA��4l�m��c}W��(
[N�j�C%îE3"�#�p���0��+wg 3�����iT��8E}T/`&�k[o`��^�I%�W������6�?1�0f>!����I'^�ݶY����G���b��bHZ�-���<cNQ���h;�f�h�$C��~kUG�����B���.�jb���� mH�o�Ju5�]E�nO��&b��S$�Pba��d�T�})7]W֧�F�4�L�G������O��7!�����|B��f�7O���=�Jz3F�g)��k�!	���usa�q6 ��j��ׄW�!DC��/���۽�ۈd[�~|��R�`^p���
����g�S5����0�W�=���{<|�D�{����Gx�8Aj4=�[�/����n�M��w��(?:�0v�-ZK�[���a$�yb�[].&��_� S��R�\��#m�WC����)d&�Z-Z����l�:�b"]������#!ѷ��|!�q��n���
����/>�#�� (�xeG�ߵ�����zvv���7Q�����Pf)_ͱ��/s[8����o~����%��)��dZ?Zǳ�'�I�7+��
v�#A�
��Q�D�<B%���[�ݨ<��q��܍ћVz��0>���)7��� %��U<�F�c�:��Mk����}�٭$vl�����l(sj k_�>�3vϒ�ﾤ��&����2[D�QXq��Oyh�VZ��h\[ǟE�H��0��)��V'���8>4 �~~S�_�	cl
�DP/�M��q�z¾w.���U-����k0a U-���x]�+i԰"���hx��94�� L��ae�����E&� �ԕ����g�5�嬬&P/&�~#2@�A��O,k)+_��/p�<���6���[�V�舾ȡ}��i���w��@]c~�Uo�Q_U_���>�X���mW��C���3�:%�N)�!��T��xo��ѣ6�����xf��h�c��^JS`]Y��6r��ì���fӯ 
���}k�8F�c���8@�=�8J#(8�7D�Ik��/��">o$�t���a���Xb�ђ��},{���+���g�Mἳ�J�.C��%�և�:��8�Tz��U�,�{��5u�0AT�e�<[�X|4�h��ږ�/[`�mG�s7� #U�S�՗2���"Bb�4̈́��s�M#�$j��Z�z@�5-��RY���i8��d�Hb~s�Q8�F�6�>���w~��(����)�x��/T������y�u(�ڦU��>$���UT��V��f:&�W[�WR�vN�Sүt6��*�5�
L�0���x���v�8�k��֟��Գ�	c�%S �"�"�� �m�л��u�e���> ����[�07�h��xVUuk�"̓)=��C4��TK�y���QL���3���a~�o���3�;�kkg�*�-�tX�p��A�B ���#�*���z+cqq���s��
�Օh4&�/ܶKf�vNt��]�C�Ib�8�$��O�-[:����D�{��	��#[�n�fuAT0�iq&�`�[��[�R�-�n�W�[�U�FI�\W��@윦�k��?o�o���� �� p��܁���m<mև�Zz�ޚ�[dG��˕Ͻ�ғ�6��]k�%&93x+� .5�P����?���O~�����G6��Y�?�{�i����+����戒�g�>�/Nna9�Ǽ�ߎ�|F�¼D� Ҷ�R�utf��3��/i8u@`9��Ru�1vSn?&Ó��v6:�Z�t'ŧVю��A)U%�+�lH�����������L��X��λ��'�*+McV(0���"�y�AE8���%Ac,nͷ�M��猈�B!�y^縄�	2m�tBQRԟ�h~wl7�}х١�*��΂�3I�&�pz �{��Z:�� ���9��e>D�s ��s�%h؁�w��⼸�@���7�}��<�qװ��"���]�D�I2) 5P�j�ۀ���
��l{Ӭ�[=�
���T�>u�Ne���9gi:�2����P��(�I=�d��0 +8���r>�Xg P,��j�F�mv�[y7�#PS�|C�,����.~�l�$�l:^�j���wXv���G�h�k�
%�0�`9S ^Y�P����^���AX�@���J��,~e
�:ZIem���h;O��W"o���E]۞�)MPj�#	@Y�d˯U/$���O���5�,4/i�aW������1f;%���<U�C�-d��8o%p����,����H�CM,��ȱR��FB���������-�c�h9n�k����až�&�G�i�D��]wD�q����	�r��@ �r��NW6�צ�n����.��p���cEH ����B�P���R�����y��s����1�,l�[=�\�o3%2ղ�Ю�̈́�7��q��U9�=$�W��T�M�:������<��o�oE��6�e�6!TC�(vw�K����(�Jd��>׈�����J���k6`��a�ooHS��S��_�+���Y�����h*�j�8x�.�*	�9�Z�G�Ǹ�M"(������8���$�y*� ��l5����.����c�WB������n?)ɮ�pXE�����!7g-��jҡ�/���g�J�2N�R���&�qBrT�h�L�_ ���ͥ�5�(y��a!T��!���T� �-�5�W�'�2��3(v�5t�����>�G���w郲�h�÷j��a�3����I���ɥ^AR��)���;���ĎƎ�`�Z�5�<s~İ��$"+���)��}w�v�{����1�N95V&BT��E�CD�'���Z봭��p��o1�a< ��Q+'ڸo�㫐��)*}�y�̲�ξF�8���&�k:�5��E��M�WY�f�
,�L�99�W��"ٸ�7���/^�c�M`��%��Z� 	n]E��L�@�c+����[y���e؜�_�c:�* w��s)�7?=Q6�-�+�Q"QDqɪ��
m)��� h�@c��%s:@������Y
���F_R�{\/�[ֽgy�M�K�Q��0-�-m�i�[�W��f�1�S߳�Xn	ۖ����c������t㊟B#���.9��!���_��N�V��	�u�T92��Ӷ�,��T��p\Oa�z|�C��"��</w^D�t�8��7S�嘪�:��� 	��>ySb�J䘲�-Z^n�=
 �(q�U���������M.6~r��v\��Ww��@>xo.�c�������Ɣ��>>ߞ�5�+0^(����P�������G����8��@2>^z���3���Md+�� �K�݃vȡ�@�G�ck+�g�5��uX�1;� =�	��o}_
��������
���h�8�g��^��M� �����p ������0�~	a��YfQ	����P������" Z��%���?�e&7��~����J�tf�\2_��^N�=} 6�N��v���Z�ZȒ�qN�2.LٚK�^��K�g߱�=�$��N�%�IVLA���Q0��B�s�[�w�&�����H��K}|���}�VA�d2�M��wb��<��}��jE�1���]��0\'�i��ꚤ�?���D
�:�
�@N��$T�]^/��'�����{O/���^i����/�OdE~���В��Y|���e�r�����g{��K�j���W�ry�Q6n}wR���O\H�E��j�.��R�݆�����?*�,��^1k�J��t�Kk��}���ƍ��bqx����Y�ա���!$�s�w�����+U�e�D�����ևte��Z/e������������HeD�W���۽�ӧ�s ��_v���t���ԧ2&%�Zu Z\Hy�G��4[g�-��Ǆ�H�� b ���	em�B�@�� GV�rs�}xWÉ�J47	���n������F��{��z��+i��պ�oI���xOhS���H�6Bӣ�����0��p܌
gѐ��6��o�D�e�;(�R�1�J�f�df�L�������)�S�4N�CU�7�OA�蠱
�1��o^���>H��js�J�*�pd2���EX+��q`�lSrPX1
�v)
����Ƶ�f
,�紣�}n��h�͎�g�����:]vgM�W�em5�|�TՋڜ���1������e�Ԟڲ�z户�����:��c������-T��\�`qo���
��In���Ȫ�]~�M��I��eC˞�)
���#��(��^�>�6)S�D߼�L�]��bFl�L��{����e)�y#&��k���qN-),D�ۆ�se�ꡇ��_�%D���d�4����=�Z�h��e��Ei.���KP$t~��m>�7�'�O���:i�p�X	����z.��)u���PgE�]L-�̷g���
�bGs�CMS� �F-�x�c�,L3��h�.Y�������[�n�s(_�r�������|���Х�`�s�B�ޮ�k��bg�=e�37�SFE ��bإ�b�`�A�l�o�T{W������ ��i�S�I��c@C-�@.<P(v�B`���� ;`�CȜ���4Bv.�c	߫Q�-6�����r�[�EG��(�dҾn1�FMTv��ce�����k� M��"��X�������9��_��� q���i5���]������'U�z��4�����Pr]sV�r���q��68����ܖe�cx��-U�!�����`�r���M�z�seCȠR����k0�t���mW�)�vg[D�����俔M�Q\��J�����%�
D�@e,0��� ���	���+��&�.t�K@ш�t+�A�a�B0"=�[�d���&.���_�Z/;z���,�T���U_�,O>���F�bi�Ǎ�4�_�@2?����BYʃ��C�L��sI�h;��>�iP����O("��cY�@��pSЀ�����k�W��Gf��䎧��N�a�Pw2���~�ͼ��4t|�D�5�/!!P69�5�f�Q ����1{�&�K�� ؂Y&��NХ'�%�ة4	���8Ϣ��9l���5[	ӌ�v��YC[Ƅ'wP:roV7�d8{?�ߋ.��Gv���{�-g׍Dl��U���^i�[fT�q�h{
ܖ`�_3��mtDÓ����2X*HT��g�慼/�~����4F�L��֢^}ccb^��;Z�f��L���&�)0a� �Oյ�����# �źQ\R����Y��7�����̀����/�|���-�ne��6u�U��
�S���L�s��lyh���/�jj&ZEQ�oKe�����-
  ��8�?M]�@�q�7 !Nc�B�ެ8)����^�.���*�Pq[� z�0	@d�hG�p]��T:�u�KwF_����3�o�Br����^c�L�g�*����+5��~�K���¾Hح2����x�.�q��{4�P�8�?��y#�4���a����J%%�����@��f���\���Mz�x�p��q����h@�y�h�k�/T�&����z򥸩~�c�zPI3�t���i/�HH��s��8I���=Ʉ���!�͋���z���g`.z2�J���q�v0�6C,����>c����.��'��h�'��Dʅ}����Ó:kcg9Ve@.:��5X�d�&�!�d�9�,f �鷝���e����״h���]���?E��\q����X��y�����fb��/�-I�M�s�^��j��2�`3��4Q^c�J�{���1$���3����/���D�Ӑ)�
Q?��%J�V|�̃����g@Wܭ��	+�V�i\ �G��������jѺ��S�^���@��;!�g�D
��=�qr7��K�F;j-j��3p*M��¿>��W��]��5#kP��";�(�n���ҥ���.���>K��.�#�����̄��0h  �;s�� ���P�=Q3�A��y)���F�cv�)�0�{f݀7:f%i�#'���ӫ4q޷�s@�;�rٯ��&L�p��5�T�ý���^�T)�-������|��r���K�=�s��h����������t��"a��zNC��p/����(DJ1c��E�4�����W�
�g���ߍ�� \�K|V��el��Nґ`�2%��q)�_d�Ye��PK��Q�1~i�h2�ySO" �FB�N�-B�{�q!��vM|1f��A� Qd=En@98����
�#rB#1��v��=bL�OwR����Nio\�����gszs����ԍs�ȟ*��<��m(��`.�mK��Ta��!���/Sy��WvkN���Tρ�|QA��o��2���͍��H���PT�������&+W_��L�#k4z�Ccs-�¨J�}�IaUL�&ΟtY#4T��:�2l����扱��rj/"�Y��A)�.�y���;�^;��c��������\����ٝ���}x �V8�aAg���Ȫ/���g��	R���i���<����2[� 7T���P�T����?
B,䧴S�c�,h՞�K뜕|y8v���I�
cL�v���ZY����>����l��y��T�r�3|�|8��9�(�����BK���Ê�{7�	�FE�=��%L6@r�erD�X!���&�(>=��l���<�{e��q��ϻQ$�M
���^̈rb��x�^P�R�$���&��H(JV�.�����p��YyՇr,��|_��nF�OhNW��p�'�d���|�p^�'	�8�����-��?$-�o:�X����qָ��4�����ĝ#�kb�(>(f[糅 ����lr�)�^q�!���6S���*{��N3�v4%��m��~��)<�xv6Cp���@��{������:�]��]+���7�;%
+�~��������<4��!�R�zs��.yl�~,$W\�]�Y"�s$0��(� #߮~>:ޢk����w��,��N U����6`F!���[�nug�~����ܠ=݌���	2n�t,��M��)�I�9 >���h�'X��ĶL`Zg����v��V�V/��XX ���ѽ�V��#Xo�q�l����X���kCb�ѥ�-��`1�b��T=I��|��-�*CR�=���WȺ����
���U���0���v���̈́�;�ض}Q^��O-:zs���<���S���s��z�熒*�1v��E�5<�q$���E	)������b��j���M�ٟ$˟�-���2*l�: �䦒�}Uʱ��%�F4�L�WX��Ļ���wP����e��QP(�D��Gz��V�������XSm�p�q��\�o}+�U�: ��$^t���g[ħ�g�!4��4M���&��^��*�p@�_�"Wp��OD[?�pc)�>�-U�1�;���3/fm�Z�{��I 0Z���2��rق
^_(�.�u$��Z/�&ǡ�K[�P:h�z�5q�䱼'/�,0Fc�Paߚ��*.Z��#7?ei?��E~��;�����8|����Ynw���}�헕��}�#n)a��f=r�����sxN`)Wn5��[�wr4y�taW<� ���Et{+h��+8����!�zb*u�[Ȏ�R�}�D�Q�ebB���|�-Z��g�-۰GS����b�����99q�B�LZ��J?�X�@x�ۃ�Y�7(S����� � �IE��{w	՜tO�b�l�O[;�9,RZ�O��8�ȍX�q5-��������QP�[�#a}�I��7a��@�(�8���\�s�ۈ���_�U}�v&-~���ԥ)Y�4-ȷwj\;�J��켷�k�썧���'W���r|�Fp�iVi����D��e�v��|��J����RC�����HD5�HD�W�����0��H3N.~l$��w�a�@@���-��@<C2ȺJvz��&����e�l\��ޫ��jN�w�[�Ʉ�l�����W	�!��ؿ�A��E�OM�ka�@� ��@5k�	���P!_��u�E~�Yl�b��Qo� K\|�%��ĸ��ƨ�1����5�UG�N����kC��E$C�X�8VZ��`4�ӘSr��S�9�7�%�����&�*�]썏jt\0���z��}��x�YTq<�M��A��:;�H�P�����[��P���5��Ǿ�?Þ=����k�̏0z����T�KR���UX���1�~��%�ρu�b����&w�Mm�H����+���B~R�r�uU��uad5��x�}ኘ��d���4�i���W�r�Ώ��k�,mJf�?�Z`�8ڃS�#2jr���f�y�r3�g`PT]Yښ���ÐY���/L�/�w��W�.}@E��������N�� �zKM:�d�	S���~�2n��s�C�m,��Shu��w�C��,�<Q dE�ڇl6eu(�ʱ�7�Vz,k$��Bf��F����s��B9X�����=�c>ᅄgII)��W��ٔpG	�U3����Qd������(&9��������.�ĐXY�8�P�T��qU:�~�>\<�E�m�_�"x���"I�`?�N�E���"��K6'��p�r�OL��׊PS���E'�UTs���u���?S��a"FY�I�̫�c"�+)[�Ag�C�Ut�J"W����k*�&5�Onˍ�P��f��O�]  ����%?l����n�L5z��J
ݲN�.�[��@����ySM�;�n&�`]D���-r�%�Ӓ�Ƴ��`��N�A��YЕ���է���p��2��WH����Ej���E��7�j��ڻ���`���,#�����~�(Z�k˗��0�W酮L��ގܫ��~2�O	�!$b�B{���π[�}FM�������U
w}��:6��c%�G��z'4�$c�Ld	�2�1�>~27�:b�b��{ո���	�D ,����N�N�*�%��*Y�;Az��-�0�:?+ �&����+�T�a3�v/+��'g���?,�sT�� GR���g�t5J�/�k�
�c��q?J����_������x�r��z����/}N�	�ptd���LW����a��I��+Gd6������i�d�>ɏ,�N��C!�?H�Zp���2;A��_��&���〱����NN2SF��`���3���R&`<� 6Z����&p5� ���F/��	>��*�Jx	�&~r�r�wI���	Ԟ�mu���m���WԐg�u�o�H��Z=t�R�p6�/���S�<�X��BC4?�RB,M��C/��o̫r��C���F%�Z�"V�Rq�7��N�r�$��?�>H!`z���2�ͤ�мI�"ﵗ���m�=�N��[?��`�a�a4L��Z�$Ԏ\p�w����@�;��\z0��W�ݏ����m�I�y��[09i��ǿ���հ�x�9��ke4
S�1]��C�:9~�aY;�*�ɥ��id��L��m^��L)�u������x
zH��_r�X���9�0�E�P������J�z��rw��ĝG����把�e�=�j�D��{slfl@�i����_���6��Iku�������"�g��-3*�
��*7�4 ��)7 ߖ��<7`�]f�\J#8���?��9�͔feѫ/b�н���bh��5r����3��q��{ 0k��=z��e�l,B��]����-�5������L8n�-1p7ܪ�� 0����O�� w�`�n�2\j��`|�4X���d����k�2����0�hP���JUk�*Ϻ��R�6>kgz�1�$��C�*�`Z��
�Ǳp&k���q�9tȊ�Mƽ�q��#Ce�'fۖ�X*?���O!&xy2�O���K�<B�����oC�����:��up?v����Q��C�է�q?zk��ߠ��q��65�A��F��BͫZ�2�Ҁg��j3.�]&��b ��ک&���C ɧ*T�8G���������=</ʣȧ4�F�ͫ6���,u��c��f]��R"R�W�k��w+��<pVlP,F}߫�h��-HS�rk�7w�Zߪ�Zv��]�ʎXC�?W\�0�?+Դf>I��O'<��hoxO8}��S�lt����E�������:4;}R3G�������!ah�'�2�J4���	����y�,+0˗yN�Y��@�l�c2`����>�+�E�ze�W�[�H�?�1��m���������ֱ�3����T��}q��XfP�kHf��[:�as�&��-n1�g<�&T�Bq)_��v�`�i��酥�o����k:]�X��Q�m�� 6���h%�k��{��\*ӗ����bu<�$S/2��u\�KV�ĭ �u,��&�>E��zx��t�Qϝ{��[�>:y��inu��x�n����-{���ݬ*%��{�
"Rn �k16�����Qv�{�]lC�
�)Z=��]��Yw�"$pK�ɩ`:!h��
s��g���]��җ9���%�����	� N�k�FJ���R.Ȯ�T�/�q����1|,���.�Au�2�	4'1,T6���7w��H&RY���L�N�밡җ��[-2�"�$N?{맡g,$�H�B�L/��������&b���kQ$p�V8��>�~��U�Q�AM�$q���"2���EX�+
�>�t0׭���~�܁�I���1xx��cZ.��	p�F� &��8���a�є|�?�gC;�ac=z�I�5����&�_d��O�:>��!����8wt8��֔�|���ޗ�q3D�`�[f� C����k~/��z�c�K���(3:.}��.`uX�j���8_�s��\[�?�$�Y�K���Z:
���E/�m�'u!��8.�ߥa�}a�}�'�a�T8ny ���s ��v�H��.cB��z�/�y���^��S�\�h�~�%�7�F���X�Q��G)�w�%H2t�1=<&�����,E6�̋k������i-��D�ywa)B,�ʵy������t��+�ؤ��бdѕx�h�`.ZZ^� �6�ۡ�;@�Yxhf���D�r�U��V'0a�y��)̿�>]�� ��4�|tFX�BFo:���z#q9�ɓ|���랐�n�Bfv�R�o%����jhmg $B|��=y���T��_��?ݣuQ5���M��d~5i�2��BF�t(z��'a���c�lB^��x2}�V��2���ta��6�0��V����p��1X�d�ч��'G)ٷ�Ӄ���O^]��r��O?H&2���eo�0��u�	)y}z�)%N�/o!�ս����6���G��u�0.v�vO������d��PC8P-$�{����]�4��ow�=�%��z��{Q�<���:)��s���/��7j�"��� ,��.��¶��J�Nh�EJ*������Z��*I��92����I��`��-�1��..���C�I�'�X;�kZ��a��(�u�R�:����[6��4Xu�xM�Z8ݯE�;�"�<DW��fce�����M9�����c૯�'-���8*����:�ꛛL���r{�����̥+]2,��_�Bp�<�Թ
eM�fK�����v�a�
I�L�>/��U��]�7%~`���aiDQ�Ko�0 ����)�����Ep����6Ńݯ�њag�0ё�O �j䃰`x�2����#��mlg�')�<QMܪ��rx��YL�Y/�6����~
�8�6!�?��w8��e�SӴ�%yZ�JPu��`,��t��P���� �Xݷ�ٵv��R��d�+��ځg�A8z0��%m!���3�f�n�N����}�Ps�kjO���Q��߄��=��ˣK�ߒ7��na�(K��~�2oǋ.�o���5Z)Q>@�|%oݪ�6�p��J'��[ό�Aae�UV|�)&���s$Lt&:�z5���K�/\�=Ǌfu0�a�;�CP�jRd����P�]��֖�Y����2P9��#A����j|��a0k
�7̘+B"��|����|�~����Ͱ����5�j,`�*f�/@�ӟW���;$Z��K���b�/�S|�ղ�	��GP�=3�&$^�L&Q��@�k���氌8��V���d8n�u>�g����e�R���-Gc�b�zo�.Z[+����%�{߁V��BPQ���*r�*����ؓ������Q2�Z���]ƨb��1!M�9�[!]��X�N�㱓�@n������B��=��=��e]�U
���;�dbe�Z���g?E,s<G�j!��bt8���0������������A����N<�"1�G-ҝc#���]�]�%r�0�$�{���K�N�����7�/��,��rs�Q/����L�T���Y9�4<k����γ�s/؝�e�cTSg/v�B�H$f�J�="I�D��R���3wh��f�$>��t�ٿ��k-b����%v3�<WǗS������9V���JH�'��9x�`\IH��0��v��-����>�{�൯Z1��b���m��"$�
��v�	 3��t���L��%�C#�&	��E�R��ߤ�lR����*A"�)qK�<�5���lQ�`
u4�Yx7�GB�*c��.�CȆ�9�/�)	Q�)��S���,���SkT�7:+��&��,�q�����0��CԱ�d�.z�����T�ː)o�|��1���@?�*C�_XJ���|,�wt2�l�^F?{R�J^i0�=!���AGsq�}�N������B:]�8j�S3w�"��b� &�f��, d���g�খv�ĹM���ь*z��'��Ǚ��Yj�]t�#�M�����r䚉�b��t6� ���2v����M��R�7!�j��B��ώ�t�qn�G���	<JA��S�l)����C�]a� 1��^���G+ؚ�'/\��ՅF�A�8R���l!��w����l�˻�����9���F�ô�ئ�d��ūn���i�'����=Ko���J2��x+�4N����ߦ}��Ǭ	~�����I��,�&��q���松���e#+?�ڸ=���B�������[f�T�a�^���Ҙ�w$��$P��d��X�7rM�A�٨�)V�
5��H�W�����ǝѸ`���Gͽ�_��Ɠ�0b4��HP�Y�3���-����{ө���[��#gV�>��M1Td��Ɖݔ���)>;�	�����v���4�D�H��">h�����Cӈ�Eg��;j���{��>�[��Nbt�-٭��lCK�Z�y+�H&a��}�o+�=�¬}i�jl@�d~vu8��$ �)��!��p�c4$A��w�<<=~�"�015���[�lr/`!�X��cHsvr�`�q�%,�9���٫xN`��M���}}�^����ce�˃��LQ�{ڧ]�aCa��\	j�B�����2��b�L?B�ˡ0�(�Q��r(y�+ah{���ݪ*�����'�9 m�	�VX�Z�&Jx{�x���ұ�/{"Y/����|�Tkm18��ɶd��%ڢ�z�8�C�D~���UĮ
�_�@TXa�w�Z��4E��8�vU*�
�!��xa��˪�7���	�Z��?C���i#�V��u�9�&�,��.���wެ�K�c�a�ڍ��ze��`��E_b�V�;k��8���7��V���m��I�<K�,��*��CH�I=�%��G�2�P���j�%�u�,Ռ7_��^�P@�cܙ.�>I�ԫn�բΜ��Fi�DC0.r�c-
)�ℐx�7&dV�f�
�s?F�#�����D����B  ��1���%<X!kUu� ��t�=	�����~�
녪-�B��`�[��7�]7�wb�C�E	p4�������w�� Ck�;��L$ܪ"~p�f)�J�i(��J��30N�.!(�"N�F�����ݎ�bS'��3���|5yF����n�_�ح��{OP�iXɍ�^Ƀg���|~���KIT�c3г'����/�
X��,�2n��㭑�}�m�GE�_��3�w��(��vAYk;��P��41;H�Կ �zP�>��*���1����xX���0^���S����8zʅ3�:%��]�[��X�A�\��a���2h�"
 �NBy�\�墥�S��Ím�XrrM4�!xk2��oÅ��0�\�1��ǥ�O�6h;�D�T��lM���ɽn滮�JuM��Ɨ�_�J�r�/+��YGb��rK�8�z�L�U��ə^���3��#��TO�K&��>�<n����M���X�"�KI��;(��Z֭��Po��1��7��!�����X[_�`����XQ�&����TD0I�o�S4�]ܜ�����I���ó\�������[���������-[�c�	P�E�2�8��tǭ@�,;8.fYx��2Ъ��&*�L�Wgn@�
o6��E�6[�؏�CI 5,��%g�ӚC�Z<��sF�!���t�����1��<�1jlj��� TD�Sk��H�cv�<ZI��]g"n��s(ͼ"7���,��_�5�}p�:yUv{�Y��1��,ӔIsļ "����>�ǅS.���ћ�m	��[#0�4�ˮ%`E:��	��K�x-��踲�u�)�a��5K�
���tqYZ�II&O��.[�y���ź�kL�$����uN@�����3�u&�J$BӲsu5����0���1	^F0�mt*�������:z�'���IQF��Y-�H�/%��X9xi���,F�;A��k�<|�}%��k�m�sץ{!�n�g񃹎gj���Ӧq;z���Ɠ���J�3���Q1��(���8�JT�$ZxQ��p��PC�lh^����cNi�Pu�d�@�E�OJ��J��^f�H�d'2^�HTC�;���O�U�ZH�G�)��J{0ό$u���.����L�n�k2��!)f��u��O-�㞌�w51k���Z�Ta��pm��7�����{��_
�t�s-lkE�W.�Pq���d*���!���PX�]a���s)�U��~V���sM	��~g�$�`�y"DJ�b���4�p�#���6�#ޥ��b8��1@l�֏4E�@�#4�u0F���{�=�6��8��t��M�=������'�x�����Q��5��$X�^��/�.���H�@/�Jo�����^� D~��.��n���n<���dd��K���)��k}��=���r�s��R��^� ��u�k�i��u�j�usMB�U���B);���4��h#���}#\�ub֥ه�D��6����G�^Ϗ����,G�m*����:h#y�5��{7�^)��e��7�<��{��Sna��Ϳ~��xUxX��~}̌CC:ݸ��׺�G'�2T-B�P[ٷ����zB;���1ǧ3�3��fBہ���Ӹ�G��yוyY�Py�3�ݠ�91�o,>Y�P���/���M��Q�w��|eN\~��D���{ƣN�!Q I�p�4�9�B(�&z��=+�Vi�`��v=5m�$՘��[���z�r�n� o/��uwxv�(�~�M�:c��4a�c�`'�D��	s^B_k����lcZҜ�����a�qT�3���� �K�irS5��-h|+c�_6<e�v�|ϗ�W� �Q����{�Ϛ>%	��DCϖ���k�:�s-�N�x�eGq)�I7r�\M�.�Լ����l�_��$��_��0�4�
m�:�R5�).�ɻ�ĩ[�m��������{�L���� ���C9��A|3��(o"�IuhT���#��!1���M�$ǲ���j�s�~�P���H��l��TZ[&�4f�|�,�2�2���tE?��	���a�#�h �e=�v���h�:`��Z���i�0jˡSͨ�)�.��=W(��1���ʼ����5�들���J����Z�b��9�v�<
Q`au�?�"�OE{�n{�U�	xT	���;M�*}��Wo�waH��=��=x�=��F2����f��K���Ca�myrPV�r����iMT����c΅x:mB�o���%NEᴟ`&*�8�"6@VS�N1 dmÖ�%Pa���1�>c��E4��m�>��r�x��>��trT�x<� ��n�^d�C!�o�N�a#���b�?����]'}�8��!N�g#]�81��A����9:�̙�K �=i����BƎ��OB�3�Ix_�
�C��Gܿ�K2���y�Q%�B�C�@�f�h����<�{Z!t��;�O#�4�\��i��xI�C9~vj��5^oy��I��J��|��$T`�
�ѹ2'�7)O9ZMD�KM=�:6�����Q�M���g�8����:lD ��Կm�����/�u�/�m�1���wY����+�n��c��r��핑��Sj34M_��8Qp�]Mi�"�P�7iD��v�$Q���'��v�@ ���԰�Y�E]V�F_˹@�hL�����Y��M4�����f��
g�z!�ۅ��?�56}�x�'�\�<�ւ���W�kc?����&��Ꮬ_N�'��qC�wH��W^��3NdΊ��om�=ћ�����X�������hN����ߒ���o,��wo�B��a�:�MA�h��:&�׾S�p?}Xy�7�XtJ�!�z�Y�x�9d��CR���WUaا
��M-XA�0�|e���v�P����l ��l�
�t���x����2�Ԯ�,R`��I.�x�����p�'��_���/exgms��W����A�J�=�/n�^S�_�s�*��^�ځ~�[ \O��?�ߖ�T��/t�]�/'�����@�����	�`�?���M�8���5a7�u�e�ÐaL�
��v����4���5�#�j��Ҳ�3LK` �XY��R
Ix����f�'O'A{=ln+�Lk��������Yj+N�˩�,å��tG���"����5t0��c�P�(�>��T��j���*D�.t#C��u��|�BL(������1!�<y��|G''������p��7g�^T���
2J�����2�x� ߸P.�9�:^ޞ��-��EV�sV��h�)�c��S8B)3��F=9h��]�������IR�ڽ~��q�v�2S�I��V�#Ȉ1��_����pw\{�:e��ߩ���K�ײ&��X���d�Psi����9�E_q�%.֥0MU�E<�m��ˎp�e�%;��Œ��䭰�x�]��sg
;�T��9�o�{#�Fx�,����Z�n&��u �!��-���)Z\���Y|��2�>�^;��M}�x3���U�V���+�p��n)jW��gu�`�"��Ֆg� C���K�!�L��|�ʻ�v�D~b9�8�%�1Mhh~�A-�xĝE�:NF�Jo��0��^N�� V�!�v�ȼ�f��>4V�j��B���m-�!�u|�w���%�0a�h�̡汕�b�D�T훗&��4�*��*�X=0X4S;��$��SF^��u�q��T�����;Y������h;��I ��}b�a����21�X�f?v�7��e�?$Zܜ�K�3�Q\�V<��]yW�#��J�?��@���Ʀ��L��+8hW��ߦ�',ukl[�%u��6�6s�<vM��(/����><��ќ�"(@l:����%8Q*����%��AM�؆�J�S޹>��ڠAy�t+y�w�`�^�Q���!!�	o���ԥ��/Ѥ���=����:0����w�Fؒ�Ȭ��KA\�y���'�P>Q�.ۻ=V�ϒ��|ZD�a��YZ�^�*6�	���͘��n��죍�R���E�%��u��ߴ�8�;s���+�Nd_��7Щ40�^�)��9BM�8�j����"���XO���%�1L7��;����Xv��zҵj�4���m����:Jzv��{\P�������|"�(�o*��>_<
��O��Џ&���8�UX���v����{�U�����w�-�W��bT�6����0KNMByd�ƙ<S�n���N\ڲ��%�^<��&��<%q���ʒ&`8  KŃ�g�;��ɍ��tH�u�(FAvF�`�P0,�NuٲK�	M��Ti2��6Чz�4p4B�S���c��V↚��ۿ��a݋���r=�l���>�*GЪ���������w
�f�MwR��5Y��`��?�	� �	�C�j�h�� �EdZ=���><aϱyk迏���X�R���օ��[�(�{"�:��~�q��`J��&��Ֆj$xmQ����O�6������>�5� �,eJ-��T�G�R�n0U��ʌ_->�R5�� ���l[J�q#8�JTz(֛��V�;�-�2�T����F<ޗ�e�óIO�C���+"�NI��g����ޙٶ�[抷.�o��9�p7J��l̤�����j�ב-�6�����Q����ܳ}�ꏰH�p����*s4b}_���3�:�Ϸ#���֝C*D�m��J��߃�#U����߰�N1�m�ۭ��
�a�R�/g�x�+tQc�{ C�� .��%i B�EK�h�Lig5ﱃ\ĎW�~�Ɛ��X�:H�?���u�FW�6{��-WkL_��NAV�$����1���\�T�,��tt;"N�]����^u ���;e�;x�0�4�/ C�p���;9�騹�N��B��_��a�@��8�����$Ϯѽ�4����Y�ŀ5�+d�6�97rF�!�cZ�2rV�dWK3�O�y����z��V �+�ŝ1�E����3��� ;���g��?h�h4����`�W�d�u�ϣ�E'�X�s�>J��q���ƨE��o=�6v��GB�*8��޶m�7�)��m���h��ƭ3��S&
XZ�Φ)Z���c;�}�=��C3��W�g�h��ގ�[?W8=g6���ZH����딟%�6���L���Ѥ�6�[��1�(��v_�
�Fw4�WV��[��dD�St��p�fX��4oE:e!��l�d衭�7��n���b���DY�te�\K$ĩ�k�%D���HP!�O������x~l����[j$Z%.k���҈�8�G��;��.c���I<�ÿtW�~ʏ�p_|�-��D/����ͥхą�Vτְ#r��ӄp�H����(�F�����H��i2�U�9��6�����������NXї�
+��܉�����OǨ&4͜�C�ަK�>��j��vΪ{�n�C��2Z��,A�c�����M?m�l����0��X�$!d�7�
z%��en٦V'�9T���l��En4���d��"핇!�1��.D6�
���,>����>�%�h.�FE����5D���+�t(��<]�Q��C����f:�\\����BY�8��V�7:65�~����+/̓�z� =�0<����Ɯ��o <S�B�u+�@�����$W��+��U�f�j�ᚉ����g7�<����,'�'>
o��ϔ%��_fF8�L����b�c\�ˮ����Ve.�W"�1�`��3����*�K������	��_��� Py�*>�ueޓj���Q{� _�W��c�����4V�!��Z��e��F�uLX(�����n{�H��<�.����9&Z��������0��\���ې��w��h����cՕ�캳�3��uO$�����)Y���E��N:n���O5
![�We�:���S���� q�]{z�Q{y� :�	P�EU�CR���L��j���9}��6��%2�|�[�7���[8��rY�j��\j3��b��dG���in݆�Εܢ ���~m�OH��` �xI8o.#�O�w��� ��q�L��L��>�����ށz���~��{�o���lnY�a���, Y�u[+wn���x�*x���O�RxR�@�{��Q��A�X��/[��9���5��v\7�OE�Pm�^��z��d�M���OW��u��⽺bǘk0o��S��-�1i�������1�y?�ц�P�Z��i�-��E���Im�X@�Zu��s��� Kcv�͉�Fe�Lp�L�� ��/��p����W^�SY���z@��`��i�#xߊE7�}(���=��}T삔�x���7�ڸ��q����dI�1��}�|�4����U���:�,�+[��hYh��(��"`�@��v���&�M�����8�G�9��K�Å7��!	q�y(��l�4/���Pf�E�)���������\��^t�����H�W�W�f)xG�d�|ϴ�&�1J�"X�:	�������� f�bH$�z�o�@1I�OE$����"����YV�e7���c���Ks� ��*w%��0XīAa�&�{�GX��pު��)���%�ڀg5%�Q��=�͔�ox��s�.�}�M"Xg
�1�����گ����1���È4�pޓB!�G޽���촔���5�E��v"��1���P���o��5���
��0i~x�ZD|OR�?��=G�m_�RjIbF��16���6��~�M~�#&�,	n��� t��b����n��Fźz
,�R(�=�X߼*ܚ�����fU��]3�0�yh��=|WMKA3v�}#�6����Qz�jP�e��	�VEtazQ(Oݍ����	|↎���0��
~�wf
�1���n���2\��������X�X��/&�̬�$/�21�K3�̰�6��Y��Hя(�D[F��Kջ5h�0� �B�j�q�ihT23��N)l��9�G���~"�|lI�;������e�szI�5�^��A�]���>��es�~ɰ�q�f5ea��-��ܣ��ݱ�c�=\��G�Y�8
8��>�C��k_>�O!�@p�X����6wQl��2�??8]WS���l���I���ݹ�2�s���3��dC	���}�p߅EQ$�qY\vk+�5/ob�r �ԩ�hRٶ����K�s�"т��ĹN��)���b�߂fHS��������{̵�+x���%��c��|/u�X"��d��k`T����*)0{��i#]\,Z�j����G8S9q�g�O���R��^��P-9Aܶ�E��6����+.��)�>U둕)�����F�B�=���ݠ
��)_ꆓ4�P��8��aˎ��ڻ2m�ƒ�7\�:W9y4=J�^��T�K��N�4��]_��0!�wBP�;j���F!�M�9F]�
&g���b��*��<��W��8����9�;ѯ;��L��*��씓Ig���7�;/d��|yh���t�w�~ #i���E���9��1<VFX�tP�*�:!�p��I���Ʋ���?9�s��y��2  n�W�`�A$�2�o��*�V�<ר3��?B�����z�	����[����<��72�4���ʂ�ٓT���Kf��@.���.i��������Lt��ripW�ؿtd3c$��v���M�E�*�KY%�ڝ�:6���5��ј��a��f�rq�K��vq����颸�1�J�D���{X�����E���ep��*w��A���D4�u�w���	z��A�
3}�ȵ���xF��3�V��;T���0@����p��|������2��&\�(P������4/�Ҟ�\�����3�T�U�bY[Ƈ���L�������~H����%B�̻�C��ќݽ�8��=���P�e3c@yׇ�����.ٝ�Krmy,T��2/e�7��������\ܐ�fQ� ��?���98I�S�x�>I�&���)����ؐ&WMR����Ӿ�.�c�W@���)�Ա^�	q��s����{�UP��8��Y��-���j�x)�@�f�?�5P?�b��/?K���F��������g�P�������=��UB�ش�W�ت���%�N�Փ�ss��r���t�uU��2	�XWZD"xn�[i���Q8��#�06��E�I�D�_C!�O�K��Nz~����\������˪�:'��5m��x�#���.qQJ����+<��_[����f�^)9%��-9w���R�m�\�-�;�ZBS���s��X�����vD��a�2]��q��C�ÀC�2�K�ޠ� j%�'��%G�y�s"�}XQ�B�UL)���W���n�)��4��e$�"z�sY�J�-�
�Ic��ĎE��f�>��50<\b0+ͻ77��Tp��0���^0ર<�P ]=����r��<Sa�L������w!�
V��
��CW�����y`���r&�Z�?ӷ����Wb�q3� /!wA��dd��Sр'��K��].��d�>�S'��m�h�� K�MA��7ŀKb㚋H���:*+�,:N���IFD!-�|U�m8+��X$�F��&2*�B����C]*EK
@����z�-�&�>�W>ך�,N�i���_ ���b�C�2���m�����2�+a�s�����Y6���J�l3�]˰��÷ X��ɶ�`�Sr�Z�g�r�r�"�O)wW��h
�4�b�D�������B0�����cQ\��3`p�����؉.�@�Z:.�,bs������|yu�~�/-�l�\b��!h*�O|��`�(�B��$�����J���b�����\��@ǅ����մ�2�݊�ۯA�0�xKB�b��#HIP��֮�g�=���|��e�>
���]���=���8VDm�D��	�d�	���E��f��p���)������S��E����4����h�����i2q�7O�m�,&�\"3<�]e|D�Y�2�t %�=�Cx�n�<C�y*�������=L����Da�a�iD_���HjkM7�g���$���{8�Al��a��|�a*Qv��B	���� z��a�`*��=lY���t�5EC�?�`HӺݩ9.�'�L\��C�ᱏ;Ȑ_�zG�G���B��K�Y_��_�I�ș���w��Љ5�Ig�αN�-����j�y	2�w�z��
�ŋjn����g�4����<	K��Z�.�͊TC�"L�{��������싣����u+E�>���=�R �[-?�g���9J_�����F��ߚ�	s�P܍�{���p0j���a	���bW��)��\�G�\�K�9t:$����@�L	�(��b���!����}�:"C��ѬyH�XO���N�\VQ�2p�f�cȱ����ҋ ���φHJ�U��`�Vg��!�rX�����K�k�h`+Yd�3`��񔈒��dȸ�����}�����z��J���DZ{{~����)�G5�E�֠2��?�����/lZ�O�g�i�ݔn�rw�e��>!�2����vg����� s]�j��u�����t܌��B�ns�C5�5C6�E��P�G;�O(`C0X�1�N��0��3ߒ���e0F�(I�Go���kԸ�����˓}�n!,݋������� ��9���f�z�������.^�5�t`��z��>��ТT���/�.C����Q���0G�3�)��ᗊ_�y����{��/�� ��+��6Q>�ʟ\L'��(�XھC,��M�\�:߃�����l	@1�F�'���K������˵�r��-|?C����(�|Z�x���2_�,0��7CK����,7%�b:g�f�[>F��\�F#�ڗ��J�'�y<VХm��5<��z�w�o�횵$IY�DCi�At�;F}���@p�=s��$q��M*���*wϐ<��#����+�e��7h�dӽ�|$Q_4�0Ұ���5@�P���Vj����es�xA��ڸq]I$y~I���`�T���	}��Z����o4���us3�Ӯ���^�{�xQ�4u��Fr�I������	�����G{4)����h���lp"O5���-�|o[c�,�b�{d��.������s9�eo�L���ӗ��V�25g^��,�N߈�p���(hT& ��66���덍L}c����N;>�5]b�Ձ��@>o��cj)�hL2�c���s<e�6y'1�X�ǫE
�B�[�{�{������(ja� vk��rХ�R��97+~>AO&�lyO���A�����U�Ls�W���9-�pKW ���@:��k��s�m���uB�ϵ��U����A�z4��J>�u�I��<[S��,~��Iz9��`���AR�Q�F�m���}���o��E �?EaG�`��u��������M3���Z{��N��6A��h��-�_���!�4���e@�������8���4��D��xU*.Ɨ����B����E���=B\9F@
w�[�el��x���R�XiA�4K�����M�螁��,(�ɔV��v�tg�>�H�D�N����DH�'~��MM���g��<ҝ��_51�Բ��� ��̀@�˝ڹ�RC��݂73d���ȧ �l��0ڄˊ�u��7�0OB� Z��3i����]T�%�槩�SB����Oa���ܸ�� y��U��cԺ��˓Q�	`�F��\������*c*�=m�	X�Q���:���3��p7a�xӁY�3uL�tV��fu���$88�BW���+�[��X��Opefb��6��������n7�@0�(C����O��J�	}�KNz4�3���! �����^y�ڲſp��l���o$h.��s����م}���cō����P�NC�k�x�h%��OH���řX�z��n�Ǘq�����V.�$Y��=U�T���TѼ����`PFi�A�+i�9���o�AWb�Իx��-�`�T/�=üI,+�8���V��8��Y�k��x=��}��[���8aq��Y�D�b*��3�6U����i��6U�x��x0��X^#<�v!Y,����)Z��D��ok�N���Y��0�Ǘ(���!��*X�Zc�l�tf�9`�l�3�M��Lo{ �`���)� K�x2kI��O�E��[(���)��-����~���bW�zRT�$yx�b�}m�\����0a��3j\�I�k��!g�D��R;�����2�ڱI���=�j���N��j��)��
�L��l(��!�� �۸Z���u>|�㯡���
�����**�Fo�� k��cr@�m�醗����=��"d��F�pJ�]�Swp0���h���wV^�w�C���,߸}囝'FK�����Gn�=�L\��[<�	�8y��?;�޺�6UL��TWR�}<M��#`�eIq�WU�|�_��q@�"���N��޻f�z����d7���܋�Ru��>��X�C�/�֣����d���q�7���ۯ=f�%�3��!aa�{Sg���b/���u��
es����Z��67�$%(�,a�3��#|���.���%1�'��gL�.;Q�v|�9�+�������>��w'��N.Yln{K�Q /�R0V�V�8����7C���űы�މ<�t�UQ]��Xd���e�RW�0u���z��z����Z�d0���.�GZ0>g�ģ��+o�(���������ډBz���3$��v-������ߦ[5bw!�2�����u��o��+=/�M�~r7��+�5�~j��8�T��@�3�F	p��B���&���\0c�m���@�>WzL�V|�y��S�K�
H%4���yL��$F�{�᥀@��}�%S(@� p�M7٩��,�`�~�;ǂ�@P�����'�B¦�ЙQM�W2��aE��pK'���E=��$��3=��6��W��ыB���q��?Θ�~��/����\��!������-/��%ҧkD��ۛ���̑����:N\��~t·�΁	XR�'�����9}#J���� ��a-������+��,B����|kF���ʡ+هU��a|�.�-�W�*��B��_���΀���̥uEDΗ8�=���������6ƙ���D ��:��T���!�ѤmnYS�s�b�2Q���Q�q�/�'n@�^�b�]0Z���4�-�\��0^'X�Lw�1�6���$%,?�,R��;�AZCa��&�-U�샕��$d*K�����'S�	���;7
M����֖��7��"�ת�}��Ƀ��ʙ��1vT����b�k�z�G'�(��F{+���#>y�����i�GXV)�)W�D�1�����;q]�M�g��D��qЏP7w�T���%L�k�e��,���*��7��KW�\�U�W[j���O��D���b�^��K%f)����3����!�Kd�;nC�x���o}�܎�ڟ�OУt�Tv�س\�:�|�+TZa��6p����4)�&o~����81����������ɕ'����g��ؾs�!������p��qB��J��3+(I��� ��{2���_a���T�U��f �1"~~����'�{ו�����qc㐉X:���Η"��8�b�A/��S#\tƨ�Ry��(!���x竑aF1�\FC+�a��aymh��9�r���Nū��\��Az��&��m`�O��@��d���Fa�ßd�C��U��F �c2�s�U�1��9�w�{H������T�R�Nn2.Q�]%F3w�Cx���4E�AZ�S\��t�G�9��Y����q�fRa)"��<��2��r)lؤ�a,�G	>խF�i]d�"ao�!~��pԑ�g����{ڨ怒�*WX����8����dm�|��\�:���_�'����@�'M���HHn�1�4�'i����va�P��Ų�������f!���r]R�B��������.E�����8��ש�H�mc���O-�P=��Kg���:��6 TQ>o��c����ֳ/��$X�m�jS$}���E����X�Hg�' ����f�n��գ�+y�>�^�p�B%]Y�|�۬^��Ǎ8�\~�h��I��B�eر��u[o����}��D�{Qz�����\���,��O,�+��T�����@�o�����wF�X6gv�mhS�93��"��%r�=8bǖ�K`܇,�G��ɺG8�1Զ)[��Y��䴑Y��qZ�#��2 X}~�7���&�rh��X��|ą�˞�?|�_�	�} �]T���yD�t�Š�6�&�L?�� %�I�f<�����G¶ӗtg�qAX��\ӹlf��HQ�3�e�$��,��.L:G5*��u��%��dy���Z��0Wj��_��.�����u})���Į҃��ә�dc�ie���c����aZ1 3}��ӄ�J)6��n��@��_[w��6��Yu�p�x�g��! �$pǺx�s�	`F%x�RrH�Wu�(�۶}�.\f%���B��_�oPY>��8�ߕ?�GG���r�i��G���#��z�J�E�2�Y����ݕA��KY:�gg�0�S�#K%�*�l�-)������>��
�P9{�{�JS�����XE.�Xlv��\v�^��~�N������M~��G6D���EDٛLAs��srf#.�)̟eb�~��U/-?X�0��<1v4�$(y}�CH��^��Q��6�^jT~�3�(<��9������I��>��[f�����Njm��DUXi�@ԋ^2�?�o��y1��B\��T�d�Gh��b��A�_���X��VUBN�6F����Z����5�\�dʃ�񒄏�~������!�'@��M�n��d�����Qsj�10Y-ޓo��VQ�����<��W�R,�O��a�5���!�y�Z��<�v�&�0��«�9��S@���^F����c1�BA�2w6���[iO�;'_�B�(j-�z�����0>��[�e�#H�����;i�	(e�se��ץ�ߔ���h�?���!�*����F�Bzҵbs�?eNr�9�Vݴ�WJ������/fe7������R�P@k ��T8;��շd/v�զT޿�[�.�?_n~�&`Y�QK�0�i�4O�4��9o4�j��ub6/yw����M�X�']�\���#���حAI�o���8�n�i�K Ѥ�]mK�i�d=��K{�2u�qB����Hr�PQ�8�������I���B�j]�[�(�b�ۼ�C��A]d�!�X�>�n&3%�y�~z��q��D`{4!..�m���qi�Y�d�����R{�?����}܈�+�[f�xW�J��|��J��#����ý.��Ƞ�e&�����#��q8���Q�z �Hf�NCM�!�,L7���R>�!�Z#<�IT��}���n��ъ�s�������ŭ���٢��\��X�k).��ͬXm�^����=gI3ө��:���l�<2s`U�� x�[��k<^�
e�WA�S�s�\߶���)�u���<iN���םp&o�v�%@Y��G�͢�A:�ד_�wC��7�&���@�҄�S��B\:_{	Ci9��H�@W�]��|�r�4��{�\n$P���K0;Q9�nNM[^�Ҥ?K�|�5-��x��[l��� �ν����q���7���VGnC� �m�j����o������&p3�Kp���7�.�^9:�Í���S�)��U+ᭈMپ�7�&��nE�6}EMTS,tcϫy2=�b�E�g�%,��Mv)D�`�i�����*���S����e�gh}��`S.���"P����q� a\�^3�s{�?܅�1x���F�;��tJ&*��?��;gU�0���:�2N��d��Ue�%�eV�O��o�����O-О�o��#�X�>��e��6��E8�?e����CZ�UB'��>��O(��2�6"��\�P��!���?i8�ꥻ�	h^�?b�3Ft�f������vp���8���.i�Yr�҅d	�꥚q[��8���n̣K��Y����hx�Ԭ���7Ƃ�t�ճ�_�*~���<���:�S"��B�b䓩�v
{��_c�޷�֪�Vz�&�6����/�����N��##҆�xx~��J�z����[ݘ��܌��ۮ9ڱ ۑP%�kL�����|����e dfghM�9!��3���&���M?�O>n)�7��P�V��� �Mh�l���ܬ�:@6���0%p�t��]dH펋��s%�"�n?�i2J��p?�I�*ܷ`=���l���^�lz]�e���z��l�>��?:+g�7ݱ������'�U}Z�Ov�������1(�g�o"x��^�HSP��`�+�c�EI�4m�}&P����`�۴���Sa�<WR�������d���塕����'O�'�rƽo:]0�!^�ms��B<Pt0�$�QӪ|���,y_0���5ܕ�{K�d���UQܤ��X*k�5P��l�N��k}a�����߬X����:�?JTSm�P��N���yH�j���p&��kWx9��Q�GqDc��2B]�l/ᴦ[��&���K9V��df$�t���K~��W�=��0���|�t'�ӱ.�ĺ��*�I���^��.(��r�4)�}��G|�64}}����~JsI���W�Ƅ��I�X�����^	����$�#o�����s	���
� (���M�;�I�cC�F������k�F5���X��G!e�ۙ����d{���	���EȜB��*��� �XQ76�WB�eG�f�8��m5d4�[��s��zX0i�y��g6��[o;i��/zaW�;ʵ�^k'��ɅM���shN���Hv��%L��A�Ⱥ�<��G� ф�qL������)O�#9K̀n���;Ƣ�w�d�ہ�5	�?���J���֥:4�2���
���"�2f�B75	���u���^܌H�V�6�l�0�\P'������8�	��)��m����,�k�Yˀ3L.��9�7�ɐ�s����ڵ��f@�(.�t��Dp�M���8�� U�ʈ���2?j��Q�1�D�aA����9�����F`���]�4�侫�X��,�W1Ϲ,�]�f���O�`껪Qݔ
�J��lM�r�{��b?>Dë�d1w�̀�XCf���R�`�.���4lkn�ws��Y�-B�nEH�e�����5�E�0t�^����:i�߹���S'e&�L����~��.���ul�Gn��c�묹Ϧ��z�)���_D݁��;m�F�:KN��Z��w\E�M C���@�Mѭ��յ� s�rz���V� I���wn�e=�TT\�D��C`�͠n����
\c�~�S�eu7Y�Ua?���>�dBI�6W��?�\>���Y�$m�d��✺b���Q�����#:ͨ@�\��O�}
|kz�����ۥH�h���F �z#,k�t�qr;�)w�4G;���@s<~y�� �o��E2v4p�V�}\#J0f��`�
3�pl�K-U�%f��/¡PC��$Dx�:���hH�SG�"��R1$��ey���{M�����j�A�T�c�6��	[Sjܝ�0�@�Z3[&���#�G$�s���� �_�/�Y�2zz��R|~�ɜ�G%���|ݦ��뀹#,�3[��x�6�`LD"�'�o��l�-�q��Hĉ�0th�v�G# 6v������s�R�c���]Rz�j�-~�;�lAY�T	c�J<P��,)�%57$�y$s�mUg�(�෗�w�g������x8�^+s�4ب��KO�Z�=��\D�����?.��la��,e��q����p:h�.'폓l�������H�e`)S��Eh�rp����C\:iI��XG�������Nxb�M��ß�@��W�ܮJbJ,�d���B�y����'V���6���yfBBn��5�ҭ(e���F��ѷ7�w�f��L�.�M�{����ħ� ��}|�~ cs��(��p��
2G"�_��lG�#��F"r���}a���E<�
�MD�KD!{��՛��N#;9wp�n{o�6�I��Qx���~MFA�9��K�о�ec~*�^tu��
���/�-l��")*�������t��HÊm8Đ�H����i]�'���	�T��L����Lk	��3q�xfs�V��l jp�V� d�eu���KK��$,�:N�f��Y$����딹��çB�a�_u��z��cEbwx$�i9�	���GvO�(���ퟭ�����3�?UuvPX��K)N�3���ɀK�'�Ń���Oʧ�׆YN���/�"Z��dm.��=-�D�s6����\���:��p����(?�̧|����2'4�y���I�]''����'�rDG�Z�*Ƒ8h�q���NQp2�c��I�P��rY�]�F�/ i���"�{��er}k�7:�G�В��n)���_����θlF�~R�j�7}~����{b9��<@�(U���#g(�/[o�b!�T&`)Y����	�f$�1�����
h��*d��y�� ���p�9ĭ�N���|�wӁ���[���vz���ٷ+Kf��5�No?�9�F*2����<�`�C����9o$�(�rV�?�U3#J��L%7� F��h�叜��	pR���ކ�H�?-�y��V�}���B��V�v3{8�5�Wz��Z����F����;`r��,�e�>4199�1���![�fU���<=���Et^6t��"�#�,aҖ�׸c��[*�0��g�B��!�H�ُW=;'�ɦ~�Ӊt�����am��@'�58�ۿ�_�D�܂|�SS3 1�d �y��=Je��w,����7����d��g�j�tX�T<�U�¸X�"&L([����rD$�cM��l��j�u+����ل�Ӿ��iX흫�M�_o(}�C_���Tp2�Ote*�c���A"�Lr�N�� q���w�X�Wr�=6ֻY���W��i: xOr�&ƫ���F��%����m_sm�@Y`��PǾ�7�+���/R�[$�%!�>y|�T?�[M��ȵ�`7C2��nE��F�qb	���9=f�k5C��-�*�M.������E��6�nC�n��a)��W���w�{唍�];ou�M�"wMA�H?r�x��0V�x=m;���q�W�߷�yʫ+=��t2���tl���}|e�*���)g�[?�Sˊ��RC�V�����Oye����T���IUz��Ip?��
^'��	�>�T�����4�T푌�g����1�	'�Ed:��0q�X����a��)����5�����9�?�s����Q��s��d�d�p��<��3���D)��א?SQ���_�b�WV�x�TQ�O*��Z�`��](3����ݥPE�'��׌UM��q󱐧%ӟo��̐�˗*�K�Hg�(e��>q���(�G��R�֛�D���,m�F:��_s�Z  n�8m���_�����4+e-���U�Eyi�;��c�w3Y擊�㡈ƍ�x��V��N�˙��ˎJtE	��n��%���
_�o@��R�Aڑ�Y�������G5t���_hce���^�f ��t$w >~�#�������1w@?haL��@ܣ�57�x3������V5OsSn~C��h�%�D����Sh�2�#'ЂJ�S�������`����_֝{��'?�r@��k5�n���\�?�̎0�h2��s�oT��6�T�B��zb����y!X���f�S>�-���^y#��-؍��n�T'��2pU�&�<����ȋc��Q�\C��FZ�ޞ���\w~��kx��������a�h�R劷�kv}9М��P�F)���̮xjb�.�]�:�J���e{kTi:���Ό!���_T� h˫�xM��0;��AAz(W�;Z2�P�c$����y�-�����Ǚ�!�LTW�``7t������Bɾ	�kiW�T�҈�E`J9X�g���_}�5F���G8�6kg+��z��hw�p��R`�,�>��I|��~G�W�	�o3�!N6*"eO��>SCqײE=�<}!�����И_:<t8
	;tqW����Ʋ����
 �Ԑ�͚��w�T]��if����b�O�]R]��x��'�����^c^:y��?P�>@�KC!ړ�ƾq��i�%�5L��h�-�8�,t����b"<J5h��GS���LSS��H!�w��ȇ\`��-�o���nE�9��7�%9�@��R��1��bmM�8�k��f�%�˶m*�L5�%C"ޥܰ�J�YrY
��1�HUE�o�1G�}����^��zRB3� �b���;qȇ�eَ z��v��\�X�%	��t�ҡ�#�K_�y�9i��P��Y�s�h��M]g���O�eςO˟�#���k�a���&轨
!IO	���2l�!׺½Ѳ���9�g��������\O��S�H�d���:��ق?Ǵ$0� f��CK�8-[�9S���}�{��_�}���D�iw`�bc�l�*����i�{�m�Rp���us��9�mV�����dg�v���	��9sª󵩃H����S��A�����;���%�^/����j��tݘ�-�����a.t��Y^�,��,�����a�+K�u�~δ�d��s,�C_A�.���6)Aa�J�kĈG��f��CN?'��D���,��5��V��1V�}�$eG:C���Ȇ���2
���#`�-:��[ ��3+���jn�	H(�w���ӯG��|}[�{��v��a�-S�ŁY�u�,ԍ��0v�Q�;�����%]�1�����8��WG�et�$n����~�?Pi�wAq���`ɣ�����^U��*F�>�iJ>�U�(�5�hBx�lV���:�ȩ�f$N��y��N���H���5M%o�a�+�HDT�l��0
�{oZц�9��E�I��6P�*6>���B@�~�Fp^�s��O.E|}�_Jq��t+������D$��v��B�V1_�Yy�,Q"�>\��w�5/�b�=&���o�(��X2���c�6������YL?p��G���ci�*Avx�-ڋ<%3Qj7��xj�ָ�CJ�9N1L學����-�$ޜ�أ��n� �;��q��m�$U? j��CS�GصLЇ��������/� u��6��p6XZ��de�~B�F�B2S��_�	��]g\�9����*;��e��>\�����5�z�t�D�'{� ��J�mq�[���G�mo��sF�a��י��d*?,�S6V}�G||t,�&��<pX����[�)�	�_��W�j��%4���Q�@D>�a�|vH�&%ʉ>��D�(�0�,��]��}64L�(K��S��er��6��z��SW�O�	�!Ai��@E�z57u���/>l���nù����\�o�͝۩�E趰Ͳg~'I�C��]�a\@9��KG�ڸ
��[�!��J<%����Ը�V܎k�yK�݄��oW M�9��Ӿ�6��:ЧzJX�M�z����@v#�,f�v�o�£�F�ֽ�N,f0���N��;���j]���1ϣ0�U�r�4�z��f]ޙ6�qkaZuy�q��_��9�ɷb�b�����9�Z�:W��L��Hk�f�Z����n�t�1G��\X�0����$���=x��VѨ�Z�;|i�X��Ӫ<�,��Y}\�R�:�cRL�G"Cg^Vt��93�}�3�yqL���|��t��_�	r�@��n%�ϻH���~�-���6�"d��( �=�lG��d#1-������@Jڐ�
Oz;��M��o�ma�V�CqfCCG��e�;I��s��)��������(��+��@Uh
У�*��(�D����ߜ͗���f@����V&����U��%�1[������.sY�/\�'�M�X�t�A�+$:r,oĲ3�@�ȍ'�>8��~�݅;��,�f�N��<�Kis����)@�Ǎ����� Z����xra�� !��h[�xg�p}J-bSn\~rc�Jj��V#���rL�����v�'�4��[앍��f��ʷ^?<L)n�&���M��7��S���{'Z��V��[��b|�)<��e��f�چ1!�XG@O�8�T�꿄��h�qz�qSvTq�"���%��˽���%��t�m�р��Z�|��k%����>�m#�$��U��P��e- ���Ȍ^Y3�G����E���Ą�_�!I����,�`ϓ|��b��GE'�N��-d~�D-x�q��&�Ɠ##�������H	!w��k�G#A�K,�;gǩ	q��5�8UPC�0#|?F�p���E��WRU�`ƷfT�dYHݮa���3"V�1_��KТ%��y���^>ǡ��0�̓Pj�=����h���'V�c��F��.OY�!s�LC/v?E�w�뭙;�Hص��:��:G �DV�v��4�+����5F�n�����?q��i�?�!}�e�V� ��G7�����l�&�-ۆ�L+�0���_yX�G�&qҌ���[��&������Fas�T���CK��#�O��C�e3���߹���q����R�x��N�piM�f�أ#2���?#��ŷZ�̀j�8}��/�7��`5�ng�(\�u!=q�k�%�ˊ��ȿ�,ZY~30���������*H/��ӛz���g fzd��Aj�R�D��N���Io��z}lu ���s�0[{Z[Z<�=�7�|�1��mS��Z;5J,E��^Y�q?����PIU��P��5�W<�v+��Ҽ�(oǉ2�my�+=�(@�r����h���Е;����3���_m�
�{��*���b���*�y	/�VXˣ��J��Ʋ��H�h�G�CW��P���?���qG�#�@����>���0�;m�Lm��������n�*���󬟪��2�?-�J�z&PKM�����K�<�"������-#�70�`��W0L�g��wyJ��0&CH%c�.ɋ8("�I����	�E��fJ���Jg���A0�>��Ҝ�D\���c��н��K���>�)�Ӿ���ITF|�XD��r�)J��O���/�K�{Mi�41��5q����)翳�K_�|�p�z c��տɵk7��l�{F��)�40�V���9�&�]j<`�(�I��>wp�NC�rr���G<�~����U���ٺ�h�$jbnUZO�T^�)����wd���gPf>?����nrк����a6H�z�
')�fץט�ED���Uy���t�zl4��!	�_-aV�N�y
�1'HF���>�K��UJ���a%X����Ң}d|Ϗx��s��Qϋ�LU$]���>��ݑ���ӌ*^���5q��6�-����D	�ޑ An�����/Ѹ5�B����E
SorA��9�I'9�T����YG�rڰp:����K�֚Hs�r���B��N�TM,J_��Ӛ�13�(���Cd1�(�:��p�;$h�p�;�b�9&f�BJ��z�<e��Sl�Wm]C�#�K�C3s��HĄ��y��IG̱|�~
w�����C}&V�A\U]�_��ـ5�������zP�d�k��z�����Ȝ�qO0ox��R��4�e&a��7�M�V��� r�[X�Y���Pq�9O���p���|J����$\U6-�{(^��շ5���`���	�߶�2�@��S�I1CB��ғ�8<N�Ibo+��,�]Sd��lfB�(8�2��;P�2X?�*f���LU���r�2�y$���l�v��o��Z�	�y�xt8��Ȇ��g�CZ�!�ؿ/�zL���@�'�q'�������ᵖH�H#QS�y#l�@e���;���D�%I\\Q���A��&��I�v��O4D&O;�%raϰ�%#}�c>�� ���Z�<!��7��"��-g�6����g�� e���vz��5����b���.����4���thɑ���D	�N�Z[�Tsm��ڲ&I��� �5��$SM���F*�R�~�������~��a[4L�b�����Ƭ?��W��aa��!�%Б�F~ˉEm��^KvQ�JK��
M�E;4�&)WH7�ٮ�w[���/K�}�:ޚ�.���P�B�i~3O�~V��0�<Ao�ot0�׏?/vT�:�}!̮��J^�py6���_���]*J�ϻ���r��Vݪ�W�rJͽC�=�u��ٴ㣂�	5^Eu�$RUKem��PӃ��n/d���И���.�D�9r��H��
�vB_</����є�ڌ�"�)_{4�H�爪�I�v5}���ؕ ��r�]�Xu��N�(5�8���Ԑ��}�bx�Ų	a�O�a�?��qHR�^��<����Es�y��t�>#��� Ǘ9b�k�� 6��M�M�7s�Q�b�G�"q�^$v/!,	/Y��H�������������[�u\e0���ly���M=K��R�+�5�8JE�-D-�l�$x�-���m�]�Ј�<s2ȸ�`S#��ٝ����$�Uin_ؽ�r���	U*ʦ���oT�C3n�K�ב!P��GZH���0̦�4�'�n�
Զ1)��ı�!��j2�%�C<�w�e��뮛��a~�>��#��*�{m2��:
���x���'�Z�[�=VSE��F�	�T@x��������9,1������g�;nbs�F@��JY�����~:�����4�j��m�kᙙ�����������jAG��=��u�;��P�4�4B��ۈ;0`���~�EO<����~75�7�1�D��mg[�0���s 0zkv/��s_n�yu��|���JŰ�i��}��h8zv�\=�%�b���
�����{��p����@��g�U$�Ϋ5���0��^���oT���ZxK�>�X��G���k������:&��tbHǸ+h.]���˟��A��~����hy�a�*��I���N�w*���@k�^K@�+1�g�I��ZV�Z��L�� 5�UxG�QU���[�h���c耯�J�o؜lX���/S��C�ۊ�J�Hv�چz���~zk\$��������	l�?�T}}-�9%*���_�*��p�@��`m��<��mAz��x����W˴�U�7��עԈ2��e�M�	ۤw�L�yg������������:�-�2�+�c��B��i��GD!4���\���<,�i�}[t�vW��$j#5�#�:kN޲��K���ks���4��GgyiP;y:���ƿJ�D�m��D� D���g�.%��>��F�o�KB���L9�~?���,��@d�@?��h=��7���J.}P>��b���A!7dL��`�Ң$�$H� �Z ,3��bo���*�\g��F�e����GI�l�%����d�U��+{P]�ӣ~�΅�"p��[|� ��E$U;�NY,�߁�lB�n�5z@��|?������%���r�Xp!��okP"R��b~1�P?�n�<�4����3�Z���p@�V&�,���d�%k^KC�g��H=u��G����E�m-=9�M�ިT-sP&�=��e����/�`�V�2]����DP�@i�I��^	���E=�3��$8Ēj���C���e7� ��c��=�[�)?�;u�*
�F�s���[_:�u�0p��x�a󢆴����tQ;�� �_G�8qft{Av�-w�U95 ;�yPI�$��%}�(�(��NfyJT{�
�0�x����W�<9h��x�n�#خpU� ���t��_5�_��ʶ'f�̇������=:>��A[�S2�n$��*k��nLK>�o�T�B_�G\Γ��mg�A���5��g~Rw��_1�f��P}������ʫi�f2g[���M�8���g������rL�o�E#R%4T�?�[&8&m�=�S���Ԕ8�r�X�"x.�ܨE}��`���g��ah"��̼�_��>1�d �if�`
�PҒ��1�q\��@u�����ewc����������� {b�O�0�P|�Ff �rO#{�懓{��h�~x'��V�6��C�G��A���9(\���-�{o�Q�A�P��˸�=�~��ي�6��G�~��糹^�l%'�W���7��s�}l}�$=���1�lO[��ۖ �	a+�N[�>�z�'�>�)8s{����7�qYA Q�K:8��f�8��O\�����Q�r(�2أ7!� X�1W+6��0�.A,���گGZ�奎��p���s
��O��X�����`��������M�ZX��?�!憟J�"w����H�f2��K�I��t��%�1�$�TuZ����ӑ���J���g��IsS�a���~,=n��JR�H��2�r{���W����k8�Ǿ�F��l�_ >
�M�����\A��@��ռ.N|����D3M%���-�'5T��cqg�h�\�FY�uL��J���tl��L/� �W��Q�sª@��������~/`[�١����x �d�m�+Qs�Gg�u�o����1X�[kS[$5����c�ĳ�p����=% �lB����Q/�։�
��L-���%~���~:�_\T��Y���#��g����Ɉ���d�JC���&�,A�s���]E��<�����|�7:��"*ma,��Fw�-Y�:WޖG�t��z<[~ֳ����(Br�tLEi����l_w�K9:a4������p	$is����S}[�݃{DW{��X�g�j�E��-bCg/��"��i��p��(�܌`�`�.̬Yߚ��n5+�B��˟���6ikp�g��3r��߬��t$ڀ	P+��*ݽݼ��T�	r,�3^�u�X뛕1�2�="3ȥR�%�l��<Ҋ����"-�qd�y�+�s4OiD�Z9�#�)��w�4��ńf,H��� ��pl�
	pO���C6�l����|�-N"�[��1T��4a��k�p��qxktBq�F˩��^-�/.T �F}����8ґ!�<�����|f��9��x$�8_�i�	�kc�F�&���d�q���M	�sr�Y�y�?�\�����)�%q��'�wd(�A�>;�DS��i�]� P�v(�mn��	�D�
���e]���o���(~|V>�V��$o�(�s�l�zw�e�_=��f�Q4�����a�\_�,�UY08�AX��g:8��CS����QP���I��r�O�f��y`.�S|/XL�\b `���>u�BM�A�)�n�H/�A�.���(XcGc�����N�����a엃0�I�Φ�&�	{�(0��8���,���8PN]t���x��].:�ǳll�����6dm�L�B3g~ȫ	���A��>:���i�68GP�bT����a-v�<u݂�Q��#xYV~�������`"(dB4L�2	�Y�����s��0�ť��2KdK�su�Z/��#�Q�k�C{�����U�0��bd�w����`&�ǵ�fK�w�jӸERI�)$��{��:�[e���=U~gB��DLaG���>�g����y�Tu�堛����ț���qj�b銮A���><ӊ��v%K�PA�xPB�s�bg���ݸ���f�n�+�a3n'iQ�/��F��^�<���p�� ���bB����&u\�P]%)*�V�k� ������䧴����r6�4���<�@%�;d��z�O"�S���?4w����4�qణA�@�)�n��tۢ��AO`1f�v]����rA��y�u�%{���fP�v%)�g[�zP�B�z[<id�JCwy_,��W-/ވ� �X��K��4tm�}s���� ��:~�<��yf`)+H��O�dm�H��n�`%?I�bU�d��I�-�gj�O�{���3�]�VϺ�[�WX��х�0����R/*%���"��DaE��!������	��Q�� �y)�����y�S6Z�H���*R=����b�>!�v7t���CēkwO��A�SD2�����л�t��q�_���J�h% g>�Fy^l��vQU>�˸�E-�3½�.w��D@�ѾMB�s��"5ژ����dr��k��J�b�u����9���[AM����s�7.��x9w5��8cF�4���4FG��i�
�TL
X1nu�Rw���nA�ȅ2��%]z9^�
Wu��j��!���d��$US)�J���C"���5�V��~x6��i�%�j(t��������Z��yX�'�T�|v�Up��7��� �ЖyK7?��Q�ֲ�.I�C'�!_�w�>ҙ���1Sm�Y�c[��������Pl�O��2��d�Qw�?�G���P�d`��0�w���"k[�&�������Px�ZB1�,\@:�
�]�Y6R?b?J�{�kY�z4�筒�,VzM��Huz�Dț����6U�U��5���n�)K���w�"�_�ns\�)���i2G��#��U�i��$#ￗu�֗tc4�� �)\�Nkr֑�����r"�r® �"��qA>n!'W���Z<;?���⒔�o`G��x��v�Kxvu�+�� �[��|,e���S�l�h0�	�Yf}v��|��ѳ�����
 �Q��qLLr����� ���	ZV�JVK��u���!_\��C_NT6�,�)���p�%6*9s+>	� =��$*���� �R2�Ō��F��I�-�ә�I�G��w�].��}�&����6غ��-����ݦ�	����Z]���y��6���θT���M�v�B����V����
!��繆�d��v�/�t?NsfQ�� �^�Q	'"s�'�@5���������m�J�cMXT�2�c�P������R��r�����Ls/�[Ґ�ׁ�_ݲ2j;�E��Ü�Ц��Md5���k�1��q�2�v����r߃������na�`������x�/;P�yQ���W�d4u|=	l%&%�Dײ��;��D\[B1� j�����d�1u�5����$[�S� B7�����r@�(��/�O�h����PHl2�՛�E���ڢ��>�ѾT9��;&��E��`T����oU�
x�P���YaΈ^�P�͒$�?�h�'�n�qn�J����$����M*�f4��*R�#�%��������Cx���8=G������}��М2�mƑ3I���!9��?2d~9���h��2a��>���K�󇎃U@#���(�~pu2U{�����u��$�p}���.7�2@�uHrǓ2�S���T�Ä�7�Q��ť���1\/��p*?@�4�����NT8P�<�n�/�lDi*�'��^,Ɍ?��˄lۇ�"^���	����TD������N��N��}ijZ�Q��gb�����+�X����3�^�Тj��zt%��V�P%FP>�z1�5�'<��:��P @=�C� ��s��c u�Cz����Z��*ş��޶T�e��s��џ.��G�b�������A+~v�e��!�&#&���4C�'O��bI��"x������T��~*�,l�d�����i#೸��l�c"�83��A�!�Z��υ2������V�6,��$"�mTQ/Y��Eѡ�ʅS+r�%�07M�����F���/8,/#';&r)���5��v����U1�!
ʰlH ��'�z�滟U��^�c�&��{��n�	Mnߺ7�/)��{)��ψ��!���҃�?U�Ӷ?��/���n�d������1g�XS�/��4�kμP�'�"��L����k���0އ'��P�fO?�A������������V��A�����OR�zN�ֿ�F���l������A�G� 6x�Ǝ�=P^��5�a|���N�*��l{ڌ��W�<�A�[���H~ ��f��}���qVLn�����{�=4��r&��W|����C-�cz����w\�)�V���������!�E��@�u��Q`	-�saŁ�&K	�������G����f�K]%����e�G~'e���V}��d'E��w��*k�jS��{dn=/lB�]L�Rp
M�MLQ^~_�q��󴻘G��T\Ub�2P����D�/
5�b<�W��1�B�+D��y\�����9��)�����=%G �;�/���y:�>�8�|��j�׾�{�H�ʴY�R�G�%2N�""�K��bg@2l�$�1
G��_lG[�S��EUn�F����f79o>���5Ɲ����-{���A4��R�e���ٸA5}2$��؜h��R����I0`[?��l�*6.���9����4�=g�F,�~�]��e�v�`��N��ug���Px�!��.�� �C�-�"���" �)�~�cu`�o��t�^nT<)�� f�<W�ΐ/>QmU=
5��#�����OG(|���ma�q����b����?�/���������$q��݈Z�!�?��b�5F��%�SE��+�V��[^F
s�Q,NH�V䕔9%#�L.(
����X+�q$,X�:�؊<Ǜ����z��ܽZ3�2������b�,@���L��:��:v2X���NmM�&%}X�6h�(�͵V}9�S�X�̻D&���xG������Ӂ���nS�:"��z2	.};���
�_��P��rw���$m�V���1b-M6�>؞�X\S���HbuG�#�x����x�6��l����ۼ��/��<�ź�1�.ˎ���n�� vp�Js��#V��Cۇ�7���
4�?h���@��"�<�-A��'�������"��u���J�����������g_��duXꄦ��U�'����թ��}C E���S5����g�9�z��9�i�L�[�����9���c��i����W���$�������gj�����g����`��W�0�5!uC�Q ���ɝ������XX]C.E�ja�,�0aV"�;�\M+\_���R��-��Crmay��%�l�5�Z�ۅM_�}�	�4��m��O�n,��Y��v��G=#�!R-���	H��t���W~�dl�e'D�9�x��[�~��c�h�z��
�v>(	�}	붡��}�w�hqp�X�\8%,S�bm\r@ݲ�3&:��) ?p�����^�爄G��Ӗ��67���<�-bM�J�qD�e�����g*����G�E��e��S�˻�/D�D��ߏ���#X&�׉�
�Zv�m���.�v�6kBIc̚���i�MU�A�����1�at���U#�5ܾ�lPH{:Sl���	�N��I7Vׅܬ��vlq�jI�D���K;�Ji��Foq�oZ�*&�\��Fˈ����D,Ͻ��zR�l�;�*q�?"��vjP���J�9��^LXG/ł�?Q��H�b=��-A�W9���������_�c5Z\�b�a`�MJ���F!��9���/J�Hg9-��_�/q�AҘ�e��{�!����&�a3�G%�}����C�P�0�5�
T��g�td�3�b�~Q�!�<(C��q��ƭ�9�#�9+`��6���k_i��\�\�/�NZ�7#;�{D�����qo�d�W)��&t�8���u�N�ˬ�dk�m����;��IP﬈�J�]�u�S���$��S�;)?|��m�]�]����˽����'���#֎N��$�+����s0=�Rj+�5�I�7�Ǘ��,sw�Hl�M���M��I)�|TeQ��,����y�W!��t[�#WOc~	�>b����?Y7���L�%�����s=ӗ�@�g�\��)_�ҝ+1��Ͻ�ڪ@��.�s�p�C�/�Z�Z�^���`��O��d��W��dQayN��w�^_�a8�ρA�<�0	���⨼ȡ�J�˨�۵#� ̕OSS+�yJ����`D���)3��f���'���D���'�9w0����
9���ys�NdO�����dCyPO�iQ�an�*u*��%�?�� 1+�ː���g�21p����rߞR�����Mr���G��{)ܡ�/�$�'Ó޷!V�-�J���|wc
ɟ=��Cv�����X1���9��Y�QӁ/pML��[�g�b:˂}��-���=��� C��u�t>���Q�o�!7�ަj=��C�C�]}#�:���bt��#^�Z�b*��c[ι���ږSN�OY�	Uf�|��!&�~�f.�59�n-��)*��k�` ��
/�
*��L:�R6˳��J�9Zꩽx�5T�XL5x�˳�l������p��2�n��z���0�wM����IW�dw��)L����4�v��K���e+���tmz�!��t��"�4yi�hʮ>�G�Aq˯d��I�?A�p��N��X�s�h�S��2@3�Z.�y��ܝUoW���9���6��+n�U��<#O������E�=Vn��Hf���z�:fB?��Ya�� #��n���"CL;lloU�+a:v��A���)�V��#a'E��zq��m�����ͨ��s5���U�@��{`7j<��5<p���T>���,b���R9x_`�)F{H�_����sP��=z�(��q���sO���fj��*g�\��	�'E;�[�8�z�nʄ��.܁$D!{�Ѩ����9���ʱߎh��2\��$6d�J;X+�8��TgK.z�eY�eN�w���ybf�C?��E���:�z�	�i�Ƈ2�����&i���� l��3j��S������A� &qX����Ю?��L%Bi�j�<=?���Q/���ے�,�D3?�� 6��h��	�������Q����}j�-����{��ȸ�y�;����t*5�0�gaM#�dL�T�?�=����6���=��f͈6���F����(���h-&KX_װ���Iƽ7�Ȭ%�&��9xG�W���E�?Qh�/�:/���9!�.��<����л�\�?��� �)�P�4��!�`�4JMmTaPյ�4�N������2�$�9Μ9-P��s���$< ���"ΉƂ2^�Y���sp/MHhU�u��?P��oia���������LM�w���e	O���r��R���̋2�݁��/�7���o�T�飻U������QF�]V�_&�{���g�:x|^,�i�%XpN~1�|��>}�vL	6 ����l�0T�t�:�J�����Āi�ZȞ�������ygy~O *� �7��S�v��������"k���$Ù��ؽ���Ƚ�gmtp|��y��9�ƞ��׶#.�ē��_�^c�*9U�D����{'�B�þ�7+�<�a��xٚJT���07���9�s�7e����.���`$N�p�Ȗ�
h���(�q�1T	E�E����I�~w��^�3�g)��"�{ZfQ͒/5��M�fU�+cG���q.��6b*������u���|����z�`�\�`�'�p0������ƨ
`V�|���Ԝ"�L�=���s	�P�.̟�ʕ"�_$G�8����L�	i0d�0O���,�9�9j������ci�>G���؈�����%����(�sUs��T�(
/	��a���,�&�Α�t@�n]��ĳ���&���a���çq�L�"c�"��b]0U�&z���<�ۇ�=M�T�ۄ���*�/���s \��n���ZV�K�2g�V�a
�Q������͛��\�|?7L��|�T�]8�E+������m�����ιC�a�Kn�$`M��I6�z�1٩Y3g36�6BO[��+p-�<Ź\|������y���l�e`��*m9*V�Ʒ��o���Vߧ���˖�Fѹ�<;�\��[#yi
c�8�Y��CԜ_|=��r{{��{�a�a��T,���O[p-�<1n.����.�!����+}j6W�F0��Ѥ?i��U��^`�z�,�u���$[>R�1�4,�\»�����H'Ǯ�z��d��	���d�!J�M�hi����u��u��rM^�Nd%*H[�7�huV���jā�����,�0_�.J������NnE�{�A�nPm<|`zI����3+��@�}^��ˤ���0v�o��߂��9��Y�����@�!Xm3zB3'kђU�2�����ӾE%�l��3;��iu�"ۤ�Pm�/��[�#��/ꡔF�"�quy�{�06G����.�Y!�\}�
�ŎW��r�e[ۓ�f���5RR]{+b¿d��Ɣ<O̼�֘' �n�v��B$���x�\�g�nSV�%�p�aߠ�,����)p
�?*<z�$���#a��}"z�{�拷ɞ��@m��@$Qu�릤5Z	����{���7uM�o�����$עQ!��v�C~�uR������`:xIyc����xt*�����9F�����g��}9���H��ڹz���ڽ�Axx�U���T�����M���|��?�;�?������2d٣^��rk���d�=���V�W#�U�}eO֣埑؂�dDոޑ��a��nW-�V8�V�=��|���DH��z��f�� W+B�(K�_�C��Wv<(�s�|1~�@!f\��H���(h?#P������Y2F�����v-5�,bZ7Y�Ƥh�Q�ѽ�a��V~+M�k���/RG�J}��-��>[m�����[����`�v-��%R�m� �g�F�8�no���g4_�\��E�� M�;��3S����֪�w_�#ah�Y��˽�#�֛�����\���E������j�u|�
�Y6t �Jƃj����lG.��2ɬ �9�	�p*~x�=�e�w&��B���/����?8����r��c���$Ed�&뵨�"��>��Aa�I<X��b)��$MW�or���~�|��El�������a�f�!-#Ɠ���h��}̅���=�<8]��>���K�o*�D�k'��U���7����fO�c��A]���#1��pi�j(W�(�������R�x�' 	��E$�'�J�0�2l����	J'\E+��,��Q�!p���7���ݥwE{+��j��L�|�S_��78���$����.�-��ۘkXo����R8��<u���uR�*��F~����5��;��Ė#�1���X�ڇ�S���B8���M��S	����EK�JE��O�ԡ�fI����F��(C:��/d�hZr��pc�٩2��7�C��{�w) ��I_4ó�����hsT$ΗـS�b)���w���t�;���-����1Ǟ Gup@�ع�׾����׏�,K�����%����rFb@}Faf�b褭��T�}��8����;��qY�n�N� ���2�9�d�J;g��<�h7�a���O�7_�#s����ϖ��Rd��8vq8^|$)ϓwq�u�|�v���ƨng��rA�Y�K�N����~Il(m��c�T�sm5�˛����sA2-��q����Ga�K��g&������"���g�,yJA"�}�/�w^j���-FSS�e�F4�Mx�;�Q'��yYF3l���m�q:�"͑4���5K�������/n �;�9�i#�B�~g�@y��QUXp����:2���D����28(i�Wϱ�1F�O����Sj!j��T>�k����N��j��!��	>�S�1�6�&�GŦP�o�59��%E�Z$�A��#OWR�>fn@��w/����6�q@n��0�,��<�|��_�R�f>��N�/�C�i��px��+�%vݘl��@��?kmsAň�3�-ש�?�h��&	�J��j�%�o�[)��6@MF����)c%��V-��#ʇ<�[;JCι/cK���_�[��߬[CM������;к��]{��o
|�F us��+����>6H_���xn�7��{�V���^p7���������*՝O����Or]�2�U�g�[bO�6���Ei6���U1��>�ul/��C!,�y��:�m��Pw���k}<$�J
�,˞c���wѢ�)����D{��y�B�3��6�?�����,#!k��)��Bў�>r�14X#a��UwY?&�)�0M�I��A1ոwT�aC�P)gyX��mX~�sn�T�&���|��pf����9����%S�(�&�9�C���8�O���Ed^���Ǩ#rG+�p��m1���.${�����{��f�n��-����CG&�E����dQg�z�����%J�4��= v��%RX�O�2C1����e������ȧ��O�AM�g�'i�Q����J����]XN@���B�rF+t�/���>�b]�Z���5慱�m��\j�)k�m��k�>��Y#s�}FgQ"j����Z�����nu�wAJ�N��nMEߢOƦ8���yH�����?Ҽ�N�#���V(y�4}���Af�N=�itu�]γG���q���c>���A��S�߽��(\}2*z��Y�Z�dh���&��y��y���k�Z(|�I�"���}��9����_wmת�,y��. ��s���|yd����6�{�X]"�kag�=FHw�m���Ъ
:ҽ�`��7�"Q}�!���.lKw	%(Ui� ��U����C��;���˪�� �v�������1��C�&\��b]�D����4ze�����W�w�Up`��וt�l��mG���W��R���C�����y���f��*y���y�� ��gg1/� ��(��b��(\
j�$�V$�)��k��[E�	@���kz��y����0��a�B�
���-����_~��S����l�,�ʕ��������{�����Ȓ�}#�W?K\��$ʔN����|�����������mx���D}�smmey ӂ ��hs���͜���Is�oZm.~U��{��M~��eՊ5���_a$��r���S�
�,Z����!�?>�u8gh�r\�P���''p�.glΡ��>^�תD9 ��¼�*�C|�ý��U@�gYt���-�#��fT�����I��#)�qvC�����������V��lEgJ�����v�|ܪ����հ�]{U��VVG��x��?yK�{�E�;=�a:�u�dh���ro�[�󪬹��-5��:7���pT���8r�ez]{
�w���kK�
/^cx�n�iQ��5�V���y���闊;a�x��!��vkpk?�-J].EW�
���o�û3�W~��v5_�rO��.�����;S�ۨ�5-�CM�J�����rSa0�[�1��j���� ���]��Mm�����~sU�s��|o��������>H@�0e�E�å��W%�!�ޔ%VN]�鹵���|��ˤ~RӨ�J�[������G��c�m$�z���{0�A�=�e���%�,�n�&?�e�}�̉���Y��M��vX�d�`Ň8 S��]a�z�^Mڀ6Y�dnX�s@o$�7�O!1ϊ�������61c�RY��<��N�9>���e_ɂCw���[�c��Te#MZ�v��o��y��q��u�8�p���XgL7N[g�6�8�ᡠg9r �!������I��ۊK!�7P
 �{AM<iJR���ƌ#d)��d�V@1MW�|��Es~���ۋ2�8�RM)��d��dq��N�{����ɜ�
�#n����n����\9�z�9>grmoVj}U$�b���Z�V6evƲf�EB/�Хg��@����Ď�_l}+pP�Gt?ڪ���Q?zW䏖��[;Q�������S!�U�#d�@\G���n2{�}�@NT�?��|��X��WD\<W�K��i�0�L`%bbNU˙!�BPjƛ����@d�1�r���7�i/�ܜ5����!����0����'vn������wuC^�k�LL(B���{/�򣅿��
˸�s��.n0��/��r�i:�v���a���d9���r���?q�;7=�mH��=n�DՍ%�J� ��RϨ�rz���HxA��"`3(*��rd�De��'��t�'����"A�V����uz%��*���̧v3�	��L!���ޢ�f�_>��^��T�cS����q!��������NC�X��l6����/�cG�ڶ�jw�ᕒ������\�Ji���ѬX?�f����:����G�@!(UE���-�۟���i̤����a�,�[5��&��{&.���DM��}����u-�8�9u�`)�+��n_��N2X�_��d^m��>V����G�܋AY��D�pvGB{���0��d��[�7A��"������� �"\��XV;W����k���.����le��+e�.� $���T���yA':S��i\��W�e%L����j�ڊxU��w?��q8<pP�e�,ٹ�]*4W�����h��e�U	���&4�r���z�~3/S+������x<G��h��,An�_���e�'�W#��5�d�i���o������?���.��O�i����>�K�65}$1�n[��Os��t>q��7'͵����̝�����R�Q����味��eWu�2T&K�E���F�@ˍZ-��㗸2K"~�#�ƣ���E�6�'���	���N/��������K��kɸ%Z8G�)q��5|��4�W���~�R��y���BU$��|��Kc����ә 5��[�l�$:@�[��r:�#i�q!���&t}w5�{��L����7�f(L��#��ҩ�f�
�'귲{9�ǩ��� ���R̜�h(�X'}7W	0���Q�6		9��3D����8�HA���yT�]խ'g+����%�E�c���tx@�O���9��%^��Ѵ�_�;�>��t���e�p����2e���_b�b�*���A��z�v�D��E��-)�>�W �*;c��E��2����|�)q8G���q��+<'�l�'�'pW�M^7x�9!.��e+�h3_E�=����A�5���n�BT
�q���7'� �gKB2�5 �;�=�������#.�#X4����NDܰ�4	����G��\ET~u��Z,F��v'�p\�(+�!�2��+4��:�T�c0794S�	��񙔆�q��{���a����yb��R��ϝ�b�M��`:�J�`�^����YaʌZ��_�x�σ�w�-8l��_ã�r&�	%��Ӿ y�\�>�7X���$U��&4��̈́�\��e	f�N,���3�Х�r?�t��dl��r0A��\@�lJY.�����)��4dܧ�f(9�V�����oi:�$B��q�/Gg�ݯ���U��l��<P�
l���,�XK>�N�_���I������Y+�j4�}����D��UҜ,�2~0����@0�P�Gw��$�o������0e��ʻc�;l֎蟕I�6�~�NA����Tv�!�]k[��w�,�U|�P�+���4��p��2�,1�����5����)��#u[ٝ]��`/h���\ȍ���z�h
#Er�N�[�)�'�Y�@�E�^c�x�n����	���J{�Q�������/�P��<��D��A/��'����m����m )D��E��J��ą��u�a:iv���X�'�a�+������~�#7�#.

0#�����Ǝ����$ ��=�P�I~]�/ݏ��c�������{��*�{@T�O>�̲^8�g�Ox������>'�R�΄+Z��j�b,�k���Q>�!�Y%'����͘�M+���Z�sO������@+���e���c(�ͪ�w���F����lӞ!�
���Ͷ�4� J�������G�o�gR �B�d����gOܕ�n;�8j� ���*�B[�</|��ڐۅ�s��T3�Q֫�>t*v���|Gck�%P�¸����k��n�fkni�����+��fR��2�į�KPh�8��*<����@�����Ű3r�gyΙ.���sV�1k/�?��L�e�8�Ut2@�����J�bPE�8�6�ݦ�-S�� ��M*|.I��J;��W$���3h����~�g�����5r7j�IS�I-Շ2=b؄?Ó�iB��I��v�O�]=l)�
�@��~�D��V��<����4��T��D�ȡ�R�R\�GbXM��TVv=�4K�W��.!6��_7Hy��>AK�GxO����=z��*�;&(��{3傆$r�A�'L�n�����.���Ӹ3����fB��U�J���0�p��ք{�.��*-n{�:�8�/�k�c�ϵ=HI��%$�@�e��
��(J|G�}L"�B��٬�P*��
8��;�#���P0~��?l�](���(��mMm�Mj��
�3G�Ξo�s�k�,��"�Q�m�n�Og�ͭ{�X�s�$�tC6�%:2�xg==Y ��
�7�z�;���| �=b��Z	W�Q3,�u)��$;i��|���� ��fX�I[D��~�b3�˃6�ڭ�<V� ���֓p���`��q�-�����6l�0U��4�4�)�sZ&-_Z���C��������o���&�s�2
��j�`�UϪH1���N��0���p�AI9I�����}loevxoFڌ������g~h�cQC�	1Yo}w�]%�|�b�i��KDp��d�MWK�FQ�ѐ) ���6g�")痶~Q�+�_��R��?�����j��zK�9��{��6�"����8��_����h���7q�m�3�#���B/2�}>�o��k@�iyS�{��E���1�.�j$A1�nJ/
+����)��v,_\��n��lIFwk�J^���ʜ������&��*低�ͦ������*Ot�>-�F����I>P�M�l� W}���Uͫ'|򑮫���w� �zЉ��) :��u{��<�vv�a"��b��;�����pM/�O_.�<u7�}}
�I� �;�S޷B�5�鈐�P�5Q��d� +&$��lm��ø�S�;(~I�'��O�� łW�l/��X��kX$u����"�,,�VD�k�>�����Ew*]r�}N^+R}�-���e.��/�<�]�99���zW�S�?��K�\й+R�Z�!�q�O	OY��<�4J ��:b�(��z�8Ӟ3&ENnT�jߺ������2׻%vY*�f��-ː
Gf��I�o��oJA(���[�ժ>۬���p�pI�^�#̓.Ǒ��V�~9�P<�|*DrM�9����)�Q�S�C���A��>\��_�h�$�=5r����A�އ���l]�פ�#[^rZ�0�q9	��4h94�����1ݫ�H#,h)q�	��qƛ��N���~!�c2 ����2�Y���Ҽ"�h�7"�n^�g��gV�5
\E9��u4��骈�b屽���Wgv�,�6yA���P�zvHMpD�:�\���A��׹�����ѭ��w���+�?��V�gc\O��7��ͣ���r���yU�:�E�t�(��/6���l�Q��#H�Q����+E9��!�]��I����j���X���<��q�^+��1=�.TI B�1�PH1�i@0��.�)�d��r;�ok5��E8:��"\�l�4AjF�.�6��¦��s��X���M>�! hW��|:4����$b�����\�b|C��Kc5Vi�V���)ۡ�U�T�̜.��Ƅ���8��A;��Ć�&�hw}cf��>
�Ǣ����ׯR�f4^� ��3��i�d$��lv�0oT�@�U��}qr|&lit�w�Z�q:�Kb@�#��66D(���s���5n�x�k#a	���;��XyKT�����R̲=e������эK�gx�r�t�Ɣ�!V 썼=�q��}P�i�h4M��/��4m�7	}�כQd ���n�����2�R(��~[��`ؤٱ)�K
�;J�;Z�w�LzC�c6׀����^��y�����b���e��]X��|%F�A_2��3C���v��}�R�Ǆz���JF�+Tm�m?:]-��Ѷ���n|l�W�M�.��n��~��k��|��T�F�9����-;6>����S�Q��oˠ�#��������d���U�����NW	���7��[�;��8N�#.��8G7܊�S�F&�'� ��e�ޖ���� � �B�s{(`ˁ	}F�{p�<ZL�|�(3��z������T�|"}��	�e�ws& ��0�YE�+4t.�ې�8��/��m=��4�E�l����1%��*�O�I��2�M����}&��_X8R��|�d�n8�5��d�עn\��Yq��M������"Һ��Z�9�2�ú�J�@�����$�T�[)�]�v���k��ߵW�id��(��2)��N�hv���+����1�>FT��g!n���%�Xg[V�9������<��3na2��xZ׎s5�0��0Lt �ܕ��68�H��8�M�}�/��+�-��W���>-�f�'0��`�3���������۩�ߵ�$�cǞ��IP�vƭ$����z��a�?}��(�s�!���ċ)ZU�ړ�աa�p���6�x2|�tuL�	njM>:���4鉛�cXD�Lj��o��63�!mI�bQi��2�?�_�cJ*E�^�iE>�
���G���|�K����|�U�nS����V�_����˕�3��Dw_�V����Z�/5���f!1Q޶/��x(��լ�$��C��w�r�����͌��ưy/�&��z
��R2G��Tծ���2:�'Z�SU8���l�4�4����G�0�GU*5�5��(�J\�9�%8���օ42M�c*����;h�N�u]Lm/��_U�m;q=�*����nh@2$L����Ҍ�j>�L�B�19��-����^Ӛ0�Go�o��M[ų�8�(�OQ�V����($�������/9<����V\L�Ř�嘙�ۘ�)v�qd�s��h��{>Uy���"���%�O��]��N� \�L��}7a�1���!�wvѓ��e�Iyj�Ś�y�S.�������9����k���W��4]�'K������D"�ˋ
F����Z�(*�$��ݻ��*�`�4ߧQ�O����R��Q�;�3���5-b������SH�� )�XF��؞.V	j�����;����x ֆL��Z�a�C�UН������y�I�gm%�;�}j\�����MА�b�P�W
�:eǳ���"�P�\�U��q�L~�)z����q�e�32H��꽄ޚ��w�(��6�2u�S�u �Ƭ��Xd�,w�*2�jqn�,��b*I���pIZ�қ�xLCs��K<ۃ>�2�����{��>��!�)�Q�	Y����}Wz� ��6E�&;�]C����>,3���itDHZ��:�Zc�)�V��΁�܌{���(�ր��9����N37V�Z�(�@S�3���z��v��Ո3	�dMK+��N��N} a� �K{�z�ٕ+�\T�B�_�vX&���J���ۃ0z<�珸��s�����Ù���s���N��(��w��� �8�� �]-+5u�LX��0P:^lha���1h3�<:��1��uއ������
�5G�%=�B��a��;uI���y�^MP�?�,yh��ʀ'��GV��,��U�N�=�����U7�<�ʹ�l&ɿ2����]�B�9���KeP񤄏�I��H� ���*5�"d��$[�"�S~
xi�`�*4V�&J�(n�?`(鄾C�[QC��}Ǟ�[���Pq�V�9������;��lI�3�W
�ҫL��-c|����l������q�ΝV2���<��Ó]e}��C�"I���E��<LŬ<A��w�k�!�mw���2cՌ���b�q\��-�\Q���f�
�i�|�<�:v��؉���Y�/*� �ەp�K��@�_z��`y#�[G�x�E����s�Y�5�B_�B��b��ف�_�"����A��S{h��us]�R-�{|��j��d�G�;�X*+L���r�r������G5���0� �Ǽ���_�e��gn��?��^���q#=E��	 �b��,)W"ʍ�<�c��S�IX^X�9T-�8
Y���e:FY|�Mo�ׅ{,����>�a��-��t��I;��%�Kę���nK*�p����"h��.���[8���B.!(�S���;}Иr��yV��3�bf�k8cؕJ� ��19��0X��4�V���F���Y��_
��[6�M�����'i���J��*�Wn�����/?�n:�oR�rE�D�W�P�0�0B��i��y��Q�UOv,�<ԗ���ʊ�)}�(���0_ \��9��|���7���<�����f��ʥU�u�f��>��N~�L��x�u;�?��>;5?�z���AE������d]$+B���]W
�ʧ�V��]�q^�h�3��F���ަԈ�r	����pn���|�R����d�J��Y�2�*af�a��9�SAH����O�����Vˏ�B�XEꬿ�`61�50h�����z05�2����y?�+
�ؖIy����謜*��{߷�E�5O�!�de��?z�_`e^�_��R��	�K;K�,ja��$N�2���� ��i��/�Jn�m��:���L]	�2�OP�zz�mF��%\1�IV`�"�oE��&�Й�#
��pC���� �\�r��M�d+ġ_L��u��p���Kb�yŵ�"���Ԋk�=���idf��׸_ԳB�փ��f�1�M��]x�/�')��lۨ�3z{œRs�;`z����rD��j2G�t��Q-�+��������Q��W�2�=�:i�dqŎ��n�+�DpC7	�c�I������ϐ�xЈ}�������:�*��^��IYm�e��q@����u��y���K"ϰ���?�#z���NM�ID�^�@��5��\��9o�+w������T䚼6��Ɨ�B���{��+�����˛�̄sְ¦L{])��<����&>_�"��4q�}�����`�F�(aZW�����m��d�|"�
��Ӆ��Ԭ���u��X�o��a��<U�IB3�^���lBX��#���)2$��^�Cs�O�P>�.bQ}`�5��,}���q�7��αF;>a�c���9�8�W��ܹX��M2y��H	�U-6�W�v���h�����W/>7��� B�l-A��w�Ȓ��P7���W�Kf��_�EC]����A��]��\�x����G&����c�1��t`D�]C�����)�G�}ќ����H�A9J������P�<���`�F�C�2c�"q��t�H��� ��!�c��	���E=NS87}�ls�ƠM��D��b�	O��{�US��y��!��G�/ՙ�D�^�۽���Uc(���/������K�`$Q�Q�О�o+�w�v`r!��a��ٟ4"�V� eR~x߼��į3͢��De�W�����t��Cj�U��վ�)I�J�^�ӿI\�a��j/)lQ����Z������P���k�{�R��7����r�S"*���W�h�����;�`E̴8��@]V2����$��� k�e�N�_%QS��P�y݊;���z�~�e2�W�1f�Aj�Ee�n㖻�-Z�x�J��y�m�<h��scb9����cIm���UC(���W�]�C���۞A�Ҭ����Jeu�co*�qRt
L4�ō��E��tn/��F��c�lUQ-p�w�e�`qM^O~�,���m(��E�oe��^R��f	�w�R�2�^Un"	kn�H�c4Zk?�adH�#PW��dǝ!�t4t�\�|�?��A��&����7%�t����a�Ʋ���'
S�̺�d���hv�o/h�Z$D�zE�W> &#�����I�]�}!x����ЎU��xv�Y�A�1G!J��%]d���;�溆~ �,�4 �I5����d��ZM�U���AFv1v�n1+���}z'h��߸�k��
|'XI�ˍ�Gi$L� Ճ����68��jP���Ժ�� G����{)�����k�_*�Ո��]A$o�aQ	�1��\�Gl�� t�h�y,��N����@��@�!īs����U}���uA���=N ���QyV>��XA694d�]�gV�#�j��sq�g��'O��D-�l1G���!��&'��m[�	aћ����y4s��k~�3h�e�� �5�:�شo�q0�榲H�#�v�� �W,?�(F�4���*1��cY�޽�{�	YQ|md�Ԗ���I����h2��^�B���������\OJ`�?~�����.*��W����x�ӻww�a�t�t�c���&�6���.�l	��󂾇7"�)���W�,��En����ۮ]p�Vmtrb����!��i�t� �WQ��Ͽ��N�)�2����R#.�NMȟlm�D�J�����)rD�ߢ+��sN�� O]�>;�]}8�<�#�;ü��T�/�]q��@�ͅ�7'R�G��7(bIλiO����v՗��F�k|Xp]�a��·O�{��O�ٿ�G�{�����=J��{4�\��:dR�����3]�`�����_z����a��L��v��PL���z2<��O$�b���m��W��".j���v˽��-��]&���1�>P�m�V�٠�S�nS4ȑ����?6	�����ն�x+��G�%.�~u�� ��7�2� �Fǚ�hJ	F�&�T�y�|2�"��u��Q��[{.ٯ:�c2��_m��kW�� ����茕�%�n<=KԽo�5�(YVcn�eB�"�0w��R�����t��g����B=�	XI�Le4����}Y�дˤ��)7&�����zʲ	�![`�\(�ps,���IvN�/)�ϧ.bC,�h;����KQl���Q@. �}�tƁ���o���åم��+�s\ل�o<36�0uRT�^Փl*�%Ú��#�'GI�eOS�������JF���{�u�	2�RRd��3~��'Gc�������ݾ�<�����tg�z"�V?�>D���-�`C�͆2��ׁ�+I]�#Qh��_G��`HH���VT�گ�^?��9E��R�>Ǡ���&kE�&�!�5�����B��0;M��u/#D��i~�aGt9��R��5p����O�w���qߣU��}M�*Q����J9~�3�6�G�r��&�91F���H�ژ�����iX��ýDe�
~�6s"LSa?�����ޒ���ǁF�"��T0ҏg'_uq���@��ap�Cu �\*ǂ���w�H3s��M������6��������Xwj��{�"y�1:7����M����`@4������~<��I	�~u@����V������>h!1����[�L�$c��?GԚ<���̟<�wy�91��EʅOQ���5A�]��]-K��ýec�{� ��ܼ�����4O!��5�LaR�iJvq��P[�m�(n�G�Nh
�!�7�L�>����~��aR%O2"M?^�Z�Á�z2<q�Kٵ�.�L?����� 5(M=�ak�_�o��]x�A |��:e?�}bA�Q���=�~��abЮ$y�(w(~R�՚�S"�}�p:ѩ['DFC/ެ��Zt;�[��3~���ؑ���Q��`@�U��Mj�Z�e�tz�;0�\��9b��֪�Z�	¾vY��H�"�0�!��F�TƄ.ະw�y�
L/����~Y�"j�H�j�@5���j�Vl����Ѭ�cf~d�qu%���(6�\��c�腠������L�A@�#��{S�F�|6�v�/@@'�Wl�`���	�+y���T���Q{�+�>�Y���G|��;�bf�?�l��_�4���{i�z[	g�Q^�|��Y����mx���Z	m�BR~��[.�g�U�S�=7��d<�0��-��D��V0Gժo���˛d��IH@$������͚��!Ϳ�l#�l��Ŕ���XA��}���BS���lku��z�ӎ!u/F���n����X�����FI�ԥS�����h�����H!��p氒U>W�Ϯ��k�1�����L#�{��ۏ �ck	�12AjXn���G�=l��$��(#�];E�Qd�B�y��v���
Z9���/��S%��3�s��XS�-�|�1�� ���*�5&�x�L�&P0���녍	(���5"ݲ������j�eֿ�o��1Y����cH�I�V=���* ���n[����[x#�[9F�T��8^8ٱ	U�%N�S�9ss�D@S�R2k�{��8��o�"P�

����:��Mu��%��v��,	�K;}��1���*Oj�aA�'�|6�V��M�9�ʈ�=��z�kop3��MI��<C�mlH�g��	�5�m�rC��]��/��/7���r��RD5��<JaPq����SlW%��]ה�l���¾�"D$��P�C�N� A5����;`}b�wx~�EM�Re�� 
f����lG�$K&��HC"bj� �g�䎴��0��(Mn���$x�J����\y��=ƍ����~G8?ϦK�D��-�eT$C�Kx���B��"v�P~i�&�͚��vݵ��^��m�h?�ZҢZ�&�c&�q�ބ��w��+]�]�|V�����|��E,?�:9"������[-���}6w'��iDw�I��b.��+p�V���A˦	R�N�H���n�z�c��Ʒ�� ��ߤV�G'��wU�3iU������,�{{�?R�c,�糅>׆����6T,A�g��!}a�kIq��I�n*l�G��A���AD����s����w�ci�,K�A[5�<�=�̐MS��ߺ���B��e2K}���;K����g룖���X�=wN.'�BP�~+ ́��`���{���� ���`�O��x�!�V'N-�!������z��SlyL� 8�A2���֦����)�FHf'�\H�ylSa�3�-�c�.*�p}�j$U\��mf��U��p��l����}2�cGa�oT�����
��m�99?��i�T��#M.�ꕿ�D'��<�R�j����9_�0@��_O�kq�orV��y�i�Oz�{ ��r>� �	ֲ��ӕA�hsI��ɰJ�4al�J%:c�B����61f��;�T����n���R�}�����̈�����z��i~'��Ì*��X� d�8;�瀼��ń���5L��˷8�4#H�Ȥ[Z��$KD�"�8l&x�YY��{a��ު*�7�h�s�ܲ�*����m���6C�w��"���
@��yj=W)Th܁~�ױ%���v��;|��eXCs5���͔�3��C�WzW�|m~�R�M�����}�'B��o�oڞmXT��������x��PF�j^l���Q+D��kH�q�wI��M�M��B4�.����c���_Y�Y�nһSͤV�`ˌ��:�����
���r��O�����J��{�E��6��l��)~YM� �{	�&ll;�z��7*l�(����;�6��+J�G�o^DR��QA��_o
je|z89��g�~AXa���q���
�aFti��u��B�p�[�){+�v�1"U)Z�	ؓ%|�;0#��5~��F�Ϛ�ܳ �*RU/* �9C����*:�ƚ[�� �¸ޗ�����)�����E\m�j�K�|
�U,�����ҒG;��zԶv��a�bK1o�N�����`�/&Wxֺ1�SĎ|��מ�oMJ�fP6O^�M�H�rةňՎ5[r=��%�#��f��
0�
~��k�a+���\d�� v��@�T�M��ZR쇆/�X�2_��C5��c i�^M�X�b����!�/+���C�|��7�G*
.}q����؟����:��ټ|�� ��<�A~/#)��Ts�ِ���<X�ܨn6 k �vޜ禤�ox|-� �OV�� (��V�����0hw��{���lJr<�����Eh��w�X��G�IuNw���HvH�8�y&�n��x/w1CF� "C@��>I�1G��	+UH���
ʆ	�K\��H��[��y1;�<�t���+zw�En�ߪ�H��U�9"�h��3M�ٌI�X�i�_&ӓ�$��*R[߀���:\F��e�ڣ"{U��kd�\����,��zs2�6�,�Ǡ�;ͳ�>�3�𧹹* �r���g��C��g�+���}U[�� �Ƞ���-�Z�|�@ p�#s�of��=��1	G;��U��E���[��4p���M�P�d�;�(qc��3���)���g}����d��8(gǸ�e��G=n�|��	�3-(Ioyd���e�#}"+$�Հ�;k.�?c���5W�N�B��}��$qM~�����L~7-���A�_k��E=�߄Y�<�l,	��������;{j�޼���A�䘻{���5�Z�E$��1�[��NT��v�`����8��� 6&��,y8���iB?;<k��s�uP�߉bd�*�+Rםt�%֭NRM�-�2���p,������ |����_i�H����uw��:_�1�0��D�r�"�XN�ܕK��!���,�%
��sm�7�Yt��� u���L�H�4���?�1�O"�-�Z��S	N���FݬL��o�f��_ȳq/���g��]2)��@�r,�&�bH;�^�d�UE��)�)��p� ������������(�^s.���|�>���Y�^�@�N�%sks��_cQF���V(�[CH�aKT-=M>n$���G�K��%�/'�'�$qp�oex�=ڼo�1��C�N�jEt2��1��C����&w=1t3	�սȑT��XG���3c���r�XU�Q[󔉎�/	m�9	���CxNn	���?B˒�M�gT�W��6˘��\e0Q�ֵDw����Ѩ!��Ua�َxv(&�b�IJy>���G1��1�=�U�Kw���N^-}P�tk��[Ǡ�,sa�lu��}��l-�T�����M˼�_aq"F����\�nDc
�."�Q0�Ġ殯})gߕ�d��A��]k���w���v~�X����{⮧g����Lh��G�'X�J����^��:�\�b����S�D�<����H����m���Hz@��Eg$��уN2�bL�ΰ��Qn�k@D3G>Vk��<9���@��D�o?;���Qz�DG��#��~FX�֠�2�ǖsVE�$T|B�O�#�!<?WD$�������<�w�d{�V�1�µ�M�����r�>�	��+x�c��ڨ�۫y�8h/�fBS7C٬{���~g���J� F���9�e����zQ�̎�	O�=m׫�ݳ�7�K��ɨ�%%�B�����p2=%F/N���f#�A��7!�*�]���;��ZΒ��C	P����	��t�z�j��nks��,BH�s�H.��QUurR��n����ϖ�T�PѰ� �:��.�%$!$iXP�Bq;�Bz�o��6���D	S��;Υ*��<2�G�N���Hg��?$96��>vn�4�vj��Gs�o���dC�{�����yh��~Ȇ�N0��2֦?9o{(f�ܩD)��<�BGbW@GǓŎd���?I��-Ӵ=i�/���i	@@��]���E~�����26��*�ml��⍯�����'����A�JTqi4Һj&��f�����F�q�~>�����sO0��������q�8��w�s�1���i�EF��d<�a;Z�q�7a���E_V�%ݙ+Gs�R�ӁŠү�ax5�	�V�d�+��,��)��e�"ci��n՝1��P�Z^��/���"��3�^�G�o�@L7�w�Nw�|!�Jb7�
7�__�}.,f�e�+�{�
��R�Zl7ʹ�R�l��ҫ���P����g%�HJ���𨅂��T����u�o*���
`G��h!�_�
݇��]*{�O����yPن���1-��A羈,�����λ��O� u����"�1�}}��΁κ��5����n)��1#w{�,��x�׶#b��8���������%|N�QɁ��缙U�0uip� *�~k�;$r�7D�(/r����ʧ��A���Xgp?��Z_"ꛚv�G�����h0<�ٵ��e�v��j�s�H/������4z���B�����^�"�3��U��=˷M{_=�����ݰ���E�Wa�R�"h��8�_����$������L"��J8�[��0�.����Z�L(�s]Bj�����ve�:��F��8@����4�Wｶj�cM��:��Ƣ`d+"p�����g�F�$��4X��(����lhJ���F�c�Q�<�*�ʊ|��o�#�o�s��.�#�t�~��AIy�W�S�����fKh�*3�7�W�r��U,������zEL�(0�R�-@�S���<�p�x�'���������}/���4t:�V���.)��_��-��ѱ�n�@=���*J�c�&��|6��ߗ���.������on0frs`��4�uoQRڊ-����d_�R�Iyiӄ�۹�#S����v��Şz�s���L����Ha�a �P9NF֌/ !R����4��me����a���w�M�\6��޹n�ΑǊ����^)�`��Á;Evz�_�SI���Uƻ4e��%��f�u�JАf���=ǝN�ߓ���ѫz1�����4I3(�9�Z���bR�_:�z�`�p�z�W`~�c�f�"�5�u�Q��ZBS*��7Q�1��]�}�2b�d/�hb��j�Y��TB�ڟw�uo��䔊�WKl�s�3ne�q�"��a�-�j��t�u��l��`]�Jg��_�t��|�vG�������¬]��� h"�`�����z�Qp�%`G��
A��ޯ�r�.�����m���e�y� �O�mX ���x����>?
d8V��~lV'"����e.!�� "�~�)�Bo%�Wŏ�]\�'"BϘ�B���[3d@��gdJ��ߤZ�6� E��K��|���g��y�".�u;�-0JL���"Mno���0����/��ϩ���,���[���Թ/AG�U�樝�3�؄r�����:�o��v�^j��i�_(�X9j�
bh�h:�Zy
a�?�E'Ƞ(ܖ�b��B���`��ŃV�a���V	���~�¿u�0�g��������Du�G�#���8��f����R�Пv]͸�8�Z�֊�e3������夠0�
�����e���?}ʚ�j��y���x��H�E�lq<�Le�P@#A�>�X��K�#�M�I;h����yXhC�h��v7}����0��`Ƶ)�.
Y��0�Yd���B�|���{y���b��]P�	�ёte�2tg ��]�1��[��>qV�wWrA�*�d��\1{p�)R��2!:�Á�,�yy�M������n��>`#��XY1ȴ��Q��C�XM0d¡�P%���������1t2��R/c�=�(���X�������Ӧ5�Ղ(s�KcHCѵ��If��o���w!O���)�������4�gz9�$-�����dL�
����@ci�2���w�ҴY��+��3g9�oi�u�އ�bw�QV
��Z�j�r��b]�PW����)�RX������0��:���I}_1l}�sy[��\�lɷ?�L���F��e�ޕ^��1��ә�i�Z뮗����H�TB8�[�ާ�Fn��S��w�B�Ǖq>���pd�V1Qʋs����{�YH������zt�$�Ŀ�~�X�&�<���7�M�NȤ˻��W��I3)��!)`���+KG*A5�z�������̪��#^�t��wVn$����$DL�e��3�p�<�k�:��|�E�0�ۆA�!w�����)�[�g�Vgc$��Î�un���Q��>�-П�QO���.��NPk���?���r���8�9߭��%�����f��g4�f ��v�Y���$n�VDN'o�Us���w>v���
R�NO��� ]�~���&R�_�X��0��]��u#�����T���z�i��bޖ�f8���-V����a'&��w�{Q7rN��.����׆Ɓ��S��xeXwr̞1��>��F�.EV'�$�YٽG��.������8$U�Ey�zFv���س#B���� ���[9ܘ@M N��C3'�e���C�~r�9��]�G��U�:��N�&��	s|�Ӄ��W�E\{VVG��
��]K�Nu���u+d�s�ϔ��(��A�U�����vϒ��j_�wỲ�]�GŒ~������O�+Ⓣ3a�?$���,�4�L���q�<*Ŕ��1��(��V��ξ:��𳺯R<�\x+l�!f�E�Z�/g� +��W���ĺ�HUg���H�K�nʞ�FL��g[bl-U0�H�|�]�т�:�b��K�↫cZ�$�H*���B�R�_�3��OfA�aZ����:,�Q+�Z;l�s"�U0���Ғ��9��!).n*Հ�.�n�����}��E�?%�V�X�;�k�ybI���2�զ��Q�8�0�Yc�.�2m��1�<�V뚨�MKZ���5=��e�b�ʩ/��Ag-l"amf =I��1}u������|8;�]wnJM�#��?:�Ŋ_�S��N
�DB�87?A�Ƨ��M�-����U@���bUi~M0W�¶�)�d!eN��EP�T�����;�rm5�����!=�}�c�4�5�f�[��\�GS��
iM�\	��|�cǗ��3B��"jbp)z8n���l���+�9:������s>��3�I��i4i�]�
4Sp��p�4e� ��9��9�������Fa.6�[��#w��k6�/��� ��u��4nGwY�������R��a$� SKB9n�5�[:8t�s)N�W�k9'�U��?�F�>�����8V�.������̒�L��5z��z��5��#h����B (qE��z�.�L�!ԩ��X�&��QJ�pV�������m~�|�
��(����KK�y��M�؋t44�D��J���z����x�IP[R%��DQ�Gt�ԀI��rF�l+���VT���V��XK_tM"�7�>@~M�KA�x�u�)W}�V��|VCj�.�%���w~epù��3��O7�cjObK���I=��v85s��;{b�8i�Ea+�#�-ҳSm:;�i{ڃ���s�<��R�D�kB E�Z<����x�_�*�;�m�k�8<��o�kz��v�\V,��Ç�Ǡ^+ ��@3U��*g�WGEX�\!��.�n�&G��Zye�L����i��֭�,Q_n�!���tD�
�tm���'�G(@Y�Տ�-��s�rw�y~��xZ�w���5��Ѳ�%A�A�5-DFx��3�zY�i��-��.6upXLA�����$5Ǣ^?E��� �~��T|���So�!E��ɿ�����D���i	��{AQf�.VF\�y�-�t�ե���n����=�n2�5J�������#��9+L�W���ֵ0iI;u����r����]����4��eWs��F��{Y�yP�(�m��}����Pz ���(�0/�V�?�<FIs�oߘ�M}O����V�Χ��o����r�J]V�}��?|K0�R�A�l6�Ω�I[o��ad�*5��򖮮�H�v�@��d'����F�T*0� �U���z�Ş�+}�W�����5j��I�Riǜ C��	R��T%+��AX'~>��rQ)�6��f� �?�s����/y۠����m�U,;�K��2�ֳ>P���ل��b�G��I*�4q�U������������Znb�S�6^�W�
W�'�Y���
�Q�t���l���i��rb�����S�\�;�934x��#�Zju�[6t�.�c�)��?�ڀm��ڍA�W75�u�k�^ϲW�n>�Otػ//����O  ��Y��|H��<Xq��v^��.�6Ƀ�]�:l>�u���t��'f�'h4F�z�����Nn� �F����NG3I��zD&υ3�)=ᨼ	���=�2wq�w?����FS�[�4 V-��������m4"�]����=��r8��UY���g�)�$p�N�Ii����wah�GT��i�`5�,�Ё���s�C�����m�=�ˌzg�l�/�\R�1��D-ëO�|�:�Ȯ�&޲���J�+�l���/ut���шuCF�XВ~an�MX~��r�Pzy�)kf[\�����Z(�vp���t����N�9��J����l�[�!�4�tcF��j5�A	�����!u�%e��$�285<��,��~us���[���3g!q�hN,�f��Ȅ�>���ֶ��	�*���E����^d��׿E�RPFv"x����x9�Q��h��O�Yd!a�&����{�����8s�O��z����|�}B���([{��' � ��ן�h�<�5���cJ��"7Y��܌�M>�<<���ʊ98��Tu@���r]��L5"S%m���!Ӎe?�	p/V_ ^�7]9ĭ����%{�ߘN^Ч���maٴ�s@�.��6�nv�p�.H�|E֥��A�N�.�����8�\w��Ԋ>�9�Ѭٰ��)�5�۱ ��硇��x<*�'��E2'ƆtVmM
�7�f�Զ�`����d�
zuD&���yDؿ�f���۠S!:�����O�a��/\FF��ь�k8�f�(�k�H�i��6��P��w��R��j4���\̆)����._f`7c*�3���>c�o�����^,`^�#���v6�k�t��	z��j��J�K���-��^�i�xđ���-J7�,E��x�S�n%��;W�Y���x�����h/~���D�p���cvO��-��Ң1�"�Bݗ@��=�T<���L1Š�O��
R��/�j��:��K�c��I>�?ń������cHC�窘�����:�D �j �p'~���c�GJ��V�&�+M��L�~{�[�K]�(�I?[��o�L:�;�
�1�̝\��\�@��k��p�3��]c��ڐ�l���j�<μ%�L��Y�3z��"��J�� �������N6��_�ԓ�^Ò4A/��h��&���;#"cޒtr��v�9	q��$�0y�}�4^!9��KAd3\1���zl]{�ؚR�d���i���b,rVZ[Q}��ť����8M��Gep[��y⥭�2�2��T�o,�O&�[���k��3�ףR��l��8��}�=}c�*���LXd���aE[|#�J�~�5&�_��'��:8Ҧ �4���n�]�0��#��\Q�ǁ/"�$w�
�p,�Z�b�s��W.D�^G����U����������AV#���h;�&��I[k�j�$~R����+��{=?%���4�FJ��g�luo/�?Uݖ�z%�W�ؚ��a>Fb���R޳���4���g���C���x���;�ۮ�[�o���T�èP�y��MLR��i#������<�O�W��QxS��~p�����0�n�:&����U#���&,�2��`�g��|@���]�(�Z��S�9����1l�!�I4�1�~�/`�kv�k�d��]`T`U��L*��5^m���6+]]��xb�4�S���{a�rV{==Ѧ��(y�a)�8�����F	z��˨?ԝ2W�L��+���.�c��gee��7/�V�Wu>0��)Ę�J�������{[�=wߌY]Z�����\Y��'�i�s��
n��c����$��b-*�c�k�&,����0z�I�u>P%��<yD\מ�WΈ�ɤ5�ˬ�'�Y4�����,����w���ET<�x��`��Zf	�X�@i{��6�k9g�5|����W�C�pT��4���p;+_X�iڤ�H�P5�Z��^ W9Χ�&&`�Ul���W���d�-���Q�?�<��߀y O�[[Zp�:~��)VO����2�U׾^�!�Ćī}��]m��������U�!�̂�����{ ���+������"���,�zx)��`N<KWڲ<P�736�K
�m�D��`���<���������f�!�-"�h��^�p�v�4���k���b_XS,|�[���8^��)]���$���Ӛ3Z�N�?'ȷf�=�X!HS�)|֚�)��8eT9'��5Ͱ�(�UX
�ws���ߺ�]�]��G��� ��w���n-�?��y\�'�㱓F�铹��}�1���˄����/�q�0��F���@E-,7M�/]��3�^-g��^X�=��Ϭ�Z9 �|����U�K�w���,������Dh�:#�E�ZrM`��@�`�i��zk-�I@��Ѐw'��0�̀��o�˺�l�Ø����kE���!Fc�k1儊ie#%넸�t|$��٠K+��À<$kc&_"K�0��q���+h9�)�XٞM�w�Y�$��=յNh؜2V����>�!�E�Nh}���ȝ+s�Af���	]TjN_L��ǁ�Si��{���#N'9Cts�"XQ?��f;��wIt0�e[�* �I��{��LZƹ��C��H�4$�j�k"7��׺c�Jh�]H�-Xo�*^��8����}��؁}��8� ��qn�K��I3T1+�Y�s(e��w ���q��0��hk��Y���IQ�r�BŻ�={5|�^������WF�1v���4b>����������a{�����M΢b�؄����w0����&L�ߝ\�W΋��b�
�A�'Zި��R��yQ8�B�j�����t�:���O%�G��Ĳ�RE�5>�JηВ= ��1������Z"��y�W
=��Uq��0�lCyǚ��˅s�����r��E��i*/��S���Y��DX���C�dJ0�҄�()�O{@(���E� 鞋�m�p���	���rL:�����4֠h�&`M�5���i�ݜ
O�.�컛n�RϺ�"҇�)k5��[����c�n_\d^�EO�LM
ًe�G�R�\$w7�{�B�5es35�7A^�!�� �˻!�`�J�3+��	{0���ؚ%FY�`B����'�/2�g2$PS>>x2:��3��ٴ.\`V�1�٥bȩ���O�4�pϓ�0�K����A��4q7�n��}}˨�]AT	��s�}��)t,�=Ӹ�����}����HQ)���J����V�Dhp3�'�)�J+����+�q�������JY��zs�'�]�\ۋz��B����zF��EEx\j�dS��'	 ��X�VXh�
ԋ[����Z�\�څ<���D'p�s���)�$��Gl� ��j�V�;��������S��hu���1���.Ha_��m���j4�Y�Bb���_�iUYX]�:�`���y��Acƻ;7&NS�%�����R|��]�{���-���G2���ur�f��:]���icG�����
^��*o]�H{�QM�y����,��	r�$3�� �ϻ�C�mY�4ܗ�ox�[���mqo��iJ�ݕ1�(�[��뀡	!p�3&�Ԭ�؍ IM��Ep\�b7��a�F��b�*��I��h�
�w�S����2���W�n�U�m$�~Z ��@p)�>�1΁��>F�4� �uNo8ܔ� �)+S�57��Q	qf���}
X��Z�ȟhM����N�(�Wof)(��Z�b\�8����W���.;�Cn�=B���6p̿����㡦�]�{�\�m4��l�J!>/!�L)�odho�S�k��T��+=�w��S��_=�右#2���I�M�xOn2>��91�X=�j� L��C�������i	�\vO���[��\e9@����C�(0����	�>B���x�	��D&�L��e.��/
d�riQ�9R�s����4b���&���C���4M)zn���2��XhU�J�����T��=�@�?�x]�э$A5��^��qO�k��@�qzOr)/�/k���ҩ� �;�N�ƶ�q�*'��V�&-�. ����̆i,N43^���=Z�5_���6���HX3M�\�7�ޱ����?l��RD�&'<�3�-��Bs~�w�}X�4���m�`͎��r_���R�`�c��q�y��a�Qwcr��4VHy�B�R���S�;�:4O�r)�j��m�PI�S�2s�H�v���@z_2i۽ԇ�X�N��D����w ���||��gB3�B���\54�?����j����`R�M ��g�A�!��,�P���>���;yԼ��b ��'w�Y���,ʐ� �M��Ӻ�M�TA5������il�g�J���{�h�uN�R%�O[2`���N�݈���Y���'P��鹲�ca��9���Zh'�a=	)�tP6�����P-�r�S�{`Yʙ�v<�5��tU��d�RxO4����
5�v�{��>��Q��s�B}�MB���PÑ�G�T��p·9��Dl��l��,�`�/=i��G���2b�ܩۘ�Y�=C�ڑj�®n�T�H�2{���84h�7Ւb
=e�@�`?�����^�պ`��ySR�Q��R���3���p$fC���z�R��p��w/�=S��lp�N����hS!FV�*XQPwhܺB]4B\�}�0^�tJQ�4wQ ��4iS�W�bz��+�!J���2���?����E�x�Ur�����MI��^��4�0��ㆷCk�U�p�Irȩ
���h�R�=˞Q�bS̘���F�1��ɑ��ZTP��睫nx���VK�2��.ؤ�c���.�e�r ��W��0��<�y�W��&��QZ���6�[��MJ�r�S���av~T_Hإ�)�Tb�O c�<�:�$���Z�6�gzB=�s�{&�̓�?��UauA�/F-ɒ��Y�������,�;ʄ�J�Z�Th�!�&���6ڢ�.�&�ǝ�8�:�]gͯ�w=u��<�uF�3�k[��u��èStc �η7��E�p�i����>6��'o~P4�����R��k���(���n��w2B�h�b)k�9V�<C:�t��D��c���$�h��`q���2 �@הߛ�c��t׷gX[a>>�|vLL�����#�~	��i���Q+�"���+v'�W!�f��[���@����pge�z�zRwH]��8[#�6�녮ܖϟ��`��!�� <z{>�ҷ-0�~z����PO�7sTU��0)o �<`�=������> \VE���Q�u]o�Ьr?�W���>U\@,t2�\�e#���O�cs�RCZ<�K?|�eM#	�o�*���/�����>跕������c���h���P5�aH%|R�q��?��+2��6���JIkA9UL��@h+x(xꜟA�^�z#��l%ߝ���E�*s���t�TP�,K�s��;�E-�>0+c�:��Xn�/��.xL��3E�۟q�Bw/ޗa�{Ϲ���U����o���z��nM[�z���'/|N��X@NN
M�5:�#�Ah��Ẑ��`�j�:tR:GXuj��k6���P�PV,�5�*[�j������q���>�`c�W��[�W�#�d�����nlRܡ�O{+�=4V��m�`�"�'c����KN�gw���-$X��}6h$�u4۴$^����NuH����B�Ғ����p���X��'˷���ȭ|�,�]z%�&�n�z�ͯsz0^,�=)��mv�`�g�����O���5�n�qw��y�Hy��$v!P�-Q��G�@�b�&P��V0�R�o 8)�*��4J3��N�xl�\�墕������#��!�U-A|��|�ct>4N�g;�A͋���$�NP�{��S��Y��9�_�`�	Sv�%m"�����8���0��-�_-hi-9P��Q�a�rO'�ҷ�+:�7���fܢ����ۜ=��B����KnR��L��g�W��GJ6�x��m]E��=��8�ڱ����}P����z�@t�8����T�*a����{�gU]���^ظ0it1������������t�*�\1Ѽ���;|�	Z0e��������f�B`������xtp�L����	S��kd5̴�$��=���ר�:9�i�E�ۭ���u���?��7Z����h����/�u6�2�>����VT�����4�c��H�IVALHI���֓�v+t C�.o�I8Vש�,�ݻ܏P��F�a���(huM�Y������=�`O/o;g���o�e�L�{u�^���j������s.�����b�������2D:3tҿ���	
ӸGC�~\�w���!��:���J/�*	R�xy����ZAe�*~������"�l�c����/E�Q��Y�\��(x��]A�h��C�y�:�"��$������9�d��]��"�^/`}� ��������J�`�{�]�Yč,jUb��W~�~ŝ���L�W����>f($�G�d�W�8{��9��끀`�WE*�ܘK|�R�w�rB���4:�zL�B�+�X����*�@��R'���d�tC"[$���r�vͻ��nb��RAC�����L5�q�ϑ\k����Z8�r�3���Q�;��_g�����G5�J������=?l�:S�݉=��\��_'��a<�B��,�v���5P�S�v3��4^�AUZ��PKr��2�6�M�|ޡ-�}���Db%��eE�n�~�M� +K�D�^`L�����4�G+q?�Z����~Y���s�
�ز�畗 M{�uC͇��́�m���ȲϏ��G,����y���q�K,ֈ]���0v�LO-��.C����[U�C��(�����[���kP�^@����wav���=�i��=�������Cd9&£�u��}�FDϒ^h�\��?�O��V'���Ϫ�X>x(�*���]�����L�O8�ĩ��-*��F�
~�1�ow5A��r�&�Ж��h6�w��S�^�,��h�r�̜u����[�[���%�WJ���d`Aܵe+�SL��fN�*�0���꒾��Y���`�P�h��&���*E�_��^����Lv����<�;����iRf��a��3�����&�F4�Y@l�p�h����&��06�����k6/�r8��x#t��7��nL#[{ �Puotr0��Dfy��Xi��jq^py�/Gg�O�F�!+?��+5��χ��'���)ȹ�[*��I� ��@��͘��h��H�L��앮	����L��j�gJk� ��J�M��ː>L�vE��,^��0���ʓ1v�|1L�N5�R��
�_F�b�g.�ѝ�f��c�$���&��g�!���9���B���`��1��tJ��tQ0�lc	�R���;��oK@SP�d�3R�/�d�k
���(A�ч���j6���b�����*��S�S�8��v������ӨqNoݕ�Bn��?���拃����Vr��_�8+���,���-�Gv�X�yG��@�>鋕}v!�1X�W�C6V�t�e�jn�"5n�
@3�ι���&��4�ɊZ��}����Ke5�Mo��'���^!�M�<`�A�&`][�H����0,��r�2���s�q�)�2ڈ��~3����#�n1��J��I��dN��y��x$r��[�**�r�&i.��HX�P�o���q�H��,�0DB����Ӯ^����<��_P%ǌ��A��o4�^YF���C�M��˂{}�]C����	N��A6�L�R] �iTD���[]�8�a�ғ�������o�+n0�� 7W�Gb_s\`�e��p�}M��?:��|�$J'<C�:�C�G��8�Y��jQB����d#����\��������m�H`�#4 I&��Gv������#�
왂I���[��uH�|��Q(t"'����m�%s4GZ��yR^{AX�M�ĩ?$����ɩ>	+�w0�����>A���5����?d������ۗ�b&��y ��Wɀ�bA���HF���VU�I�SC.��f��<������@��v���Q��>K�����:��>Ӹ�R��!�xTm�Fą��a<�t��y�m���*�d��X�����B�3����1��Nk�>kk��mGw~�|���`�[7�C�����?�F8�!�n��ř��״�	~GK�A]͌df�Je,C�v��b@���x����0��
<�-�d���J��c&�k	�N2��h7j��)�ǏIR�W�7�ɮ�'��;��^R�����C�
���K%l�r�=� ���%56G�*G�k��k䒔y;f��U�?��!'��_>D%A�-�+Zh�d�#\������}
 �!e�&�('��F�3������$�k�=��"9�8#�NE���Q6lf�V��O����"�?���0`���g��>V|R�P�(m~ie�_;��;�Hy,j�kgM�O4D>���EXl��lt	�̬�R�ڗ��Y�6\��p�u���G���1��Y�������c�?����X{���d� ��ڧ�$��'�,����.8S���l٬�������k�a��L��3��8�!v�1Y4�J�FD�5m�J}�%�B I�*�F�lq�wV膗��5͌��ZBƟ�2�>��o�W,�dC��C���~Z�!|�����T���Om6�G�ά���9@wW��L O�3��H�E��Vs����NS-ȹp#�X��.Ana1j V��� ���5up�qN̆ٔ-F�Jz���ܢ�}PS�~�*�r�:�]���5�Rl�K���6t����߹a�Q���A��Yx5Fr�	�*�=�&��	�%�5AP��w�4��.�9�7dk�����D���0mA���1�'�w_`suM��f�E�EB�|�l6�k��5�5��=��|��7�Nߗ�6���s҈ُ�,�L̅�l�N����6�n���t�����v>&ʢ=�R�A�R�6�w#B�/��-���E����}/�QYt�w���pf��`T�O$��S����}b	=�H��~�P+�^c��X��鿘�jh���VU���<�!�8�VZ�ҹ�n�E�����7f�2�P���	��H��$EQ8Ok�1��h�(�/�,��3��Ojۜ��g2gD�*aTZe>�-A��ǵ�]�	�C��Ā��C�;�yg�D��g]	���}���8�D���K��!�.yQ�)�?󯻬p�
��6,�	�7�U�-��ž��O��k�Jڷx�;*t�N:ʉ�?��Փ��gk7�s§U/�D��B[����X�.[̤���'p��PM��N�z�7}�}�on�:enk-��5 ��],^���1�{|�C�!����cF���q+�a����`��F}��F������Ĵ͒󁿆/��D�D���;����b�ݢܺ�YJ�%Dw�՚�P�}-���W:`�fz76z/� 9W�5ݝ���d�.�g��A���x)A·'<o�0�ax	�ê;�Οe%{`�ݛ�E=�jkwQ�i����ƷH��2�(�ۚ����7���/�_�"Qk���L��I݉ @��O{cyF��>IP���ڜ ��*���'U�.���Qtβ���]�c��dYLM<P�Mq�'SB���q�Z%��!GU�js�.3�u��C>\E����P�O���CĐK��U�>l: ����WY�` ��Ɩ4n�!�mQ󭱶�~�ԅM�+ѳ�@-��N΅c�P���˪6��^rӍ��tm/�Hy&S� �Ub�Omk��?�������B	R.ː����nw���0,�!�in������Dx��#*~`;�		�4?ŉC�U8p��5EXj@���`� �+�A�s��6�b��H���f�������S{�[���(�B��$W+��$�dr�/���p�abo�*<���\d8�8�o���X��UX��%lP���fz�&ڿ�#�'��sP�c2�q�b���D�ҵd�g�8%�D��0�h��Ѯ���[;D*1��F�[����_!��K��Sz��%�GKI����3O����Q���$���_���5��3���MM5T���?>%��]B�9����K^�����W��@�EHjT��(�d𼣺�w`;�]���v��.�i��w����@��^�Ʈ�p�?LY�I�	7��_N&۽��R��\< ���0�F�A,���,����$Ӵs���>͍�ʭ�2iNV���Q����" ����$����*��(����G�G�"�G���[{CU�� �ߊ��j�o�^�`r?h��Pi�ziʺ(������V�k�
���Z7���0�������v���xf >j^̠?�"_�F�����}���jl���<YB�{&��i�h���M�@���A/�=�k���=�5�:0�Q�q��c���JR�]�L4��L)h���+$4��->a�NU�o}��hC�#/��L"DN�8�ч��ɓ6�EP'�0�-
k�͸��0
ӈ�6��CV]���CG�ҮV��_���0�f�p��#��~��c���q,ȑ�&�U
��ri�Մ����r|��?Z@��e���C�HjA� j�T�i���)�e�/!쉰��8���-�#����|=�7����Lb����_��hv'
�#�K��h�|��{��T�oGUKE���
��hI���E�R���(��IzO���$N:��(�ݐ�]����}������C&�,��]��W�4��x���+a�T3y�c�i���j_}���^��)��U�@���}�Z�C�^<=W�l "H����w^�l����q���e%	�d�Q�cC+խ��Xn�M���r�a��X�g镼H@�]�5a�%/eڹKm(���Q���Lո������%����yɢ
�50{S���l��:d٤���P�+�v9��N��V�P�I`��@�v�RY������zCJ���Z�)��zG<�BOfB\�$.�Әl��όb�� *�ҕ�f�����N��*�6!r7�����a�Y��L�h�b@r�I�A������~��1!n=�z߫�&�kP�`���UP�-��t�t͆�	�w�_,Y����a�&yo�]��ٚ�vpp��b;�K}_�2D��L9�8~��"s8�R�˩���7�ؚ-Rʰ	�B��1:��[/���� �.@�*�B�#�͛%߰Ll�,��)���}R|2���	���h�Md\(EO�6�ƴV�oL�a8��c�R��%��X�q�I�w�����"��4\VyYnX��9E�zQ~�9�ka�����?攁��1H;�o7�5���Fށ�ix-�A{w^��P��`t� �Ԅh��f���G�Q%�!�INb�~�5px+���)V�H3�׽��َ_�W7I�Ld�b� ��җ��&a0���)N�cr^�� #S��s%���c��,tFS�F�ΦΏy����l1겔�B�;A�?��G����
my��TՇ!�a�{ob�Y��V�WcC�C��PW��_�ۭArK�&���U��/�r�SPn���m����⒋u\ڌ�$*/W��S�a@��򪼺	av�)�>�\�x�eu�9�֧K�)��|���;|�O������Gh��V�q1Q��(��j�`9���`� �Wk�U�i	ܧR��4Q���L�)�q6�3x��I%��}N<���Xm��Ҍ�Y�������>䋚1��|^�Ǩ2�
Q��h�7c*��r렋��Vj�fU���л�U_
���qG���_ �F[0�N���rm�s�Y�44�ɭ�vWo��r���_	Ɔݴ�B��8É*�d��C�:bq {�b�t#K��a�X<=�
+�7�z��a�GΧ|U�'�����iPp���bK2��8��9HN��[=���}��3��0�u`'�R�@�k��|޴��-�Z�%e+�Ft��\tـ�mbμ��V��5�I+�����.��Y%��q(�Gd�U\���q{�v�!���'�_ W�/���^�8��+��㧬Mj���S<⼔#2r)�e�x>���*�)����+���|����#��~��:�v��/A��� AV�>�۷�� �[5�_	F@*т,�4�MQ�f��Y�	��R���f)��������*9Fi1:xz��w�qII���e�H��Dfj(.C�fay��)4�Kл�v��s~9������匨����:N,`�c^�d󛬣>ވ�1րD�_���y�������Fl�*����.?�w%���!���ݸ"$J����eq�+Pi�5��G����'�]X˻,l3��vm�+zO,k]db�H�@�*&pT�:�^gcB�n��2pyP=y��_}̦BԱ"�ٓ��&��9=&�)-��9��3=jhmR[���8���8���4������@bV���W�N��G��s��S��V�J	�4,r�yn�zQ1�c�_{xv�e�����u��RrQs܍��ee��/2נ
�D��!g #�ú�D��Q�y����H�QV�Ǣb�!�c]�L�	��+��#����wq�}ە�;U�����N���ރ6x}\�g��E=}/�Y(��$�)������{���s���a=���dv�yV�6
�\ �v�G���w;�k'�G�D]	]�"lel�viZ��(�:�:����f\��T�ֲ,.R��o�a��t�11��&[�� n<��h��ټlW̺FUs>RN��b6���<���S7�hxWD'�Q�PK���羕@��=�&�h�/����Z# ����a-��%s���`b?��F�:�NEoM�1+іx��\�a;'A]�d4PhY*cp��H� ��)��ݒ遀�{�*�IE֑f=� k';�� 촟���N��^5�;��E}��9p�W����(��dv�6S�������FSW��6goU'�ae������U��^��Pl/�"����&�\�!	�!�]@]��0��8�|*���9�Y:J�m���Q/�"Q\h�n�]_^��q#fʓ���]G i�{��+Ү�cB�
�
�������=�������i8>��TCv�=yF�kUoEb��"�i|#�gv]� �K_�vj���U$A�\,�N�%/Rz��,�H����=�Q]{����ll"��\�k��#A�6ے;�T9�u��j� _��e�:I��� � Jx���ιm�ž6����<��l� �.�sC�j���}G!�Oӥ_�&��$k(x+n��l��G�ܮ /{Cu<O�IG������LWc��͓LaZq�8K&��U����S���{x�����|u{���F��p�a@�,M�S�?��H=4	�5'�<�$8N���_��OQa��S������z��y�}[�S
j4J4�df�HN�0'QLѮ�j7o��zBU��b��(	���?�����L�-�h������i��INg{�{�\o	7�E���.XJ��A�ǌ�"2��>��Qj��� 2������`�()`U�yt��o��J.+D:��4��� �r�d�?wq͸���&o�s�� �\�c\�E�4Ĭ�W]������muYNH������A0��z�敋%�/9���-y���?��]��&Լ80���+K�	d�V�/~[��?2�
/���8G
B�]T���u�{4�D bf�hI�[Yk�y:p��{�v��Gj�W���ړ�n�����Uj���ŸJ�2����t�y�B�v�%�?l��Ou��_mJU6ja�ĭo�Njr�rV���F��
��s�b��K���
;���O���-NZN�@#uB�m�5�����'�WL�I�pLT�k���F�Js���h�����*�w�e��֔��a�]�t�D�7��]���$����5��;V����.󆍘�W��Q5���l��(iK~!�� �fϯ��}@��Yj�3jx�9��A�%��񚱸�z�+��+��|��������!/Oi�Ą|�?0�#H$���k��"��Ԑ.)���5'�	U�֭E���P^9:)kX�M����*X�mO�k���R�e�d	������J�"K�|z棕����곶��Y�^��3.���������:p_܇� h�Ԣ�u���<c����t�G�pP�M�|����C��[�X9V6[��Eާ�]����>G[���lC�h>�No�]�yw�����Ⱥ<�>
�ٗ*�Y7�@;'���A�^$����$/(�].�G�~Ko��}�1�������|�֖��,��7b�	�td����b��)��:1W������W�@I��ϽC�C�����_`�������D�����/*M�ڱTl�G��}jI�Þ8^����ܕ��N�Hz#��,��|��
�����ز���[A)'�.-qev|Ҵ�� >�]Y��3��-�?m��e�x���xӞ��^PE����q�I�V'P�AXJ�W;��ڤ�2�x^�X6I�w#���E�a��75��/��7��N�4�:Q��5|��%�Wn��imS��!PD�����#��2T-���9�lsf���3V(��$��Yv�����@Hk��K��FN�`s0�^>1��1:���P�)��X�(o��i(��t%3q,�8@�Ĩޚ/JȔ!���P�.��*=�}�y��&�B���@��.��ً���5��'"r�2��-Uf��Pl�u��c�/8sxTD��]Ro
��&�S�MA�j��*Y�ï�sY>�6���r���JZ$t���H��?O�+)o�|�3��P�j=(��Gf��:
�3�s���I,%��q�e08��� �K�]SS�g^��@�}�d�0��C5)������^g�:�,Xb�Yq�T���l��\'	��,�⼢��b*?�UJ�ԍ����OU�
9,�P������^b�$� �
�3�`ZQ��K[�b<���/�:�: 1@��y�E>D��\��M��˝�X�E�ė�֍��T�g=�SYe3w�, J�w3`�4�����N�b�|�frb �$�pa��G:��	���^Վ}�_�w�G��E�,�>�̔Y��8�/ND��v�p*Ό��螳�ޠ!=�#)ƴb+��jh[�̑��O'Wa�,k���p��g���Y�i�;��@�eX��q�}�∭^�D�ͱrvA�Qq�
���i�NIm���Τ��B��r�W�l�r�ع��A���HE׎�ˇ�(*
�y���e�.ҁ�����4S�#����JEڹ,�kMYlA��� ��r��������KC�d��q�0��:3~��ܜ���ƍ�s��n/l��㚘���ldz�
i�����:�X|Z��1���sr�3?��-�R��>��nG�"��y�Z �d�\;	, �?�^]�T-���!�N������Pxk� 槻F�,������P�o���\iWXb�2���c[��ѮȚiP��T	�`J�'qu�S6�����C��Lv)�yK��X�/>6�r�2�,��'�ₖQ����v����=n�P��ㆭ��+2w�����y�\E��u|IVS���Seԃ��kBVvq6Kyz6��
�$bt�,���;�V\����V[�$u��ø:,���]�(y!w�+I!j�N�����bɅ����'��9<�.��~��~�Z�[�z�6���k��W�u{�Gi^��C77�޽�_ɓA^�͓�]�Y�LϦ{o*u��Z�l_X(��~|ZHtr+�mF�s?�|�Q�Mr��0�>��1��#O{uwAk�5h�z�n�Z�`��i6?Ͻ?���#f��C���nv��ES�Ҹ��]A{����LF���`��7��h�rۜ�|0~C��
��l��t��O*�[�ڟ}@��bOr��ԁ�-z�휧��� �TZ�N@��*�� Ss�ˑ{E��<�ֲ8T��R��&�����S%��CW�H:��N�_`-+�V�_q���5+�I��]I�7��ι�{��I 3����dJ�Q"g�8�W�.����Qx`����@Oء������|O!�<��X�Ф5_E��4�y_U��j��Z7nӱ]�9QƂ����E<���L��Z�$���`v�77��V&;ޞ0㳇�<�k߭�x�k7�A��K|X�p3<�x6~�|3��
fz�g,��O�s!���m���?@�C�z���i�09��|�:g���$E;7��w�P�^�����O؀�tF4���r����[�?0x�K��WJ�J2ə�C�ƛ[l�G�i4�UL�8�l�g�a t�ͧl�
��O`rjG�Ҵ,�̩t��Fr��e(i�׳��X��[f�b*�ծ`�W��q�EE�/�D�a���CYؠ�.C�ܰ�$֢�=N��Ѯ#
}�.�����[ �c�"��,[�DM���!;��pW6v����[���W��|�k�  ��{K�oud��4�TL~;�Q:һ��7���K��6=�	�?��z&������؆$�JI�fF��Z3^G��u��Xa���&f_O��y�vMe�r/�&J	e'�^l.��\�-Srͣ�F�Zg�v�%ؼ���?K�N��a�0�?��XP���d���b:\��mO&;H���y��y>����*B���\H͌иT�PS�2����.7_��X���<*�a �G��iV��5rhUT3ՇF�>���s.\(�|�(���������2;K���K"8%-3
�����j�ԅ�?���¾�BJ����1X#�fx��ZQ5`t/8;�#5�p� 9Q��h�n:N#�3�;t'��4��7��a8��A�I�&��:�������EM��~�n����#��O=]pȊG@��d�� Z8�K�%{iO(����a��tP����Xq�0ha�fg�;��hx��t#G�q !�~������NZ皬��X��,
f�lQ���	k�2u�� w��$z�y�;�Xػ ��n��3����N���ܶ���{7��xuh� wz���e��X��6���Eif2�3��@~��U��-�O/��	F�qF���D�	ߣa_t�FI�BXJ��o�ӈå ��N@I�9g��L؉���S��
&��S�{��g�t�3������o#v{���.�����Gu�N7�4�8�E�ܕxw�l�ڞ�
P�M�FN7�8g-l=�v�@�wH/3e�}�/�7ُ�-���@c��h�X-���s����*�}�)Ķ���s�'�Y�e����BV��-����^�m�n�e�x��|�������b�gǳ�Èg!`���Sw�S��v�������Xc�e���~�p]����HaU�tol������ ��&s7'��#w�H����罿Yr�yL�9P[v!Ѵ���� V��3JQ�X9w��] q��0��h{�x��Pϻ���
��L~��^W� ����3�w�������w��׿56�#��ؤ��X��:���&��-�3�Ӕ�7�2�K�KڕB�+`m �Bh�ʇ�������{�RߛE�y��"h�YD��I�Q�����eN?qou�����h����Z���M�����.+�Re']c�m�ތ\
���+�j9��;�n�_3��liA�g3`�Ty$%�3�k�[���#�z_z���*�ڰ�X�h#�m�nuF	u�N�yr72�����L��<��q�^�f���l��[��tB�����USv��D�uD������Xp��ڢ<��#H��^+l�uĂfrI��'��95c�KS��"�Zߺ��Pߤ�B�kէ��4�(�%�2S�&8�̄�[�zW�aG�"�ynL�ƛ���ke�!�j���	�k��!d�"�<"��0����*�$>}�t��88��H����r�����������ͫ�@�'�m~�*�����0�Isl-�{3�}�(�a,��;�t		�h�� � VwL�>�T
N��J3k�S+��q�\TJ'����H �7�	����+�`���w��¯���%���KW�
x�w�������i���!Nn@bU�p#$�*2E�n����F�c���ǧ9���o��ok�/V�Ef�m��$Kz���G^����^r�|ۘ��Z�u
9�N&�����XsI�[�ف�"�%ra�
fw[ӓz�]�Q�϶fve�c?)nh1�+��E ��ʯ/=�^i�f�VP�V͇�(G��Q�@*����� ��h��Gb��j��܎,N�XP����47>P�� ����yT#m˿����D�vkJ�x?՝�8�2?�ZfU֛�K�F���|�?�0D�����q�?�߉=�y ��Φ/E�a2]�g����
���i���f�~G>�����+�w�AJ����W��G��'u��~�Ig�7�~�:�i�d���°ne�`���v��a���U��<i�&�v���K��� �d��0Aٖ��lJ���U��K���}��n�x�:�p�{���Q����7�$��3q},J���;��Ѻ��fZ)��<�ɀ�`A��#Dp�\߂.7ڹ&Q	S�̀R�ۈ�j�� 6	�X���h{�y��Xa�p����� Ԍ��ݲSnŔC����;�2F{������$}�v��f��]�&,�Nt��+����|{أ�zS2c%&T<[���4;h��滲Xď������~7�+DJ+�����>���'l҄l^��E�L��9�0=@?|���_� �~�B=8�U�F��D�2��L���	ٷQh�g��C��r8�}�3�aL�I��X�
�ƫ����
��Ad���m��{d�*���*���"��)io��9�>Jw\|.�/�W8�������2��e�Tw�x`�Pc���J��Ō4���M�f��t�n?>�"�X�[ �����VzkN���Y+��ճ޷Y�n
�+��j9�����v7�B�0�Pc����ǾVB�����w�2{U�!�^�mnSL+�!х���i�e���d<�AyM�=�V�h$�����tt�mH9�@�\FB_�]�&%�]�<=�!�e���!4煉��!�{+U�?�{}3IP�^�.u�5����d�l �r}�;u� �#�-�Hϩ�tD�Y\��/����E�<-Ɇn*���a��qzM�ډ_�+���(7����OS�-r��c��fIag��<�c^��3lG��7���o�]����\�zX]S�ZO�w2{���F�7e���!���4ϢgN�Ґ�Qה���9�!�8���/�H���~��b�� ]�O#k���s,��΅�.U�060]���\�~|IP~x��$����=��J`X�p�F�ޤ�����NH���ٔ�6����]\��q�oF�ھ��ч{����@S1Js���*��]�������@G+�jnVJ.A+7���퀰�q���e9 �e�x�0fDa�d ��J,���o�l������B�8?i(%�����%��n�Ic�Pͼ�zn�e���i�сH����нvw� �ǲ��.EU��p�&J���
b��_�i�[z[�+��<���ҫX��8�Ϲ?���!�tO����K�ʁ5�K���T��J3�p�ҋ�K��K��G��u�Ll�&�r�T��� R0������Dú���St�{?�ߨn�k�Q�xCUBf�z'�ݸ��n�nī�{sǼ�����? �="��d��#3V���/E��7zg!X���}��0�"	7-JM�u�Per�*�
�������Ӊl��Ii1��1�ן8C���6�ԨP��Չ 8h�o�#��v����Aۊ�;0]�|�%Rlg"��ٶr@�$�	v��ޠ�?Y�p>b���.��b?6�N
I>3�5�1
2��C�Z!�u+��)$�r���
��x����������d�#�|�G��sD�u^�V"�'�K�GF㚡EH���
����-g�P�_�LHh����-~���}^�<4u�����\(��*,y�dO�tmJ�VLBc�'�[���݁�|�H%��M�c�<J����c��;�%���9�xIg��=� 72h�������(F��ە��V׊$Be#i�m_��+r����ĩ��B2�n�'�Srla_-��Q�V���g�����)v�N^5��-GqQ��}�StK�H�޹`��I���MO��y,G�Y�Q1���:a���D�<B3�!B��ғ(|ϕ��H�O��{e��<Y=�ȕ w&�śt�	������A�܅R�X`&��~���!��+�*�웇�C���`G�l�Zf$`�8x��]���FLzw�U҄sŐKu�CoA���IK�to�T�h'PgQ���d�j���>@�Ϗ0KG���ޖ��J�F7��A�\����������Y��n�D��ma쇖��Q���[D���i;�d��Z�����ȫ�H'�f�}��'K�����@ݷ�\N�"E���}��n�@� �Œ�'uZJ�)[��2\D`
A��gH [a{)
�b G�эZHZ�E�m����{��l�wd�F3�d�g�s}%ܑ��/�wq���u����ܝ�l�B���>]8�H0���r_�Rf�`�g��K7"}�WU��W}@te�n���}�T)���ѸE�{?��0�$sT���Le�zdҳ�|�h�E,�Ơ�2�{�;Dy���p㺺� ��Ă�T�L��[l9|�%Y�������Ͻ8U�_}�ˇ={ �^��O�m��$iLI @��s�����kB&�!c�ZD/�����m�v&�թWԱ`��)yaj=�yW�bB�l)F���ew�0J�]Ծ$�e䈁�+WM��k$�AQ��}������'8�n�=���!��ZnR�Wn��D`�|`��芿�?|�͹6�w���a�P�ߵ|�AI|}�Y�|fޣ��T��t�{�g!��0[��������l�-���=��N��;�6'�����珈7�����YoF{d�O.<�d�3�u�u" O�g%�Q����qi2mHϊU~�X ��٣�;mQ�:��[�`>sn{Ȅ#�|�k�<�>��C����L�)�
�X��Nj<<Nwv��]�V����G?uVB��7Ӵ�ɏ��c'����v���h���� .�	�z5�I��c1L�>HB�]��g�e[:y]d �F��0�JP�Z��*|?�I]3��6��䵬��3[-�hm���_��[o| S��=��/���/?��1�����<AӋe3D5:�0�9[���q{2*0�eȽ8般��m.�]�o2Ǥ:��.�uA��W�M��Y×�b�A_v�p��j�L:�$�L+������9Dۤ�G��{&����2�>�0�X��6���& v��oo�,����3������|p�/���ii�F�4�*V�)��\
T��❱���gG
uѕ3���F2}d��H�N�1(�%:��@� ;k�!�'�p|I���
_e��x'�s\P�z�L�5
�ofP�%� E�e�'IV0/yB��TK�6�x�HBj�1��h�����e�iPHO��ģ̲zu���b���ִ�Ƒ�Cȑ��a>���A:��,|4�|(O�@�vyLZ�u�֤t�6���XB\�OKpE�׮h����Ku�
�bD?��X�Q��Ә?��G���r���z�%�
Y9'�Xx&w�h ����l��6Z�5Vu��}^���E`�I�=�>������ֽSx�H�'��ɭt�9�����aI+M�X_�
o�	�)����(d�)IΤ�E��V����{T��\���)󽎽T��x<��<�}u�������(+M�|��c�ŝ@���R�1��h��猴����sj�B҇�K5t���()n_�O�������u6T���j�z7E��_����MG�Ai;��؄��*��b!���Z����#����F�n&!>�ҕ���-m�T���!�ډ������"��SN.�gT�D�ð.}'#�Yţ���7
�d�=�̪���}sOP����:z5 ��m��=���@p��gaY������P)�D�͘�t:��fTm� q�,0D^#������3���|�4]g��U�`��u5�^֟�Y!��1�H7�XZ��V�'��n�>W���������X�O��NL	��wO��������ߡ,ܣ�>X�і6ig�"g$j��	߰��*+^�H�O�P��橇r�TC��J�*���
�^P7Ȥ�������D1����\`T�5��a�m}?_$�Py�F�]`;���СS�;a���O&�
�����iӷ�(i�� �u��4橋j��#��oa.��i����*�ِ���w��j����ׄR�(�O��bt�1���%}�Y�t��"#Ov$�=+�EɔLR�U?Q�5�E�L �t��ڥ�XC�0���R��ej| |��rĔ�m����KPO�����^��㶸7�mO�+��xh��h��Md��sŋě_��ݣ���ڜ{)���6f�M�	�\�5�a<�A*Z ɢ�3�ڋh)��H����?�%���G�&�%J��Vk�?��_t����������"��SƔhH^]��j�����&T3�jk��.��Kiۚh�g�-L�.��eFD>c/M��x�A*�]֫K�Y4lOť��<޶\t��ԥL[�|�+�h��Q�Q� ���AC{l�(�죡�*P�OQ�}�z����-���@̍�7J�aO��B���
[�?��S�oV��9������Y�Q(�p�L};��3�Nf;��DZ��{��cuFen�	�8�^��1�&���`3��U0x6��ޜE�~%�𘎷�Zү8��I�8�R���.�6c�u�q�yک��%Q��*x��H.��N���ݪ��Ć?����&� ��UK`Xw��i;o�����D�wq��]�e-͡�R�������+�\W������S��-�o�����)<c��g3?=��T�[�f�ڥ ں�����j�*n�"
�C8QGT���P���a�3�Ϡ���� �r�_4�T4��S:�k��uW�����۹���		S���5��M��^ؕV�����[�-�"���o	e��x��MF�h��E���]�b0Z��vkg�ȥn��,8Y��%{�֍��z�r{� ��t���4�@[Y/R��D;0W�������GyV�8�.�+��2V�j
��GI�V�T����M`v�a��qy�l�,Ǫn���r��Z���疽B�E�<���b���j׭�M�����}E��t������=H������K���BĦ�g�E+�F5L �&�G=�>�F�ae�츔p�!b���Hs����f��m7PW42�����Ҡ������'�/3+S@�5}(�H���,k���C5����-�.�R۠�21"�~~>%�S���ɣL1bv�$h��_��
c��?����;.}F��A�(��RP8�)B���܉ZH|�S�ߡKW%
0ȣH�#o`�[��.@GjQ����m�,�R�3�O��w/N=�&��ur�����f����� R�0򹾀 ���'� RR߃W e2[
sK���o\o(X�f��H~��aQ���)3�'�t)]�"�����_!r"(����Ď�f����O�	I��!"��	�۵�l?�������"�R�˧����Ժy�Y�`�| �����6S���q�j�C�g��+ܩv/;��3g��%�O<2�O}�h���}B�R�e����]��^ק+�,կ'��e2���	�V>{7�Љ3�'�Lc ߐ#H�&�=���~�!	n �@&�j�Y90G���(qz/X�n2��[��J��n:|�	k�<5�e~�.0��ԟS�]��/+��:h^���:BD�N�5�߲)���ԳU��땆3��[�'�I@�w�f���]9���r�5gq��I�m�e� ��ϓA+��4�=
,
uPު+D��tj����f��q�T2�!��T�J]&�4�jŉ���Ȝws���� c�̲Q|�]
͔#�F�u<
m�ϴY+�W�b�������6Zu�_=x&�+�����<U�1Y޿�K�&H�4���>/�kP*�Z�E���D�z�\f;��И��BXẂq�q	b�.(Pm����ca����g�_�6\P�[e���ۊ���WawN*����)�Wk+��X.$�eA��F�$ϔ|��Y[�:Z���~�%F��)�o/5�q�܂��F,�fC� ��z���r���(��%ц���IK�8y]��M�B�+�K[�Vr��N+���ݩ:���B�ھ��AV���r��
=�_�\s���tݕ�!��	��d2�'2����&�R��*8�/
9O8�J�f|����m��B�_�z�+��3�û�G̊�2���=�x������d}�}��G5�x��{\���{��YĿk��$�M�\r5p���٬^Um)��C�.L�m�VD;�����Х\W����Q��J�zW���S�8�j�1��Y�Ѳ4a6#Er�Wl�w�_z.�����n���u�\�ja�Gw�$�G��쟌'�#��e�k�\B��n-�>a�����ͳ]p`����V:�n�9�f��زG���G⟈�!��i��M6�a�L(9`wo�l�`�PCݤ˛���pM����e��ř(\��eD�Y�!t��%�u��G�&xaY��������{[P��|�-�(o����Ｌ�뙤�8X�"�����󒼍��C�P6VB|5�l�9ܶ��_�E��X(�<��խ�ԼŲq��S7�n#8K�R�<!�_���?}�E��d�
��+$�Sx&�`9�̎�E`N.<J�d��[�����>�2�K�K6R)�+���t��y����;LU���9�����`pH���u��=�s�#�﹘����<x����R�]��Fq�ZE58W�Юq'J��f����Tg�^�h���`�i ?�D���>t������@Ia���\���)���@rX���;���[��v1����WW�㹸���Z�{ĺևӿ�u��}*t��lC��*'�O�āI��f[:h$��'�!�J���z��b>��ҏ��	�Dˋ�X��h{Z~��c�傻��Z;{�'�����`���sw}تL�o�bb ���OZ�)�F�\�L��	A-��z�l>0y15�4bxഈ(T�z P� �XO�.@k�=y�o`�&Z��f������q���K���ޡݺ�~��}�w�ǂz��^��8�>��O����
��c�c�`���{r�#h���D=�3R`�xj��
�AXܥ�b�Ѐ�f8��3��-�yΔژk��@mX^J�~�'�O��>o3�;~N^9�}~�给'�CD�?��m=���l��B5�;6��U����(�3àv" Y�#������`P�
(p�?3��
ov��� J�?O`�����y�u��:ƎU*��5P>`U4�����/�5� �Q������D�u��y�����z�G��^��Ul�F�g>h�߼ʹ���dt͵��@4G�n�?�jg��\���Ae.g��)K�BE0��{K�~�*�����������ݹ��@���=d&�[c"�s�$t}���<Y����T��2�5�gz#	]�����"�ȅ��
0cq�����g8`)Z���{f��f�+g1=x�CY�Tu�뵥ܨp�����MV�����_�!�h)|���
����%;�Х,�jI�2o!�a���O,��@��������*T����$�z����Ɲ2:���VQ��g_�H�r,�K��U�D�������t��x���.�Gi��4��D(�N� kz?3ύ�ۣBe�5��u�<П�N\�9�H(9�u�/�Y��/뫾�.��_`vm�x%��7o�u���KY���(��8����(���,���~ �7�#��7�C��Bqg���v�,7����WEw�1Aj��k�������8�b��W��*[�䑖3w��T�5�h��>��F���emS�+&��J�*�#ͧ*�8��)�0m���pKn��v=����p��P�/κp��	:4d`P��Uw酓�����,W���ި�:S�U��*�������g�'���'I���v�$���w��6�O���~t���u�^Ns�W7R�/)I����R�X�y#�z�\�ڌ�e�L�w��;x�(���h��w��;�ժ�S��+hҸ:e�J 7��ٳ�%
�������l�m��4mN��߯��+���jכ��|4��GX�[���\��-P�Jn���Չm62_�r��|(�� n�K��2|���N���b}�"��H�ɢV�5��9�6]��=(Ҥ �i��D\0t�g]<~�7�+	+{�K�5e_q��Wd�� d��C �R�`b�w�����w���1�J�_��;��|�G�d����������!���4�4����--�<'�G�̐�֡��+r )4B�HGԼ���#	�� �����Ē���^�p�m���嫥�Q��:WTO�8��Å���w3`Ҹ\"����<���k�d���k��ӶnQ��6�H�eY"�$�!���_>�S����j#��b�(����!�c ���s[�����L0&/�樇�o#�Ҧ\��r��c�J��Q�nc��]�.ǧus�=P������֕U������m^��]��5�k#q����oh),�rݚ�Fo��qq�'D%���Pq:�6����w�?��E��<������W|�H���NK���o��."LW�C���g�S�Ĝ���}(={F�/fA�YX����C'R�h�a8�h=W	C̻|��^�v��]7��³ǐ�!q����KnʰP�����:uF��4�!�S�y��������M�`�7��O�^�a�q5ـ��N�;�Ꙅ�rÌ	ȍ��q=#�|&���ThQ$6@f?�W|�L��|H+I�BH*�2����q2�Ɇ*1���;��<z�pE�֫½^8D���C L��\�k*sO�}�X�[���'p8���Z|K�Ǧr5LP��X�{����)�.���0u-"�����:�3:Փ
�u;$#��c?�����S	�`�|�%̓*�4&�V�
[�9!0S��n~�n�D�'}�w�(���v�-����\���ob��v}&@��D;IY�
�<�®Rn�i|c�2زm�-c*ۻ8Z;���W����\=��̫�~z Ɣ؁�=RMcw��2�M~r�k�I��P-x(n��J�Փy */�̑�)B��6�{��5�P��}/igb���)g�#��N%����������I}2\1?F�py�x�P�r�7AMaá֔���*���v16T��A����r��-/�n�{����a�z��d�Zh�U�n�b��i͆	����0���L��4
;Xt�X����́躊~��>��2��&f-,�`�#t*�#�Oݻ����n�`}���C��ۿͷc��.�XE��j��=|�Ml��'R�F�u����o���u�!Š΀��ю6d�w�j�Q���X����q�b�_�YQ�:lP(8i���R�n܍K^��}FL5���ܑ,��4�m�ȸzL&������EJ���t�F�m��}HT3�DZU��=�H�Qk������������ؼ�
�7,Od9�#7��]�hݍ�������`��g/��t��YK8�@'�0���y�T,��*�;� �vm��Lc�������ߢ+�p ��_K�K#0<�!%�F���1(]4�������2�RY�c�w����B�v}�YhMZF�)�y刞���vK���x�����ռ�HAr�L�Au�g�T��]y��[G����e�ӕ/�D�9J���4A��k<�ȭ 7�wT��Z`i��xM4%�e? �8$�\���e#�P庻���ȴӈ{�z���-7Ӳh�镭EV|N7-E{Y�to���RVnVrs4$;�4M.ĦLZ�˘{OS�SHגOQw��H��KM\�Vւ~�S�m����Fhڍ�RJBc�����\e>�ŭ����~���P��T5�H��#O�(y=�;n2��f��(��M�&9#]K�n��d�{L"!E�(<�[xmǱ��HD�<�p-�p�*T��d������U���3=.�� (�9�	c�s�i#M��!��[���s����Z]��{	%q��p�<�B���ңcL?D��j�|���������;U�l�>m��Q�ZǏ8�pL��]0���V�%�ק�� ��0D��yڱ�1
�k 	���w�5��f9�w�WDi]X���j"	&U���H8����5��l��Y�P�yt9��!�D�T%�u��֡�&N��Rm5���7�AL�b��/XZ�O�_$��ƘA/"7��:�M;���w~ M.3D.j��;t&�l��J�6�!By���#`>�sax�eu�5?am3�_�3�A��s]zJ:�����ٖ!+��n�KV�R��:���,q�!R�ob�}p���_e���։���z.��]|c,`���@�Ws������r.|H�P.xZξ6�����r6�k���te7����jB)�i�N�Q��ʻ<``��J�S��|9�O|�3(�	|"Ř����သ�,���,�`�O曞≟=&�2�
�Y�Tɶ��RV���랝����k��::��F���Q�#�����e��<|�q1�+g`-�K�OҚ��|H*��nz�����/��W��tL��jx�sQ�i���"��w��� M]5��5���gNw�z��n��y�W0k����
ocC%YNu&�'�M[�q�Ts��.m��?v�!F�I6��?k>��`e�J !����[�A�h"0���<�ݯa���38va��Z��.z��0JP$��^�#J'W�At��XQx=ݒp���K�lZ�-�t�q��d
��_����Ў$�p��
!���V�.-���y��Pp�c6���7�%.\�$> q�0H;���ɨ��-��+�"?���6O$z�{���� E+#�����B ��y3��8�vֺ�\����k��3l p���S��h2{=f��D��=�_�x��mL*Gv���D�i��u�  )��%���h$/��U��2��[7��,�v���Z�����ہ�@�)܊�鿂bxqh�����:\P����k>`�uʐ��ߪ���aķ\�7�[�)r�(�t9���]|{֫�Y�f4AVK�,��Hu*�mY���N	��qvA�\.��tޖT��w<� ގm���6s�#��|��'�^����X���#\5o���(��ΧĄK3x����Fd;D�,B���m���'=�L����C�*aO[��9���a��y�/�T&�W���>x��hD�f�=3�n�����*z��|g�-Mw�֧JY����R8ૌ1��W�9�{�5*���5�z��,Z� ���x} ���3/��T+��DJz�e�����B��r*�!��²b��SjRn�q
�&�]�e��V�w��x{Թ�N:�;�
s�+�I_�x֡��In?����V<�}���mۦ�=B�c��6�'/��>�z��v"�v� ��X�Rum���q�'�:4��3wi��������ر)�+��hY��
�s��dH��T�"T�\d�d��[����Q�����q%��̙���(�@Y'�M�b�kd�e;]OX��Xz�]�l��)oIfv�`ق�؝��CA�$E�D4�u~|��8���Զ��3�௉��u��Pϛ,P6�ʯz�&J���Z��,j����Po�f��t<d70�? ��Y��?�� ��R���ÛRg˒ʫ<��[F �F�9��u���TD��8��}U>��o͘�c���mC@6���79w{�5�M[���%$m���t�n���
����o��e}�AT����ΌKl�C��l�L=�A���4���K"zyx��^z�s�M�`��Y����o�So���u��{\��E��	���O{T���W��"�h.9ﬔ�"ͳV��YSI)�K2�UR[�\
�D�H�}�W�G���cFS�O��{/3Q�RAsyq�rnI�"�9�h�VO��}�ě���������D6���aQ��"�;���h�8j{�MKWp��(7�Or|jW�Re�~�Z���?���3G�rS�㨾+j����xV�j8�^F�C)x0�^�+g|=�j�7�s��hc���y�aU���Q�G���2�-_��Or�T��OV�#��YB8�!�?����C�ː@���n=��8�"��Տ�]�~��ҢVv���k�@~<5ܽbQ��Τ�(�������cPĠ;�6O�L�k���]�o$�E�d29)Yz��ء;��u�l��<�ig�?���>_B>�Ó	���j_"��t1��P����l>s��a��:G��lL���=Y#���}�(�=g���D�]����J-�g���̛�sl\��g[�`Q1�w��¨�NZ���{Y�z���m�T�V�xi� ����R��  eX���`5y`�(�����%�g��3c��{�˝�{˨%�(�<;C�j�mU9e�oR����!#·�'oP���1^0 �3B��>B! ���@��,�N~h&RFh�ţ��fJ�_�'���^{�W���^��d!� �5l�p>�T\5�$���Zr���������t)��ns�*\"[��v[Ѹ|KP�R,�tK��ejW�T�Ai������0�1h:��R�@�~���y�4kF'��lz�P�F��Tx �t�9�'���B$+���0��Tn��BR�u�g��Va����Å#u�@L��=�2��Yd��M�e�̱���g'�f���r|��p>E�0.=�L�4��?�R�r
l�d����;�sU�M�4��v��Ys�y�8(���D�u
�Y���p]�@ ]=SĒJ���Kl1[tdpx.������/�,'���r� AR���x5�
�i(s�oU�>)�M�^eO�X��i�A�l�.H5 ���f٠��ήr�k1�5��`Έ�_ �S�l�U��V�B��l�8�5��/�3���#��/�����=z���Z��u}��ꓯUW�]���zC�PJ��s<~�q�� ֤������qW�b?���L�5U_p���4u�b�X���P�$־��B�H�~�	6����SR�n�m ����*�kW�_OۜPT8Y`Er����x�aAN�^ve�>��!�'���O����^������Z8� ��$�u`��&�D%���Y�C_�\ζ�ly�H�����ܴy�M�EϹ��a'�r[m�I��b>EA�{ɉ����9=s��+��W?���N_K6�K8K����ŉ`{(����ʷ��ך��g�q��s�A_���AP�"��MQ�9!�IAm��t��}�YWҥ.�����Q1�+��p95�'��.w�&>qU�\i����"x]���!9t�����t� ��=���6��b3<�<�e��*�	�̖�HR�s++R E58�.]�㠟�h�r>7�E߳�Xf6�(�
N��"�^.؇��ê�>�f���6A�2��qa��L���H��cA�J��PG��>B霑ĉFOVg,2���X��+ .�LtpE.6�ݿ`�X�R�sm�@	9ga؉�s�����{�-ڗA�
��H+�"�Mj�JT:�s'�`nŜ�����Z�N�.6�s��[���DA�'�	I[y5nɕ#֋aXޮ-�[�,U^��� ��)J�� -���ˉ�e~�����\����Z�uD �q/�-1��dx���Wv�<0���p�H`o�g*�Q�+xh���l3��Z>{�T0���&�.q��:�I���� c���{�5#�EE{$�dK� ��!X�3_�@����f���n�(E�x"��̭��`�j��#�/�n?O\}<�t����f<��ի�����>������&���[��V%N�0O
3�h�yڵ�y��u[I��'=v�x4 .�jrlN�l�ĝ�o�3���I�.�:�g��B��]k���-9Q�,�R����W��s��
�D�)���z�rN3K��j��,U�n`xn;z�z�����km?C��<~�(�Ƒ�ܵ��
G{��De(��+�_�4�RI� ݂�8�Ǹ�;Y+�G`f<g+���M1-
���;U��44{[������q�$Ϩ�S�s����Ѳ_0�����{��!�5��d�0`*v���_����fV�{��%xDb�_�f-���,	�)�X���z��@�9��|]���4,�4r��]�����t������S=��UVcݰ?/�Pa�**h-wD�V4����Ǭ�W�f�6��q�~��ͽd��y�5,�:����zV5lM��:�1��1ht*zoBՎ�YY��
���*�]�q�V*g�BV�Ġ6ς`�,?���r�zqkY��Mu��n��-7�E���A#j>E�d�͒�w��,7��@�u�y�+:�X<����U!ğ�	&Zn�g��$���(��z�0�6Nn�j�u�1���iNb,������CXD��C$��y%��k�~�q��l�,�[ZK��IWFh��#k*���S��t`Z��*c��'���CØ�igUĬmw����z��߫y�){q����Y��}����\|����m-m�eX<��k:OV��v�#�f��������ۡN<1K�ݻ�Mz�9s~�R,�1���J}h���V��� ͲS�]+(I	9�!'K�$̈́�&��d��R!��&����G�'�y��-����()�4��C�:�|���	 M�Z���nbYt
��i�&��9�ʞ֤έ]Ѫk�R�MECf�E�ypHC�R�9��ˁ���yi�C����+��S
Mq�{�3�z�ޭ-��Nbz�Ka��T� �>��)|�U�}mjx|0��@K!��<o�t���~��!�Zm-�%����Zo������(���]��j0��R��	U ����L���ƽzW>\{�/��"5�=��t�9�σz����R��6� �ߊȻ�5��3v6hbZ�quʄ.�ڞ̞'�)m횘N;�+9s���>;�d9 WT�Ve���'�+�N�A+��E�>x.ٟÎU�6�JV�������g�I �;�/�ɝT,���Qcֺt�~��d-��dh.�K�Q�ֽv�>'d�l%�%0PnTYh�v�JZ�ߋ���C�[�����|�bo�G�7#_s���Hr��%X���v�`��Fy;��vt�K�f�^�M3�w'�����1S'� �z�
�fb�/��fOL5%����@w���q{{����^#��d.eGDX&��� 1`���|X R]9:�婜S��x��M����-��D��3Y��*!^e$�ް��L�e;�~�;�	Ū���A8���6�������@�O�֛���Y����(��H<���7��%�ҭ���nSbM��}��+�*�߁W|�zܵm�����?*��K)�䕙-Nq�8A�	>{H��W��Jb�^ĳ��}ܞ�.{PI��L����Mt!��e"�Ĺ2ӳ����V��# �@$%�9i׭�e�o@#�zi)uޑ�GV�N�[F��Ied�����բI��?/�_5�4)��?��>6�vҰ�L�#�ގ �C��W�A�ޑ����2��(O����'b�����kJ5="���*^�_,�6 eˠ��<_�/�mΝ���.�$��f�O�#�W�F�P^�&�%9ʔx���d����9�'_�f�Ow$�<˵4S?���xC&:����geڰ�Db<�|���ʉ{S��> �H�7���ƀ��"Z��@Ʀě0:�36?��_��Nr2���a���f}�aw�=�?w����њ)��&V1������'�v�ub�2��?��=�D�&���e�6z���Mn��� �=8q[�6XFh�@��4-�B\�?3p0��'�hKl�,�بD�E��\lI�kO��	��T^�`��%��-���*�T|��L(�oP�jrJ֦��"~�B�C���oZQ!��ԏ(ynW@�\>pG�4Q�kC`:��	�&���˶��L
v�Z��-�Su��*Gr��@m|���K��|��vu=+Q�)�����ZjZ��H�i��U�7�|U�n>�1�3����4��v9�ĒA�F<���=އ�q~?B���q[�+{�����"�4c75w4���X���o�_#�0_��U�8�XC����L��w��B��L��);ϵ�z6%���%��p#*�z���Sn�pM��:_��d��z�<j���������Q��)*��o���H�Z'37�=���?�pO�@��86���T��;<�N��+%��.���휿��FdyuG���F�/'߆JKUC5/�I\�(\N;G�%����,�k���qmے���$;S�`�  }��)��1cB�1s�����i��r�Ё{`\�g;�t>}D��a�Zc#H��5�A���%� �?�.pX �^%�b�l��� DY�2��5H�~Z��~��I��H/�ً(�����;�"�J��jywa���d�p�����K�AW�dS�,<�S���@C~��v�ĈsE��b���m�cT��XP�k�����ʿeϙPޤ����%�H:��N^���~ܘ�HX��P��VI�W�"�ކ�X�|����`��{>p4ε�z����#z�p��|��O��Nݕ�L*Ƕ��o���ݩ���GqC��u�<��u"��F�;}��Ä��*<0��m�4u���pꧥ^���򫦖LZ��Ǻy#�`b�O��6}���&��8��Q0�T<�ֶ�y�����5�ͳU�Ji۾:����m����>�_Q����]�i�:�˦����9�{j�yT��鶹�Ar��{i�䥰���ʯ2�f�!ⶼo,c$�7�M�"�$�d��B��V+L������t��B�4�v�ڊt^�k�ڹ�soc�=��2���ɭ�qt�(GKe��&����E��UP�Y���L;�0V�M��P�t�!�"�ӗ�o���o�$�;�M�(���7�'�|����X0:���<�� �yFF�qHPT�D �2���"Z��&q���ȱ��1b���~:9�O��b�.�2�C�_[���4��dx2M�R2#{
�)[ϩS!U������ a�iĜ��(�c�-n1!3W2�����MCe��	e܂=l�>�[B�T���9������P9�x֦Ř1iۙ�u��1��gZ�g9�<�-v��Q�v��o3½��D�k�1��o�*G39��^��E·�����V��kH}����@�����օ��w����&
yfEi���U�%^\ N����l`+�cQ�c��˲�h3��[w�>|�����yp�ST�%CU��Xy��vL
Tw-JQ�~�b1kp;��1�Է�K���N����]��;	�!V�w&7ݚG}WL�Kt�+��/!,)��:}�ׂ��q��6�Y���ZW(��>�5�?r�T���q��ƅ�/�����g�:��7�V����2�g�7���Ki$H��^3Xs*{�t3v�K�Z�q�r���5%!�4��:��r�yq?: �Bv��Ԭ�0�;W5a�l��z�O1�sy/m��%Rz��G��ڗ�)Y�Mm��H�L����DO7��p�6s8b�!U{]�:�}7U\�-���.���A��1�Ljí��e�7�iR�&�����^�&�	�-�a� �0��hsПՄkga�g����8���.p�ѡ䈂<�wjJZRٚ�] ��Ios0��W�����6Ω6<�}�-�;���%��h��%�K�7<�C@��rަ��bf� 3�8(�1Ý>�����ҏ#����L���~�k���T�G��#��E)A0M(U����B��C��z�y_�Q��&����O`�:)��(��=��C���E���C��ü��X�5�ō��������^�����l�G<&�+;�9�+������n�@��	F���b_�޿{��,L��g^^D@��W9�ӿ� ����8^��
NjpC�����5�"D\���Aa���+�����;�J�h2��ͩ�)�UX��XJ�{E�^��iqd��oŋ�h���ygf��˯o�Z�٣�a^�V�UqSd�X�\Č���X�e~o�vb�FƤ�5����
��+����d�ʂξި]O'�P�����|���i�N��o�*2�I�q+H$_1`��)$�9�_=�}9����6�����+���*�0l��q�)|uA���n�gt�"��s����J���x5iWx��Y��S��.�Y��ƗX]���~��?$�O�U���&��������y�bb.dn�4Ր�ync4��S�j����_q�D��� l�Iǁ�P�����r0_��5)��)Mn,��>ڨt�7�䂩<3K7�j���2dz�q���cb�v��)��X)M�<N��
�:&[`L9���S���_@r�7G���e��>�����o�R	fV�R�}�x�����5A��Ŋ�V������Y�O1cЛ7e��X����g>�}}5&O��l��b;ZV@� TJ�x��e�C����ဳX�j�U� ����@���Y$ģŷOjf���p_���9ե%�#Z��G
|�rv�Ǳ{�J$i1����2A#d��@��@|�'.�\���ɽ.��ogc<�gQ�@y�\��+Y�T� >�Q�đ��	��OqRe����J�PP��f�<7{��p�y>3�r��W��&� ������8g��:$�S��]�e����K�21��d��zє=o��+@�kŮ�������="�~�������˩\bSTڍC}W.�~��<�8��!r��)[�!�'*�8�]��]B�0�^��3>�0���u���I�����j3�(����(���z>� ���3ˡc�/j�����tLaZ,���C����g�76&�N���9���WsB�7a]�j3�jm�J���Y��UG�k�@@�����v���GL��TPўb=3rq��i#ǘ8��y<#�L<8��^�s�s���m�ԉEB�)�� ˛E���s� �o��Ҡ����t[0�#M[y��aB���H�'J����������j@/��gcC�`��հG�����OȽt�S\�l�簶��:��F��J��B��iB��ń�j��~�
A	�oF�ÿ���ꦑiy�bn��p���/z�^����Y��B)��{7E���*i����v�i,�!(��	�ۏ�h���-���+�烲�z:gJ߭�D�0[��Z�����]��-E|Q,�P���򽩬�������o��~%�����ͪ)ʋ�-������g|XY{�>�ݱ�R�#�]Ǻ1��EwF�>,L=_���M����	5QM/��G�����l�ϓ��3���2�,78�c���n��C�@�PN���Q�Ap��@s=}V�:��6��s�����#���"��3��E�c��+���#����uI�M�U��?�Z9
��O���-R���l%�aT�v6L��\~i�˕G�²��)豲�Ua���ՖPg�j(��K�P\z!��S�c����%������� �ي�z����`��|�8Д��&t�H���h�:��|Chߡ:n�!��
uss���2�s����@�u�z��m�3Ǡ���B� ��qg�L�k!���:� h�(���ڞQc�,�����ln������W)+$��fѲ��-3��<S��\�ЛH$W�q8`D%�y2�[\�����'*Œ��t�%"���v9�=��7��qỊ���m�V]:	^����u𙸄#pkb���M����U4hk����/�$P�d`��'���E�*/��@�HF~�&^��@}
:*���н����ygQ���k�VgU�5�1W5z�r�ijJ�E�G�I7@�mc`�#�5IԔ~�8hø.O^���r|L��*�u�Iȓ��7�i�;��E+e�e�H��!VZ&7��+���3'Љ�N���DO-P|�t���I�;V���]@D�t�� m�NP��c�4S�][�a�Q>r�M����X�Xz�&�S�����o+vk[m�&�D�.�i�"�a�s�� ��
ni�#�K��n�g�%��4	�W�� �ӭ��XS|����D��8��o~�t!<�19˸�q��LWn{�g�]�s�b�����.!�2�IR�"�B����Y�ep�͜Pc��7'���s�U"ck��ʵ �Q�i�L-�u�ˁ����j-��s?_iM�����2tT�9qi���U�8�?z��6���زHT����E�Z�ݪ )��������m�K_�ۅ�N�k4������3�x1�z�ru��;�Bc�6��qd�#̗B��!�(�m�i���x�L��O���C���e���ӓ�.�>>�O^��F�*��d*��tU4�]^�̚>�ڹ�+�pk�'�4A�%XSkI���	��bd��[�<�1���$Tr��%1���dR�\&���Eό����叙[��H�!��Q�3���b �ݜ�y;GX�hO꜠BG~ڲ^9.h�&y�uA�,��>K�M�<�n)�y#�MQՁ�rOh)1S�zz��2C��@⠆�(٥CulB�J4x�CZכ
����<B����rI	�Z���6����3�w�����G�w�A-Oŷ�r��o^�zs��-=��)E�Ʈ��L��<d{�9����7��51���?�	8�Y$���,?3��n�;Y&�80�
�/�Ls���c5i�_��V=�䆩��F
;N��ȁ�'e/�E���G]���\w,�L;���QEM&�eF�%Ϡ��%���L�IYx�v6jE
`o�ՊM��2�UJ,������f_�?x���LYǋ$:��R��yOCgw`(��1)C����Ã��j�Y�A/˹P�]JAxC���Jc�3�[�b�lz���M�:��:�q�F>��A�������noza�F��a���!�X�3��Xx�B�e5�M�ڕ�*]�À[˼��/ �Ġ�_��{SMQȀ��aS���11�m����T�wW�f���r����c|�;~�͛\i;
����5��e/�7Q�O�<��7M�%�V��[�Nڿs&gH�H��}�=��t��皌OD������,�XgSZz��j��n_^�9��WR�G�_)[3��`��^�L�q��o��!�%�	�3�$�@��:Wh�;��/ ��
��,i~����V$F��7�4�����g�:�0|~���]��\����^��ՙ�@Y�J��wU��-.��)���ә;+Qա"+x�8n/I����"�]%�>��)�t3��%���Og��s�����܍%�i}�drL,�K���P�5vT��6�(����vT�%�B0�q]�/��N@���O�`[fN`��թ��セ���M�]Q�����d���|�c���A��Xd�3º��bM�+���,
N��$�h-�4����{�3k���_0��?BRT��L�|����ѭ�1p��Q<�p��^U��e����s	z6�u�����2�6O���l�[w
�C
�@s[�ҟ$&Ӽ}e��3���=E��7Qb��Ui�X��BVɪ�j�X;�V��~���r�P�U��/V�OZ3c���C*kՎ)�A�r���qE�<H0L�)�� �Bx���2f_o1V�S�D��댁�V��
GWHєVlۂ�M��]ݹ=~���14��M��h	&�t�㌷����p�F��̿BL��t�7q���`�t<3�e�^����+x8k{�ll͂Y�c���T[E�>�ဟ�7y6���,�$��E�0PHϳ�o��|�_�����ƞ�ߺ�*Y��v7Ϊ�O���������7b��d(|�Ѫ! �*��<\F�l���pU���.-���h*�pM�6�͞'t+��\(�<N�	>#����S��̃��-H�P���w�p�@P������@2�b�_Ө0r�fI�I�!F��p�{�D�D�ֹڣ�i�e>��c�]�/�	���d��E��L�i��E�`�B�IT���H �Ur�A���ʬ��^���ų��H��Q�����Ǥf�pb�Ru���bpe&e�`eigH�l�Wnq�����u��殹��m���Բ�*r�m�;�C1�����yЁ��Vp?/���d��, �y]�h��)�K0���
HFPl���B�K�K��?O����ٴ�b��Y�N�ت *%+�e�c^�<;��2ѧ`�Da}�pi�ǗL�ï4wV*�W뽎`�*h�L�nǙ��(��D*)����L\D��,�g�Sw`���>�m\�ݕ�긹��`�L��H�Xu�:f��@
���M��U@�����ⷽ�ӗ�Ͷp /<e��3�ߝ�*\%"�)6��g��'�Ws߇���KԺP�	���]�<�AH ��q?�V���Rn�����+�#����F:侮Փ���ٵ`3�ͅ5ǮW;1�u��f$$e[�7�s�6�������K�l�aT+B?�I����['����[�9W���T5���w?@�@9�mcMw�~%,�j�O���H��|\���gzM+*�N����=.�ة��Ӱ���<�\~�m�Ёi��"i�g���h��=v@�9�*:D�m��_t�{�V.a#Ϊ{[SF}t֛�\؞�	iCk��r�>.��r��W���/,Nc0`��14:����C~$yw{�f�3�Zn�6S�J
�8=;�޸�2�ւ1s��+Z�o3 ���ZG�8셯�ģc�n&&�W�դ�^�VQW���C�dvUkU�یU�K�E����sG�k;´L�('wnC�o�ً|���<S�o���h� M�8^MT���������.���C��
�v���ky�-�A�l �²��R�����SU@"���k�8�"�Td��eh*�[
���Y<`�ɝ��q�B�?�o��'H9���WJ��x0ϻyr�@�m*����FOXiM�_y2�z�*��� t�ږ:�5!dX��w���~*�[Ҫ�m��1�Ե��ĮsTar����Đ�M������p����dU�$��j��T7EuGKg0����&¾S7~G��qd�AY��d}<�������է?s]�� �f�zL!�2��Ѻ�j���
�[�SV1��y���3�Ҫ�&l�@�^щ���e�^�=��1�3Cj�]&2`[<�\D,A8ױ��
|��J�ڇ���*�o�wʓ��ja0�O�����Y��!�M!��{Y}�M5ߕ�n���{#"��Z+��ډ�����Þ�H�E~���Bc^rN���E8�O�9h�o�� _\̑�����ԙ��{�������Hg}�@cX��N3.@�o�E�sv��D(�Hߛ2-���*���U����$=K̤;��g����*�9N4�+$#���A�"׶{��'�qqn	-T�O���Dvr�$��v�xNފ�a0���l���-y,�ڂԯ%��z�ѰȚ�A�`M��&���'�"�O��Z�m}3r��z
�n�P'R���@$r%F����� ֞
��8AM��jlQN&~_��GT�Pɖ����;�>��������i/Q��J�7r�a�E҈�'�"��^�:,�fV1./fm��oM�����O��W�,?ڦ����sl��5~M?c� +�<���@��B���qs��U�ݠE���zZZ��q_$U�yi�Ē���������#���M?�%uF�,fV{�n%1�K��{�"H�]Y�����NE��|�n�'A��"=bd�D)�\>H�_����'��KG��v�M#WqBگ��-���[�6��C�9�P/�Z���TRB���d7��e2;'4��d1�������W��'��𗠦�f��vQ�/r��A�l���70�v�v��}�O����G΀J�DF��5�8�Z��7j��M����9�Ȣ�M�ʁ���D�zE��U���Q���E�i�����Š�2j,2ǻo�N��2)
݈����K ��f���8�Uh�&Z>ٓ�u�]z��2<�q(��ɀ&̣v��E�^���O�t?ˡa \
��Z>#�12:�0���#�sĺHI+t,G�0�5�J��l��/�W��ߙw�ԙ�
��s�/?`���7�2*���!),��\����� �d���n��G����ЀMܶ��&'���ߩt�Ym7@]<rLiي�ba~	u�Dڌ��]v;�|�G �vT�@L�
�D�L.ߔ�&�)�z<�u��'�ϒ�3с��U٣�� ��)��,ä���/�k>1U���5{�cQ!�7������uz	5JB�,-��|.�HZU���U����.�����R����-~�����	`���'��Y��R�^o�9�Ls��������<c\�E���,�P�����T�!rd�]J����V�Hq����h��C������Ӑf/YY'��?9sn�Ef��S�G���q��mPw��s�� jX$33�}�\��^�ER�@�v�>]����T���T�C7pg�G�u�FӖ�xF��vӿ5<<��ި��vRB�Z�"�P~�z�䁃�	���,�o.T2H�>�DP��C���I:6�q���L)��⫚X�24)�t��^M	��Y��$�\��6�a�+�DޜfOGJ�&�=p&~�����Gn���r^�$�Ɏ���t@핷n;�9w���{�S�Q�Ŕ+���U`��u�����b��$�U,��\36�&B'|��0c`�N� � 6a��ߩ�������y&䕏Z�QP� ��Z��7�F��&�h孬�:�T7���-N�Cq�n7�|�"��u��q�c5р">�׸}`'i^�*U��$E]�7�1H¸²��A����3��-���k�Rŧ���x�N3g�ݤ�/����l��蹂�� [|q�.���!��:H&_�-��]��Y9�cL;�� �ۈ��h��r-��U�ܶ��\�K������8�O���s��goQ��w�,;�ss|Y>�a@�a��Ź�]�&���:����#�+b�S�����f�z�����	E��b ���Mw�{3�̈́�c9�Kp~�%�9E(���v}�O�yC�@�Fl����z�qL�$��������?�+�N��� ���%�W�E`�k.�E�^����6�jf�u�%vu'�Ot-�'�(��<{���qd��+���x��cJ���0�1cQgL�"�Uϡ7��ߢ*�¨z��!d�^4{܄�@�jrM��[���"6}�N0�p/tQm�\&������04�h��
8��@�e�p�4X��9&�>[�^�c��ѐ1���,�����~��
dK�ph�H����J�~<���chn������S�Vf��V\iw��xVu��,*�3���8��Y����e�l��>�q�/���Bȧ'.�J���#{��^RvO��Q+�(�!�ڰo@��D9�ע�|�gʔ�`�q��J�����5_`���Ez�@��������ݪ�%@b��t���΀����%�Z�(~�����f� �$|{�7am���[��=����7�
�Аy�؜�u��tƨ��f�;*�izC$�	.�H�<�o�r��.Y���RI�(���z�J�m%R�'���@	/&�@��������ub~F�4ˑ�Î�N!)M��1��G&̵�*�/s�Wl���v�㙎�G����i�m��kUk8��������
�h�cA�-Xd��@My� kk�B?�Z��n�ɯ�X�r�٣�)O�X��X�����V6��w[ꙑ:(���=�ғTׅq����\q��]D�`�]�f�p}�<R�oE#e�#׀��F%*����mUw[�����,��^����8a{�����>�c�-UxMڇP(����#���a�}?|��Z?��I�K�k�Z0�H�J�����V@�(�=V�X�h�= ��x��Y�7�?�}�@Anz�jiV����("� D9zb�u�4OO6�H��?��%�$��Lx�w񓸆�zy�n��=����Ǉ;��'��G���vf��C�r�A��2�O>?��On-��%(Z#����c�	6*Nf(d.1�[l0��I՞y�@ř��]��N��-@�̽�<R�/�5�`,8P�ǥ6��ۈfp��#�ljv��F�D����F�*hY�xk~4q�\Cd�j��=cҴٹ$[N�P��ҕ5nb���`Q��i���5۵oy�h��tr���{�TQ��5(���C6�K%��_��e��&(7n-��(1Ȱ�T�B�Ԅr��CcV���4 Ja��x�&D���_;혮d��ΐv"�P�
="�M�P挿�N��K�ȅ w}�m(�w���_�b��lԃ� �Uٝ@n�;RG�1:���< ��OL�v��=�H4C�I�j����+ö=b7}����6�ڪ�܀�%(�뎭�{��޿!�;/�Gz*�����.j�S;��e5D�_��,J2��Ö��߯j	2n�x	i��,��2��d���_1H��6w�g;���S��x�r(%��h�?&mp�	�:Bg0�� j���F|�#�B�<��Xw�z�XUQ��SՑ��Y.)�8���H��ٯ�z%�S����	�HǢM	�2J}]�#a3DnȘf/3�6�O�A�q%�9p��h���r�����ޑ5����8��oXn5�St,i^X��๻���ڀ�q1M�0��
|)�/���߆��|R#�����O��j�`x�U�v +N\�I���Wy)�HI�3;�FEP�|�e�H��.��!���5�E�L��UY<���((=�h̠���$�`d�wq]��zV���ۓ#V0o?�ڸ�J��0�'��tΏ����o14k�&�t!,��PY�4�M�m������b0���%��yW� �N!��l8ekt�h�cUM��\���
��4��#α3O���L�{��C�MeG��$/UU#���v����ez���Hk�kx������^/�y�K����rgP"�*�U2x!Kk,�/��hR�# j��z�|U�r�c7��L8����!�	�6�*��%&P�;ҷ/�7��|���� ��kJ[�ZJd%%BW �wH�xL?�\|Z��F�g k��S��<�-�m�������aY�ll,lqYD�h����C�����Eg\��I��x� ��ټ��B4���,]� '�z�����D%�uTL6f��,"�ZqnՀptz��P��h��t��pWiS�lPҥLǘ�R�Ċ��M����A[�q��D��]d	��,���ߵ��M�2E�y�0P��s�t���4��eE`2�A��ȫ)W1�\B��J_�E���ʐ�Z�,�W�b�Q�9]�@C�q�B�z�Q�ߵ�7&�M�6����&!�I � ���D[�q�b�۶.H��?��b�23��i��9�b�̸/by���1"}���Lk��t������P��qt!�guS�.�u)VHzȹ�����ǹ��`/��}U���J��.�g!�F;I�Ķ��o3�z�����<y�G\�j"F�Nɢ�b�-I���w3If�*�����"����j�z��`��@��x)�MB�F�s"ӭ�#�0b*�O6�w��:v�_����Eu��\��-�,�Pk��.!������?�N��t�����1�4����O7r������( �m�����ޠ��>6�ݒh6�B��x��v��g�i�ߙ����a=V���ύv�Ї�s��"1�x.))~���:�t_d�T�����S������"`�F-K/\ػ���W����r���h0�-r��X�d����|����s�&��<�Õ��bn~zkc9�|.s�����ڢ)�ML\�%�lLz����;#�E��)R�~0��P��&$���Ad��?����Kaɑb�O�����G�`�%� ]�x@�=Wit��f�u��#A�3
����[� �M^���t�Ԃ��2og<�)�|��9��̢� +Y\V?�y�����+��3zc�McDґ#;!�F��!�PT�c�ߚ���D�ͷ1� �P1���'�q��Q�Y��#9�/T����c,P������>�
	!tM�!�R����󜙒�W����	���#iD��}B(�`b��_h�9W<�w��Y5p\tZחH��My�Z���6[�eu��Q�����-��/��M`}�Ř>�\�1K\`Z��������܊`��D�
���rNV�Vd�L�*]B�l�L��5.2ܙ���mM%�Tq)G	c�&kB=?3%�wΆ��&�h��R���~beL��$��p9����0�Wym��f=XP!j��_����5;EA��?��#�\Bpv]O��-�����(yb���ԙ��: �5���y:R�D#p��4�t$\���1�c#��q}� `%a�r��֡�.kyC�R/�)���n`�����z���ު���r2aH��[��H»DG2�F���������M����CF�%��/׿�#��E=�@V۝6'���3�;pu8�+3���WV;M&\3��QG�v�MS��Mh�M�,=E���S�c���Y��ffj�K| � �z[�o`��`��p
�m��]�E�,b�#c�� &(�����󖙡�����ե��%O@���-ҿ|C��j��S,��4�wY��b��OG@ ���1h��Pm�P>נ�����M+�gE��`�+L�o��?"s=���[�ĢE�S5
9�u{4��a�C��b{��k?��PV��,�AH�wW��2e��9iMz�{P"c@�Q�be8�t��>b�pί���$���&�<6����X	#L?�!��y.�q�N��UPJf'�9s��^�Y���`9�����.��}�?k 8�Y��7�h��e<�VXcaӳ�V"��ƜܑE��h�<����N ��At�v�	v�J��Dh�0���\��	XG�U��m����TeQod3��iJ�8�;��&Y&u��� �
A��";M�C��D`ʷ�E��YR�[,$M̥��y��PP�/�{��M�^L��e�U[�2nW������2dU����y�*߮�����t�,	LLK�a����톁�8��z��黰(�#�2�eM�L�ŋlوچ
�E���+�z�xoEU�˗]VLL�$�2F���P�G �!�m�ԕ�1��9&��}Ǆ���6�+�ư�ʖh5�O�;�d� �m�zD�tau^����|�0|G�j~y�&\��l�o˜atQl����z�|w�iI�l�hh{U��^��h3�[Z8Ɛ�ۿ�e��A*�����Ն�9����Q����N�P�hs��6_���`b�шN���>��W�8�,TeM3�;CTBٟoK���U�׽>�Qnō�X��X���B�g;lL���孺5��>e�&Wo�� �m���q�!�Є7�=���b�m���k�3p"E��^j�>�Y*~�{��cK�s�.��Ca�]3����9�I��1�X��� �>o����L$a�[�t<HW7��>��z��6|���RZJ��#�n��8��|��h�a�{_�B��ö�(������d�{Y#��(k8�Z
�X��h�̹8=��W?4U�A^�{�Y�!&��	�i(o�ᐸ ��[u���%��Q:��Q�>���W�f�K̕en�++���+�Q��-��YS,���{�X���\:���bG4�!��o�vR1s6� 	Z�B�P�ú�]�P�0��$��m��^1hxG���ߗ�+�ŊL�D{��&��4 _�f4R�]Gx�uxC�۫��Ru(;wU�������<�;7�K��q��3���C�2�|&6H|5��d��������C�U�6������Edy�fV�>��c�����VpB6C8�AB7G�ӹ�|'�}�H'g�$P��ЪO"��L%�o���*�k�8o���v'��lTH~5�_��w�{�ͣ	$�\U��f��O�Ŝ>�i�;��$�H#�OU��+_��+;�{��Ѳ�~P���sOd��f�ձ�L��b�ݷbcDh꨷B<�Z@��3�'�G��_Ʋֳ��l�YrIxvmv�G�3*�� +}���\~����!�5Bג?��X
�J�M��`��BЭ_FoI8r�L_�湛���7m��L6ps�pi�����
�ѳxק����r�З�Nf��)1�ݕI!	��p��t��E���7�d ܯm��Ua�m\D�I@3)�͸P����ƪ,�����h�x3���UКC4��È�"�E�	B�K�\BI�ܲ�y�'x���+6ېJ볶������c_Q֪(� ���7�� lǛ���QȘ�l�,41�j�F�adKo�nG$�$��:��0IZ��'��>����DȰ��{��$�˱}&�ph�1Ni�D���-�=�������d�L3J^(:*���-G�+##�Bio�;��B3�3	s��2lJ�,�\�3]��AA\�n��d:���w��G.��c_����Bٲ���%��Tk)m'����3A7������hY<B�l_�:�"'��U�w����v��lZ�d�*e$*��$���2�Ff�jjf|���!�a��"�jy�Tb�
��a�11��E&0]�L���4{ڵ�;x�C�>�ca��g��o4�_A!R�M)[,�p�( �*�"*Ƕ5i�Y<dRK��qXԋ9~_�R�4Р��F��#+h��� �/1�8`]8B��;��7��nl���
,Eo�񨰞��D]8L-O�rP~�<[hz�v��X����`r�Bk������z�����P���Y�òؙdO�c�E5���^f�*�.�(Db8��ȢVd�ٵ�T�����P4��<MZ��Xi���
K�3�D�\�A��9�T,
��Z��}U�|"ˉ�)�@ �-��;�p�9,��u5ܕ����3mC0h��Q�h�2)<���=V���0�3�	?Fi�g���Ε���b0���=�Gi�4��Wt7ٻ��ͯ�ͧ~2sH�`�ٵ5u�S8�/m2W���'��t8D
x;w��� U����(I�#5z��G{���1���Z�@�}2kYtA�e}U�mtO;-ȟQU���(�h&v@��Md��q�C)RA@+9��z�8w�T<�p���Ȟ���r��8E��]��-�����x�P�B4�%�r�{F�h�3�b���x���Z}��~���{����bm����ͮ�|~�A��uwH ۢ�0��s�>lu�ֺ��A~dE�I4�b�rO>�mKʼD�Ѡc��[V��,p=Տ&W�E�{h�;�|t��"^�<�<F��\2��A�y�^��1���<�Xf�,���o|�ނ���'s�k�"W�QUg��?�~���P���Q ������]�-��vd�&N6������h.z3ؗ�"Se�PA�`nv���3M��� 	��!�Ё�*�9H����nZ.�HI�v�2�)v��y�XHC�1L�a�J�Z�1Y�
�hF�I�>���r��V��WE;��3l"�[�����߄'9�l<!FO���T��k�D8�;����I��_����i@�s?�^�����V��V��3s;�-��r``�步��w��0��AE2��u�:yh�]�,O�h:A%��PB!Rri��H�N��A!���:f�Cp[��?Q#@͝OH�u�0�Q��N�f֢�$Z)h�G����TyZ*����a�ppR	��,�zQ�b�=����w������qǤK�	c�[��|܍ &,�7�d�����]��=�+�=�a��\��f@�B�~�R�j��s�&�2���f�^}E9��]�,%s6.��و�7�
��1�/]m��#�.�������A�m-n��j�N�!S�8v���W�oN�m�9L�� �:sqΥ����b�-����&��a���n�tQ^{�`���_=~��Y\�ʳ�@eG���H9q��v޺B�L�a z���dm?�� N�3R�^��AM�P�5W�^B��:b��R�ktu(�Mi�/(,ؓ*V<̚5훂���v�SԤd���L�!��.	���.�NT�˸/�X����� ��K���A��9�`2繆���?�)Hk�+g���o/�	\FU�rj��	 �m:��J��ھ�ٻt*�<	����(�ˤ�zgs{R�!$�:��Dw��=�7�<C�lY��_ N�6)�fU�qj�T�}����D���	$cv��!1a�a�.(�Xɮr��k�����`�s�@	��ڸv�r�fm_���aD��r�;��,߼��k�ii��GC�H=Wi[=����t~S�'��^��6��f=�otnNb��h��',��E����g�@1�J#��qH��W����c7p�tU��G��qw_�
 �����j�%�ɶ&!jþo�Kp�ׂ��u�½�2�}�ŉ��<���T5��GT���v�w��7�S�uϤx�ҵ�xj�(>}�]�r]�9	��u�q,�6�������fM�E@��#��0�d7tdd�(佡������L��de�D18E�3�7�LϺ8:ħ����'�F��}��!~����0��6ж�`������M��1���� Ch�ʇ+�j�V7���|���c���G/+�y��ė�b�9:�>9�-�~����	la'p�S�y��Z��g<9g#�eq-
"�Z��Y7�4ٛ��<��M��|�L>[��♭ ��8��1��kg���m����JN�\o"y����n��U�ښWL�������ǫ|�4�������*
�WԊ�9�E�g�gef�_�~iH�0��_d�SdnA䖄9�C-���җZ�h��+B��ߪ��*7�#��A�Am隼F&;����?�_���_�&��A�pL8�B�z#L��~����-�!�o��?E�K���_4��ˌsQ�ѱc0!��LEm����5 T+�8t��Ş�vَ���X(9�LJ���5C���䉓֍����AT}�7,M?w]!.��g�mr���B�0�,��Hzd��8N���AH�����_>������̉k�5r��/�I�t+iǧ0�i��H_��Z��r�o]]� ՟�T!qH��9�2���xK��w�٤N*�M1��2aK����꾿�ܑ�9um(C���}YN�fn�u<�K�����h�Sqȣ�Pغ�]j%���ŅxUHG���c�z
6��S�����
��@[��Wc�F��/�I0T����"u����	��V��h�.�.�I(n�K1]ϻ�_�9�-w����ǡߣ���m�@嘐�`<q���W����$H�������t���f�BQ= J�ɽ�I,�TpZ�GWN̤�mͰ��b�W^r��>C�ڨ
21����ޔ��^o�;J�64`γ�O2�Yc���e��?p��P�A��')������&�XI����?��`����
��+ �Й+���k��>|��>���e�簾XFKjTgܧ�{^�@�;�b@#���y����ԁ:���wE�QȎ�ِ
���z1�H ��}��m��{�s��؏�g�!c��3v&����NU;��(%�p9�밀��C0��N���[N߅t�Q��5]�}\�G����.�K��������ת:�r�B�3A:��8��Y�L"s��Nr�0���善z�@ه�>�'�H�t�A=�Jx8�@��F9�լi�)��W2=�>T��{l���"�S@{�/z*;�'R�7��ϴ�F¼32���zcO�f�R3���޹IH�t]��ߴ�0����E�&K[�#�5���;��D�I&�w&�"��4��+[�w��
���:T��eM2
�+HŠ���8D�au�op�kTU*L�liً}:@Ʈ��ٿ_)��iJc?�l4@y9(��}+,?����$5�g����M[W 7�խ���a���mi_�D~ס;�!�
vo��Ƅ�_�:i�P.���N����oBK�����>��uPiK�b�p����<F��Ө����G�	`�~į��M��'�?8�m��x�Xy#��|$}� �)x�q"� ������D�8�
�؜Bnh���Gm'���R>��?�;][?;7������rA���!ټ��UE2ݥ�m ?D�n�h9��:��w�c5���H��%��d��n�S���䩻�T<�dy��B1�,���/��h��1W8$U�����ǭ�@Dti=��{�wpP2Z���F��'���%����YRڌ5E�yV���~>��$8H�����ѥ�d8Q;��\0��W��Kh;�/�H�6�;�>���{[���
;>�[0������@���f����x7�I�F������q��1�JG �t����1����$�U���g�@.�]�?N��z$;S��X�<*�����:jF�쏳և��gx������O���m��"n��8��)���ʪ��UM�z�Ɋ�}*-��Z�J^ݓHtN7��P�/�������'JE��N2��@�
N۾�V�u���ya��X�3�``&�C�!� ����g��t��}���LJ��1���^��S�,���ć�d! #.����bv�����5�w۩�D7�"Nu-���П��~�@r�JN+�z��@ѓFz���g��!�KD�w�2<��4$�Ei�Q`3��ӵu���*F���E�F����m���S���\��%,Ԗ'�b��uIQ訬��_��2��?{��F�����*�����1ٿ&����}=���g$���EBK����OX�w��|B����m�����Q1����V���Q��ǥ�{�0l���C�����K
Y�~k�!���	}��ʡ���ϴI)�pB���7z>���Y��z�$�<�����2d]��b�q��ܸ!�*F��Dˁl=pcG�J��٦Ozf�N���[�ey�O,.�ww nޏWmn�E`�-���y�d� )OE�{�t�	��Zs�TV3̘���#,�±B1p� ���4�[�6H��Yq˸o|IS�P�>�3��b��jt�=וT�g�灉�4F�?�B@@����6d��*f�4?< �.��S���Ľ���058'�K�&l��U(�� n��>���G�P�T�r,�aK3�$|_��D	z���Pn$�u� �WD;O�6+�)�T� Y��{ĚBMk���/���3"wE��|��@8~O�
H,��7�F�Z�#ha;��DnͲ~�	s롥�����i�$��J�����-6!�B�EL|��P�u@~�b��fl�ُM��%��g��̠���Vv�\Mt�a4�[��DT2(#2�62ٗ�G3���#�#�������Q�or����dU/o�Ւ�j�[։[Km5z���IW�#A��β���}'��	����w��PPݫ���
��F�Kh�*L�\��Y%qM�$�ֆ�<2ת� �����#��M?�@��W����^�;��q?�Ԍ�vͪ5�.w�fɳ�3r҃t��d���$�����
ڑW�Lmdw�:˜U˦4T`U<�(GP�����8I-cdR������6��#���aW�҉[ �m����d��j����+Қk_�3�}�yÃ�+J�S��H�������-�
���d���h)��i�$���`���<����Ӥ|��	����q��V_�Zk� w��~%�+%�X�$Mc�S�I�'z��7 rع΅�]� t�UX�?Dؖ�ql螝OK�J�zQ�v����gT��XgN�"UL_�H��#SM��5ׂIq��`���e��
:�YQ@���#��ϧ��{)��8p�g�qB�J�J6�ӿ�FD!�U��u*���ӟ��!�d枺C�n��[����C�4�Y�� A����?�}��]�������yNw����a���'2{��������QDG�'j���0���j�N�G�|���C����L�<p�G��+��oT�񙢎{-S+�M���+���%Z����i5q���f�7�:ygوx�m���4���0T�0an}���D��@N�$l@���y�Vp�� �.��h,"&S*O<�T!_\���J�3���tU8�eW ؔᄱ]6�|�$��Wi�i
n����?B�r++C�"�c&Ƅֈ�i�O E����w�Ǳ3mZ�up~��j�|�r�W �1�%ݥ��-LV�K����#��aZ��`R��r`�0�\�Ҡ�EJ� ��v:[�>�,��Tf�����WK��G��%��Y��l�9�SZ��掵w�Ͻ�o��3�C��O@ -Müڕ�o���m�4/��������<S�O+bj�$G5<�_$�Ć��@�ENPm?�a�,�.�j����2��ƽ��s!��3c/�O��]�p�Xs/�Ճw�e���n?��|g5�	�����'H!3ۡvxĭY������ɳ.�~�+;'��n��U�������4d��=��V�#��.CR=)���P��c0�N�YY�Cu����f���Aƶ���7pn���k]��D�~Bb�cf�s$�j�}@��̽���j\u
���LE�˗�<bt��!n��[AL�s�o(��5�̤�=Uw���3�{*�F[�En��1�k8�K����=�c�lL�X�F������l���{���Hy3'`�L���q5�gi��5�֕`�a��ꇒ�vI՞�ݹ�H��2I��l{l\��U����������n1ѭCѳ���n�߃��S#�d�;����awJ���m��;�(B<�v�������*߯D�0� 6�&$whv����Xi�U�D�w��"�ϱ�JF� �j'�[X,HG��U!ٺn���q"H?�3pAY�΢�(��� �4Q3Ң�����^	��G�!W�~H��T��{��K�@���}%��#~$�� ��LEYcU^��OY=E�Ɉ!$~���J�����^V~C��r�:��R8v�de�4��h*X�T����k	$��x�q 5Gg��e�<�cf��x�K̈́���9�nC��޾)��%ק4&������9�6�1�~j@p�a;�w��$�!��eWf�J�:^�W��n�1�領�!��ڃ�pݨ����6;ڍ�cb�*�Վeə�4i��D��9�I5��K��j���P��$���2��YF.`��AF���:��`��UlON��	6�����KVJ"�9���fEt���ynH��ykL���g9��b���&�Z�ڛh�KMe�pcC[Ϛ+�Y��{�Ӳ�3��5�3J>��������^�����4S�xoU�,�(S�9wӳo�L9��eƥ���^�*��R�v����UAħ�/����8���Wh��Y����~���Їޏ��9g]1	0��)�y<�r%"�P]N�k�ޣ%�w�F�9����
Zϕ$pB]�b�ږR"�)tC�:���z;H�)�P����9�u����z���VD�&��:o�7c�F'�e��|�B�c�_�׮�Y��#:���m!s�?���&Ǡq���K{6A�a�)	R-���	X��>�bY]���ښ�<�t��5퉷�ϫfO�9rw"k�-��i��ŕ��C���t4��N�F7%�e�@�s&l*�cW�c���P7�ӹ+&k�	�!�U�f��|���"X�4�yS�d*����v���2,J��M@�X6�pSa��ls(7����Rv�"\��|R�,�4�"��6<	�����S�ٵ��cZd��ς��gw�q~�pD�B�)���cY��c5��㆐5�����=v�LX�zN�k�..�ũ�+\����~�)�$������v�4��}v�1�ܓ{�R��4+���s�k�g��1��'�
cMQ��i<	x����aנ����C>$JG�&oXvsF2����e����Ԛ�o1��Ц�4�����Q=��\E��^�0A� D��wT6ʈ _���+O5\@��@Y 
�A{Ƹ��c����q�%��6Dͤd�_b���0h�oH�E���Oy���V�	?Ҽ8�7=������%��7Kq�/��^��z�.�i��i|#Ȯy�������`�� �gzd�n��K�ɕ)bW�E �1K�F�>�is�ƭ�!u��F$�SšV����9������o�%a��3m��[�3��&~�ӝƱE-��̄ҹq���,=�L!^�Md���V$+��E7�g�ޯ���l=I!��G6��[Qp�bb
�\���YK��|v'������VG��l�jz���J1C\,/�� β����٢c�E5u�1͊�+�5=g��k�<��*z$��P�>{r ol�7KX1��ټ'0�_bk���/��ag� -��ɲ)FZ�8i<��;I�6J
Z
9��O�^�|����ގ�zW��I�(yp�j$�8���P^%x�-x��� 3�H�&�5A�W��F�`��-К���ag҅-;Tpb�Uh����H�����c���	@�W� �<�乪L��1��s�gqb3'�`�C۔��c��<�z�q�F�d"��%I��|F�|d����r��E����vw�qP��3G�Z����I�%�*�Z+�MYe)@>�i���T�$I
��|,��m�0=�����d�KD�H�Y���"�N������!$��<�N{y��)����w�-�J�d��~R��@�8�����8�K:�7��c��
UЩ�U��_b��j�zA��j���6Tp��/g+D	%`p��S��Z]�.��2��@�|gD�}c4A/���I�L����hG�~�Iս�5+���2�ߴ)J%���$\��)!5|�L���X@��YX1���笾x�n�!��	+�����,έ&Ա�.j�ߠ��^�*i�Ꜩc{�4�w`��*ַR"Lj8��'\פ}�E9{�������4*J�ד��w�0,k5���(暗փy�j;�yJ=ڼ�Y�8ώ�̺��ܝ��b���ٖé�p�`t��ڰ��Uh��x�F=:q�܀��`<����1��6�_��Zf�*�����5~����R��S�i������1 ��W"���2��b�:h�4޴	�n�	�I�����)�q#�<W��Pk[��~�	�øۻ�Ko K���]Y�z�(!�/�������3�H� A�	�P������/x���w2�G<�AE�0x�y�F��:�P�&���i�9w�r/[�|c�Y07pȤW��i9O|1;e^���*5��6�3{G��v"{W�&Hk[��o	n�zY��5����g����H��0�ΐ�	��ϝ�?u(�!��W�.��b�>?;�|v��á�Z!AmH�:��{�����Z�6�%�4|���*Ӎ���^�|TCN�')$�_��S��E7I4� 4����U�f|:Ta(z8gM_;ȿ�r����jj������/��Qvҽ˟�5˯n��p (��{��$B�D~����R�D�~�B&q��/���-�4;*��A��*M{�������\�J�{_onO��UԖ	_�O�9�xU�0�8�>�F����ή6z����X$�'�Hc�;R�✗&�����l�r)��ĕL����̜���A_V�StY*-�$
������,C^Eʓ��������,͖�G}�@�~�T9$��n�h.⌌�U�!��¤Ƣ�E��(��7ը�?y�g䯀���w���،]��}0��l�](W�s`K��{�W'RM�ZL�7��G�=�'ٿ=L��rQn�L�m������Z�*/�-����
}'��rǴx�*��-�����W��-Pӈ1�جTג^rc�b����V�蓧��)NVB*Y>
�>�Fʺ4wEћ�����R�r�k��7�L2wvCՒ�Bl){Z�4@Q!ϣ�Sr&4:����\N����[Kyq�2�<.���:�u.�,t0e��k�a������r8M'x�NC7Q)���k$��5�{EM_��~*=����b�hs���{�[q=�<�� �S�϶��Q�Y;�||o�#mP��7�0�T*	�kш�Zx	C��
1�7P���3��$���t��% �ƹ~Eju$���k�	6�0.L�^���c��_���a�G�&�I��0�vF�tX�,�{D_sO�X���d�^��ja�]��Zv����F��
�kCI�g3�̑���x1`O���U4?'�t�*�JOY�iCA�M:�]�kƺ�T"B��z%�-���e�������U̇k�,�T���h�̌$��*}uu�O��?^���T�뽉�=�d����Z���)���}K_�����sM6�Ge@�נZ��l�dU��ކ��o�6M�"���fW���EF�xW�D|vvm��N�J�1oWoZ��YWQ�t�F?c;?-b��8�.�0@�U�׭^�K*6�`�"��x�9����J�r��/4݅\!�rH�\�\+�����!���Kh� �����o�i��pu6[0(Mk`͝4��uq_]r��EKS��ֆ��I�P��.�*��
����%�ϧ\����ʾ�����:��*�ʦJ�!��j�濱>>>ٷK�$����o�
c���z��u�E+�?N ^ۉxz�x�|{<7� �d�ܱ����5���-}e������(u���b��V)ܜ�(�FJ�E����Iu|5b=�?u�6X����Z�U����RY?Xf)aN�I�8���Y��<�����3G�jZ��*E�K0�D.���ݞ>)2�bLM�}�8�t^��eG-s䭷�QjW��{��'���ś�@��KX�&6m/be@z'���guh}_�{;����.�
�H�m{-�B�50��������+5���(��V�i���F������t!�#�~ʆ�h��-mɬ�X��(�#�27�S��G���d���;�G"老3�ti�2Xc�����}gEKr�����:Wp�b'# ٠�d��#7��r�m��G�� ��D�� ���1Pݶ���X�Xy�୿���o�����o�Pt�Ҥ�2g\�!� ��E�?3=H��:�n�Q{v�S��t�j�$�{t�!}sM6�]�ל�Пy��W�@(���?t���w
F�qPQ�[���^ޚ��K@T�H��� XK,*B�	���tˮ�S���o�POA�0y�����e��V��S�u��>��޹7�K[�م�(��kAlnC�f7ĝ߲� ���*#p6��_����K:��L!�!�q�^9��a#���~A�(�-0dta����;L9V�Q?81:�I���jA �s�/�,�.*n�/;�B�#��/}�x�����Q�QS���OXqE�M�"�x�$ĵZU�J0��J�"�GF��
��8B��tO˨�\G�GӐ���PY_!/��5���X��xd��\�>���h:�d5��9H����{� ;�K�uI �%́���Ȑz��ʧfF���%΂T��1���{YN�)��G#�ZW;�|_v��.�r�>D˘����11��jc�KFHlw��"g+��8hwd�{ b4�
���Nu;��
y1�N�V�5��������,��4oƈw;t	�=@W@��hkL8��ֿGp��A�Qb��u�P#�� q��E�q�?@%�U%d ���D�k_�#׳�^�?�d�����h(ɩ�/��
t�M|C�ɯ!OW�,�u��w�c��P�t�`'D�#�I��%6\�/]+sҾuhT|��?�R� �Hs�o�3H�Q�B7|�+��p�d[���(XF���[�c��/1���֔n�jо�� ��y���b<��W��#�6Z ���ϼ���dy`]�B�+�@:��k��(�����6/�1�+MH�x�%�xg##��/�>rg��E%2��t:���۠ۘ�U�7 LЊ�N�������V�&����I[΂�s u( �-)��8~I��l�(WQ�wV F�W��M�R�u�Qy���4Ҙ�:"��0w@�Lc{�'i�I#:S�9)����e�%ܵ�U��8
7��󌲴&�36�f7XavE�KS	<�Vj�ǐ��R����<C?�9
��-A&��I)�+�]�S_W)W����ݝV� ��pq���U�<x��#M�ߴ�|�n�ޟi�	��������/�����nङ�V��u��>.�M�����r@\�5r��kǱ!�l:嵍���K��i\�o|���eA':~P5]ԩE���O>,�m�|���K�rH��W�^����D��_y�%����n����g�w������Ra�]
O��a���ݚm��>,f�����,	���Z��<c٘��'ڥ�1l&�oW�K-3M�BW����$�4#�h�UK��Љ���>Ƴ.�:�Y��[JEq�~��f@k;�,�ܮ|��M�*^7���Z�R�	/�(�����F�T��x{��S�b Fy������	_a�,q��� �aĢ�:bwV�����!_r���~�	2er#~��i��e8e�FC�&M�J�Y�[1#�S� UuH"�]�F��o�H�=����4)%ȘX����� #���*VE@@��_'ҟ[����lI�����\i�s@�e�XU�q�OcA"-]���~P�b�pc@������nH��� 5xҐ��׾���V5� A�V�&��Iw��%��}��/X�Kи�i�P����l��M� �f��͢hGo�ɇ?E�������;Y=����#)��oU���2�^32��߮B��>��Y�莀Br|_�o�&�����ኻ��+�T�(z��
l������b�>8������a*v넞�D*]�j����<���Mu�{*<k���7JQ�A9`{�J���;B3�O��)�n B1^��8�=.G,��1�����*/N/n��&�<_(r�,��8�d�����Ǩ��X�0���h�/�to̤�ظ�*�ܲw�m��$�������@+��~@\!��Uv4��w�$R�j�[C��x�6��uk|op�ln��jfwD�i1>�Tؔ���Yn��>����r��t1G���Xb�/����j��Zz�ʯ@�>������ibW&wC����1��EW�}���-a8���)>p���*ЏU[:��4d�r05j��\T�n�Ѷe��f#������Ct�o�B4����X��R�b�ū�U�vmA���F�*�Č�
+T�X;��Ӛ�*�j�X�,H�_�h�^(�V�׮N�n$IȆ���:>R���hc��6��V��16�� */��	�,�� Qb��h�w�ĉI���g�4}�PC����_(����"����}�"���җ:����m��Xί�.������	NPM�S����y?D]"���x7����	״����bY�y���( ��O#$G��PZ/&1ʑ����5����%�c'k���ɹ��?V{����=�T��V9��U�<z<6�o'v�b�,���`�S��~�$��F���r�)���*��ڏ��!��r�\��ᔄ<����BH�֨X*���:�@�spB�Y��vA�+4 �K�8�������%�#����6N�#��>�.t���꼙����Pr1<uT���	@�
;*�R�f�\ǫ���B�\ʺ�/'%n�!bILnl���a�Q�I$��ֳ�	J�T���fcDPݍg�w�Wq�r��Eʆ
%me1���7�/�?���#$��ؖ�DX�'�>MS�Օ��Y��y�,O9Q��#~)��@�v�<z��-�.0ZE��ybR�Ǆ�X���{��*� �O
���\������V�|�{�k7���R]~���DЯó$��w�|�_"t��Ybə���=��30�>�G�� �1�gA��5��C�[�A��7�T�TҒ��\�Fc/I#h��\�~�Pjج���Mf�׌x<^{9A�U�f���p���)\�IOY�D��%Gv�1�G%��Ϝ�M��_b}�H��+HD�h��b���پ�s��k�w�e��z�2��I8(�lo�U}�,x�l�g�h���O�i�?��q-͌J�'x�ܱ:	(O�KHt]x�B���J�g�oۉ*1�j�*<��3'�#Z6�R\Kl�1��k��w�=�8?˅��rtc��eY�j�	�a�x���0`(��yM����e���	�q��6��x{P��Sf��������CI�ɝ�q���:�o_=�]���喵c-)q�^�6(�9��Q��� W��B����,P�7�ӷ&���Κ�Y��c�χ�,/�e�J�
��y�9�qͥ̔hvOy?D�a��^��D��������1[������G�P�w+3�)��� K$2by�RM�d}ik��k�2hU��;��wl/�	MZ�?3������Sή�@�l��a���o�v͟:>���>[��V�䚊�H̦���ӹNN����Hz��}��[�@,��xe1��ԗ&�s�0k�������P�.|R�jz����+w㊛���D���/f0�Υ!���@A�oD.�����0P�oa7O0ʬ�)k����!���_	!UѰ�>��i�^�	��ЊY=�'��S���5,u"Fj�@%�f|
p�J}X!8�{��6�_}-����>T! Y����L$�2� �*\��'��P��©�⮀3���G������Z4��T��T ��fa�zG�oWQ��� @�7������s�H�P��N�w��1]E@Nn�.�������^��G�B�:�ю�cb��������ɠCr���.��%�w�l��$���u+ł�G/ߣ\/W�ph��˶�W�]֎��?@&>L�N�k�������j�[��p19�4G��Seq�g}�!<2��I-E�@�C��v���*
EqL����Jxh��W��b�܄��3[�-~�P�,�Qd��g�}_���!�5E%�Z�%��5v՛Q_j�J �1��f��heyNp�>C����ܞ�j9���07	Ԇ�1�UB�=��/?c���5YO���l�oc(<�&�����4S�e����%MS���t���=s�M�^Dȼ7n�P2]o0�7�SY{�͉ �,}_2��ֈ#���6i��or�2z�5!���G#>˥f���үuͺ5!�5�.��B{��wR���U����9n�K����T��8؋C����njp��]$M�b)��}��J��������nQ'� �@76AH�}u4�\Z����PMH��_�x�%�{�2T	�Q��A�����I�3<>k�T��!bkQ��c%BlM<��p�P�W�Պ��i7g�����knD��@���M}d��N��9��O�oV�}�b�`̽�3�Nsrf�����z�%0X�uu>���οa��u>�Ͳs�\Z&��7-��uh\�c>R������h,�ڼ��@���!*�
ӗ�d��{��c��*E�f�.��X<��e���xi�*�Whܫ����,�|��T"�f���mXX(qxD�{X�Oٯ&I@ޒv������Sr�ͣTt��0��ev<S��Aq�q��0�V��@�C���׏�T_,�.�ƀ�X��j#��k�ί�B_�R��oxʶ3���ʹ8�Bˀ� ��k(Xo�����|ś:�^���	�*��h�e��b6u��Gy�⩂t�q����47a�&�җ���������U�4��J�g���L����`+3	����ٵG�n��tPq�]{zg�
�bM�lj_�7��'�M*�f<^�[fLݙn�|�򦷩c��`�I{�Q}��07�z� F�M4}�v�,ݧ��Y� �R�9i����G��(�N��o�����&�+�&�w��k�<�̡��8іr�'��������?U����Q�1\���#�
���ѩ[ �=�^����׭%��İ&�����H���A]ERr�pӂ�;W�x�O#d��{DZ23k���)�e�mp.C�����-���1V6T�&u ��M�	EE҈��X]�c�P�j5���H�P����˟�*��R׺�H桳_�f�e��͐CGv�+d�v�G�|���@��Ũ�m�	��ꁅư ��F��	YB�]�j�]�H�"�?��Ҹ���I�:� /(�C5����Ek�:��>���X���A�G^�8:]c�684De6�s��4f���zi�!���ĕfo�貼��
�<���ci���L�a��#�X�*H�/r�*��1���k�6��\K,g��E2��;O�(pЏ	���?1�4R��?
b�|�n�y�ј�x��z��G��/��it����ֵ��6�����I+Qn���6�����K���MSE�xOώ�M6��Q`�K�$�U4���S��Z8�Tbz	�/'�D�ZUl	����u�YX���%��
E��v�Pq���x
|�p^yZ�r���	�J�W�۸�m4W�d�w֙����B��,���ܦ�UY���$5�*��PȄ��7��H���ʹ,]{ي<ei �j~F����>%�CP%Q[��I�a���~:4����Ei6�~-�f����QV�<?9���[8��Wu�,a|:Ë���nB�� B}Y��+s���v0W���Wp�w�T�S-0Z'��݄��Զ���s����	f㚤��5����z|���R��׸����[�k�+��L���?��:��? �� ^B�׀�g��q0���H����P.���f��[h�3���;U-  ����7��Ѷ*Wq;�rCD�j�V8����M��Z�;؜�B��6�-��جOiHN���|��Pc^q�!Y�I�E<g�ы�v7�XW��U�_�{�a�
tă;���Vv��co��5P�J�JX��_ug� ��2���u���c�6Qnn�H^�A��ǅ��#C9��Ji~Ѽ����{���/Z�/zG��?�+>���TY�(���IO�A�����B��2	�c��
�q��;�sɔ8������z����`h��c�X�A쾜z%�jZ�j��{�-�'�sG7��^�&��KM����*�e��c�\���
=��6 �����6���ͻ|���G��oʅxH���Q�)��z�?�$Z��g����В_X�,|�_+\dR�\R��IMVb� �f�%��?�bo�UnM�d�T@61+Ο˃�t�|������#��m�߷rp0F�n���孫(��O���ZSF�l�T�ZԶ�I-!��f�1AP�!+��sA�CH��6�BG����.�3����X�.L�;T��>r>����Q���3�"�x�)�}��)��j���B�¿oL�6۸^�x��חvI腌�:�ZԽs�a���0��S��$ϧ?������f�s7�����J�OH��~ҵ�@�b��y؀4��ѧ(�	�~�c�R�,]�p|/��Ho���n%�����,�&��J�xp�N3�rs�P�IJRCA���q���=H�{��)���fdK7#���4A9��'�8��0��j�\����M�"Q4�o�$š���Cu%���п��W�)#G�������?<»MH�ع��e{;�����@��]�~�K�R�]bJ�ڈ",��5���u���S������G��{ft��pY�8��hK����+�H.{��ZGWʢC^�*���EYwmڮfн�`xmU�:I���w�i�������zx��E��aR�M���d8gDnY�ް��'�-�Q���o��v2���J.��>&�#�jz\�gWg-�e��qj6:>���Zm6�t��9���Ug�\�W�"w��hs0���}�"�W4�8���~�HI��u�a%��LL�!F<��e
仪��?DJ��c�����h@�G��C����%5�Ln�"�;o�|2k���&=������e�{෽�)���e��y���`H�6�Ϭ+���=�9�3��W�k޼͍u����]l��cA�=)�J��8'�Z[��]m4EF6F7�h�OSY)��J�3!r,C�Dȳ���X@/1���h?���2�,Z҇X�f��Eo�!���)^m��g�yh��$�@ce��K�\�,V��t���7FtD�c��ܾ� Z��A�ŵc�j�/"�>I�+c���Κk�m9���{�XkA�!�B��k��2�
ZM�z����o�����?$[D��۱b���!��^�@�;�$�@R��|I{��{e*��c��QQ��P޵4�*��+��T:!!�S�����PM�@/Xۯ�]�ow����rB�����tJ
<��"��o��Rv�6bZ�Ctt����/����`�uz�E�c%&����jP�i#�9O��t��n��+����}nʳ��Vg	ʂD��b9�Vj���� x�������]�J}!-�ǯb��zY�)�kdR���lEm��-.�Oj�T�D«�!+~P���T��wK�<����u�LH��wbJ��ȞE)l��V�����Ի�����~@}���FL�����9�}�k�X�Q�g>q�Qv�:�z@y����3~P~�'=��/����=Ӕ�f���H�f�3���ҹ�r�q��7�����߶+���%�ޚ�{.�UN��R��|x��H/�;��5������Oza��t"��mI��#E���S�ό�ö.�M�lU eՓEg<�U��[y.ʔ|�u�t��(5?����ibI�.���nJ��3)���z*n�!Y����<2Ц2y��a�.�aشl[��9�[���ʪ���s�n�G?��e� TJ���~���\�f-��徚c���7Y���?���e�ܻj6X+��r{c�ӹ���#L�ѻ�ns�$��,Y/k⪚�=}�RV��'�S=�~i	K(��6���T�!^�M'|EMͧ�q�D蚥Q��EY����t�~�V��)��^�HpF�R�E����Q��:oivȫ��(����t><�F�NS�B^���	�^�㓷����[��ߗv@M��\��`�^�6�.�%�(��k���6���&��k��?h���Ϟ�3J�9k���o�� '3W���-�$H��	�E2�ժ!<�/'o��覯+F�"5Y��~�b�	�`> ����|����<���嶠��ے��ϻf���=R��9r�~�3�P��9���AD����Q�Э���w�:��K<�/-ܓ�2���9ߍO]Y��靹���2�'�b�N%���?�5D�H���E��s!*�Cq���U��3ٲޜ��?O� �(�A0�b��%�������8P���='_���rl�S��{>��ykR�#�ϷEmȀ�U�p�����aσٽ�ޟ�'�2a��*���8R���Kdm�m ��	�{�g׎�������nx��~g�@�SB��W�v&�c A��F�'�=ƫ�@S��'@w����s�5�eЋ�(}*E�6��ə0��)(^�\c�FW��x��8���q�x�D����=��(��}\q*l�o�f�B����U0����e���hd�e��!���}���!�	��ͽI�)pT�d)l}�4l��[�HX�81m~�$*����e�,^>L������JcΗ,��R�s���_x�yEjش���̸�s�g���i�������[)/��q�n�1芡���T��)]��D���~fBDMr�֟�GR��ʊ��䊶���y2_��X��qtg�=�2<��+��qu�ʄXX�7�`�}y�y����9mq�,F�������ݔ�b�h\���9E�L�
�ml����d)j|��_���r���X
��6i�\Ȋ�df��~L��C���i� ���*p���I�h|�xU�0��5�[Ot����Z~z��U�؞�sᨍ��o��^e,�&M�?�I/�U���l���-K;�����H�1���>a�ϧ阴���Jh;���G��0��au��S���y���@H\�4���*����Ȯ�nx��m��\`?ۀb",�w��Е�F�����)��z������M�;�){}��T�$BHE��7�Փ�R<<���_�{�j�'s}�9T�����JF��;�HO,���p��/xc��*��Y��s�;��FV�25�Mk�q{�s��Z>�j/�����W��������t������ 8�aQv�R�{��D�Ի���) �� F_��v��X��������)� +���O���x�u|Q�I���״������~1�l?�+��:�]�~H��]w:wS�$��0�K�ː'���@�ǅ��@�R!��c�n�D�@)���[�r�	z���l��g���1x��R$�a��wZ�K�&}X�Y� �b:����HG�F<�6R����n�@W]P���
w�#&�٬�)yM(�=A����X���dE�U|%�����`���@Q�<�w�*�o5
��۞J	�7{��H��Ä��VI�<	�uz��]d萍�n��9!B���=�����g�Qy<O�$?�\�;Cc�p��֒n���Q�]w��Z ��+�V���Y��T�AJXS4��η9��E�#v���ͮX�޷&�b�#�?�v�S5i��:��j�0���?���>�"�3�FP����c
�j�ԟ�C�vG�{�YmJ����Dp��,W�V�5�.���"BJ�y.M���\��R�Vl��߆r8���T���i�C�  V�%�vs���XI>��οv��N��šAN�k��e����ҺB���0WZ��U-Ҿ����~xؓ$�343��պ��Vq��H_h!u�@"��/��Y]o!C��۷Z@������z��3& ��c�h���7�CgA�L�˳�{��<����_b�����ي����[��+\YM1RF��Iߟ�^��R�By��XDN��L����q�F�����:B�0a�dq�3��8f��8)���dFh�]�"�`(,��<���X���l�a+���S�(\ A:;|˃�i����5#]�������(�G��q+�.����E�ʊa�;��Q���ZM�ET���e!�WH"ywZ�A)�)�t����3�%��P|�=	ݏ<?�l�(�`��}�������/y�ırV"Y�w��Ϸ���0��d\UvF^`F���o5 �0S�@Eԓ�H,�-��hV�sh�B���~�4��x��G́���W#[�� 9�m� j���=��BW
��8Ir��j�;�]����� ��)�i��Ɨmb3L,�Zq�m��j4�Ag!���iUq'�����"_?��Ŭ�L���E#��F_�<���0.C/�R��w&Yʽ�r$�Ϲ'k�P'�xEeFX�6Ե�}��zיj��Bֱ�t��4�Z��*���)�(B%���<X|��#2+���km�P�a�g�N�����J��.~IW_����x}+�$^�`��n�"�JtWA+���+���Kx�)#$�e,�On��cپ�{�����u��>��C�:���h��8�/����;��n�r�u�}8cHd�P���z���@^J1�����{�,�r��c58~Q{Dz�)8�\�١5�~XC[c�K�d���D@������#w��������	h�5JW��`>�\V�c<���g��"`�J�oI��A�C���7��u�0�E�c ���@2��V,E��0�7(��^�1ΣL�h�9���L}�G�f�#Wif|���Гv��6艛���3u�i�Ϯ��G5�+"ڲ.:Y�9y�A]2˪��j�z���	i¸^��� �LV2 P�����ݲ��ȗO��Fӈ�wK�?�34����	�3+����¤�z��n� �\iI���N0�[��7P����$߄Q2�bT�}��M�F��v>� ׻<�Ke�ø\<�4�y�"�f~���P�R!���J�7���8��v�������a
�r��*ֵnnC,�"�A�5��z��,��0 ��v7��h6[� o����~d���g��p>ħ+�FR��,�t��k�;��,fڦ�@���ՇM�ܢ��>	�pۡ̓^�E���3���[����f6<���P
���ˈ�>nJ�a��|VN�c�i���	ȹx�Z���&J�i��z̆m-��9HI����>u�.z��B��.QH�����60�\�>U�]:̎ٝW�نs�Q:c���2�p}@�+4H��Eoj�<�68�t1;fڃº^{�b����Ovc�gm�hm�Z��y�	������d�y-I���('���F��h�T6 ~��`w9}�K/�^���`i�č��Z�*;�G
>���FV��6xb�A���F��*�o���⾫REp Nco��!�S�m�#(~p�:��Lh��н�I璽�Oj+��h������������g�ɵW(������9N��O/���nkm^�Zm��2nD���W��تّ�F��`���-@k�/΄���U�y�R��ߚ8$���Cc�A�X�$#�գI��c���J6ܾ\������a苸3�_��ՅU�Q6xR���;��,���ژh��ɘ:�tT=���I�-�K�g��,� V�
���)�q0���Q�wYXp��^��4���z4]{sd�vRr���&���u�5�A��;F����X�$�]?kq�DVF���*��]瓐����dX����l���w�4.0��ʵc�fǸ���2{P�J|�P�_�)'{��Tb^�k�@Cj�����wb>��릧��E�?���WuU��Ĭ���+ˢ�l/r��WK����.�t���?J�&Ne	��S��;�O�.g�����j^X�]��Y��(y�Ϙ��,i��^sP��J�A	~$>�PP�����n�L)��#,w՚9?f�'��NB�@g�C��~0pCMz߇{��QIMn���و화���jZ,��u�B���,C��U��b;5V�=�Q�����J���[\���ۤrd��|��'��&��)�ޕ �BDr[�/:����q����~�Fi\�D�0�n�d��5�
�(���t<��
w���^y�T�忂��V{]%iy9v����3���%F�?J-i�����+��H,�L��������^��{ӗ&�0�Q�#2�"ʚ�e����G��;��%�
�f���$���j���#)x��Z�-��6�a�5�7Сy}�ق��WK��3W5*�E�=�x�����l�^Yjb��mI����8Xe#��Z�qy���ӣ�n`~�=���3��t���O;�d&1,���l(���}�U��6		�{�%E���a/q���Q�3�E^�N����ƽ�R�LHV�A�k%v0Z�q�"����3�#<��
���W~g�˦�k�R��Ųw�@E
#�|��m���=��{��E/�=�蓖}���/�td� �I<	]ۚ����`8I�T�Iݡa!F�>�o������T�5?��/�3;h �+�N����7*�_�"�뚷]C�΀�k(ْ����`��)z�ƣ��=�>VLw�^���=������
(2�ROğN�ћ{�v��S�y߾�W8��{�	}�����u	
�����8x������eS����U�YI`��'��ow��l3B��H�O�f9��b�E		��?�r�S�����lq������8d kv~N��'�̑?�z�{;?��J��d���lѲw)��rI�f�~ �մ8���Яj0Br�(�����P9�J��ѕ�=�,^>!v��bR+6��^6Vہg:�.jHg2�и֨�|���)��U>�ofF#7��eLb>�A�R.X�>���ѿk9������ŉD�D��v>b�ƩF�sd��մ7�j�$�:�W��2�96���-�K;Z�0�R�����Y:E���/��
��̭�t�|o�L����R�S�Np7��_޶�t�c8Ʌ�Fjh���̋q�����.�QL�l��=M��vj@���#}�(`(삢�(BL�,,E��瀉��%�)��� ������������N��88��:���v�=���s�U1WT.g������w�#Ef���'"f�Gv��e��N5��0+SA<�f�Pg���R�2vE����YAd�E�E	��73������w���9�V��U�4�
b$����ѩ�x.��*T=ۈ�ѝ�D�����c:��4���t�����	/{����}��FR4,=9��h�5��@�3���N%�4p�:�~A"�_�g�y�OJU��t�tN�0�:���E��3z�#(����+�i���'��\�`_W��W:%7�N���.K����4V�����^��eP65X/���{�ؒi�t�#:���s�"9�<�J�=��N@lM�Ro5dꍄT� �n-w�o�bh�,	���ʹu������~?����"O4������/ 	��lzT�YxB*Y�>Qybx����b��J�����g	K��Mp��'gI��,��+-�]�#?$���7�%�G.[��1�;v�]����g�wV�+}��d̏��i�ɏ�nA�0��|�RW��=�񑊈P��7-��MP�����(�\l�GZ���{3�7�SD�uؓ��I����]Q�ܺ�1ҸIH�4��,��� �w��<MxM��`�J��U&�Ɋ���f�҆����l:U�%���=�z�H��q��#B�Kt�%��4�&�Y��I�Ic�~�K��_�׋3��_�b2;�r[;ɏ�`0�*S�w�ޱ�')�"�<׮_R���s(�C'؃�k�����[oDA�Yy)���kT��p<��㾓"m�}�Y�p��k�ߵz��|�Z�^�r�6�m�'ˤٝ��H��T������q���gmoKb�lШ��gÕQo2ʻ�bR�\h��+(�ߝ�mTV�����Wǥm|Vtr���̯�����V@�t���Q�����>�ӓ�c����G�ۭb\ȁ,����¦!��/~�wc��" Q4�B&��i3��LqG�{9 �������չ�-FѥXˇ��Rȟ�M�B"_��w����(�S������x�s�A��J��)��~h3�8�%�񆻒J��9=�WZ)r��♄`uO���HLd�.[{~`J�Κ^��݃�������r�|���R��������@��vN���\�C[uԁ�U�6]�=Wh����u�P.�=�~:'Cq�C~�����GY$(P�ċi�������TA!�V��|�'C��r��E��,��M����N�yف�/�2.\Ax=�ڸ����	]�i$nIܩ#�f�x��n�*���D��~�{��id��Lc�B����&h���YH��J]�>6	��d�OaLdA4���!�*2`t��Y���X���7F^4���ٔ�� ����JHC�(<�ΚA|�"I���`�R,z�n{�+��M�B+tWߵ�-]��a?#�;dǃ��4�
�u "�����ŝX�s�m��)�.�7L���5H/�Kg��5P�I2��Ȁ
^䐂~� Kr2��S[�0�[p9PPxҤ�Y!r����o`ڗQ�+�� ��7T��*!۾�&�;4i�C��9b��|3�Ųmܷ�bUd)�jjd�_=6^���%���*�~ MMM_�^:L�W��HR��IG���U��.H��̲�&���ɓ`}v��$q����tPDa�ʢ#�n��Vm���jf
���-Aa2nP�k|�J:{��f��gy�A�c��lfl_�h��E�N�B�����U�ړ�:C(�À;��A��|ٺ��,�VR�	����ҙF�*_=�?z�)��\硵��>��Y���~0�ф�G�E�K�v�5����=��ɦ���|�G���2�������ުڏD ��{`SZ᧕ ���nϞ��cܴ��$�*�y��	��=%�[�E�o���rgi���m[���y��-�h���'��*�RN	�~�[���Cv�i�8F��U�W5Y�(���xQ᪵�hgDց������H�*�{�vƈ�C��B����EDr�l
��/עPk�J�0��tHT�F�-�ٲ�KH�&�����B���&7#�oύ��Uk����c>퍣*]�S������`�ߓ����+�?I'_�J�?}�-#q�v�J�s��_N~�Zo��I=��ڦ�瀁����q�%���\�aW~�(}
a�)����t��(ˊ�o=�G�D�=��Bu���!�0-6�E)�6'1�GYj2�E��U�xg��b���M6d�����~���m,:��Y
1tV�Q�t�2��8�t�r>����Ǉ�n%��.o�چy�l���X�R���D}"��鄺� ;��1�b뗤߇_���֧�$�o�5�Ԭ�W��ךNT �ӳ<E���`x�ʑ����HRCY�B�%@�g�S5@���$s��_��3�B/��MB)F@{�#��A1��B�{�f[k���%s����͎�CP��q�λ�N��ZJ ��9�ٿ�j�c�D��4y���T�!'c�kZ'�>�����q��oUmog,(�[�cV3���Mȁ��Ar]��Zh��8��܄����j̘A
�%zl4�φ�:�%p$-��{e�����z��^/�Iy�6��k\!�i�ɯ}1��!��������-g`�M[#��[�I� �idV�����;x�&�dB��#h6̒��S;=7wݷH�
k�[����d�M=R��'U��s2ڲ$��s��$^|t�ͮ�>��r�:�]��}�N��UنF_�T�v:��y3���� �[M�a}ӄ���gY5�y趴��Q�6=�����Y�u�s�R�k��	?��U>Ƽ�ǎ�������gt�#�����������Ø�d(�@���+�]#�\.O��E���2ٗ�8~:ȌV�;���s���/�*c���l��l�[�N<,���I7��m�����'�c���?��oG޸��;�#���IL5̊_�ާLp�4#Y+Mu�d�&d�����ý����o�A5��7Qp�������t�5�E}&sS�+A�-�\��H+�}�pQ�fN��8¯ӂ2" ��F�ZR�p�3��H'e8G?a�/۪��k���!��Mh�c=��!L��:��T�n�ɓ�9�fL���*��)���I�l-�pgl�HR � ���po���U��~��9܁�	/���r27���h�.v �����"I�~�qiS���2��'��\��R�/��#�HX�E����(����9=����C%�^Q�<%LԻK�2]i�X�l*��>��سq�W�+����S�%v�pW��l����]7wB���I-���hxy*dYip��{ي�M^�b&[�6�XG�S�R9��֕��,ʓ!_��윟�B�݃��u3p���
c:��b�`�o�!������g�o
���;Gؗe�&�����M-�$�1���q�i8; �9)�~�$�����r�5��ԏ�=�8K�I��C&2b��hB	C��b�o��cO����LDh��.I^V���,��oH�ɎM�AM�S�cx�>?pD++/R,�Q-�d7*"�0C��q�P�Ax>:Wbݽ.���Yr۾nz�z�^`�z�oT�{�����l���<a07+6D�M[y��MQ��;��%G�U�;�<��V=(�|����T�X|���w$�`��:�\��:��|�h��#&�[�II$��`���'�)�|M���j�d�C	���߀je)��I�\��Y<t�^Yļ4O&��qYld�bz!:��h���ڄ���� �AA@���@�(t�ɷh�1����k<4_�I���2�!'(��'�'&J͝�E֓���i�D��­.�C��]$�!��M���//�E��5�2�q*'���Z��E�X��9�Q{�S�V�-9٢�w';/O(��z�_�����5�����m��zƑjyΛYrm$��ʤ�@�%��*�k��H��0B:E����/!vSY�f�c��� A�|�K�<���m�1��z���s8��Y���Q.	�(�}�\Z�B�����huK`�<���.��Y1B$'4VbϭrI�}&�Df�rV������*�Q��]N�8��S#��95B� {L�	l�XqO��|[��^
}5q��.�Y��}��fA�X�_��r�*h�gF��r��+���&���og.����Ǯ�ėnI]ә4��Լ�!k�e��<�8u-�����4	KH(�����	��Eu�h����0�v�(���ec�y�}oXp&Ir�����C�E��j�ԋ��������
zwC6�&BW}�2o�)*=]'��88��;x�<M��;��҂�����@
��,oL��~;���Sx��:�X��h�M�`�P]���+&����k.D=�$�������"��|�O��o�i�IRR�\<Y�a�d\D��� �HnEh�x����������Չ��n�V:$R ���	1x�eVa���W\ϸ��Xo<!C6��'�u�F7�R|K�����Iv�XQ���@��V�VE��ҔhF]��A���z�.Q�����V�Z�艆�V��)��-�������-��K%�؄�On���]��fC��v׵�p�x����fh�����7*}���!
+$U�O͏��FeIR��|�7�k���blHL���@�i��k
fѽ^b�_b�6��2�~�?4�����~���Z�T�)o�\�����g|g��w�f�����}�&l��R���S��M��WXO���o��%�gy�\��5���A�F��dR��q���������
N�aɚ�u��u��^4���q� �9'�^�r�KRU�Y�p�W	"����|x�"�| 
�J�Xz��%bX㸼'�i�8�N���Y�Hu�	�(a�4vUΊ�D�#z�-��Gzt� 2�3	)Z�
���`h�%�Kf 7��}�h���֒��x�uS��ȉk����|����A~�I�9��D�t���28И���,@��F�`zu��P}��~8�8+�Z�0_��b�S"H�*�\�z�Q|���뇤��?�u�����y�.���p�>IPO	T��صzۓYe&R A�"`!]�V�>�ُG�	����?��ߌ��̗ٮ��_��etPf�M�WW�J�3w�vg�G�_��O��R�뎒Ԩ��_8�'������x�.������ן�Y�<�\T�$<�72$1���VH$DT������f��V��#X"Spso���=,=Y��P�`QJ�
[Xc�ʲ���d��oIih�l/!EP�?1/nG'�s�Ek%k r���(-iHh�Nn�܌oWx+�8�)�.�Cy��;�Y�� h�z���z��ũ��~r�iL�Y%����o֎/��Xf9��2=|ۥ����>�֍Ջ��|�@��O8�N�H8[����d�V�L��k!q�q1�@Y6Q�μ1��e�#[��1�0՝x�+�懨�ד� �?cr�����ʽ�2NI�0��Ǚ��}GBe�M�A��S���*i?��4�9�,t���%������
��������2��e]��6K�fʲUx}�-F}�l
�N�`��͠�ǒgfӡ�J�n������3�r�����(��T9qj\����ÀY�o�W{�L����M�v�ѹ���.�H������E�0%��U�[��{R�����0	���p��`_���[� �W9/["�h&�h�W��o�ks���QP��aR]xc;��6�G���& 8��O.6�q,����@n���q��iT��0.>��StF��/%�~q'A�'!XR>��{J��h)��פ�74�:f%E�?��ΪYͤ�p�h��5Y��Npa�B�q1����D?h�NM��\긏ٓ��L�+����X �Z����T����H׌�����m&O�e1#���a�Ȃ�W�`I�� ��ȗ���pf��>
ĵ�[Ƒ�
�3&��Y����:E��*��;n@L^�A{�Za��D�k�={sĲ����4�lp��e��e�p�i		�e�:���HWi>]��̖��_�J�=�����bڑh7Q�"�ť������Y�%��/Y6䵶2�T�y��	άҽK)��N�~+�7�Y{y�@��� $Dr.�01�, �i�p�sU��v�.�k��օ�����^>��Hljn��y����I��n��RS=�T��<����D���	�%��a&��SAXmK�7������=��'�GjhXə|��H�b4��n��zh���M�9z	ɭ�94�H��F�T[�+��Ĵ��q;�7��5��h��[IόS�;;��e�=��r-|��{��\׷��������ݧi?�i�s@�
�D�G�%�����f&�@�<���~F���\Q$��#�ʕ���Ѓ0� ����YI�'�
W=�rKچ zoa14�O��η�\?S}���Z�up*���In	��'w#N�4 (y!��⨳�׻��ë�L JK�@�q�Scp���y����dsɵH-t��F�]�Vi�Q�%���"^�V�	�43ܹV�DEi����y��~�o�jU��kj�<�
Gl
V���k��V�jdņƌ+���oh)5��2j����d٥� 9�?O�r�y�{��ׁ�{��0~�@o�(�ځe�{]���zt,^�;	 �G������R%�`d�'�3LϽ�FL����x͞�9��?.�̸��-o-��+�A~a��S����d�؅D�y���e�ץ$`� (�]>0�3�Y�;C?�8oL7����T���r�H�R��;����jw�چ��ݶ�pE���z;�vr���.v0�pZ�
�3�9��fIf7�.�(9��ܴ)��^���Y�
qks�FO]����ϓ�ӆ�{�;�ˣT��#���y��5�z���޾u��G�U��DZ�gR�N�>�U[��j�t'���o���0�f��� f��Aʯ&�ǝ������ս�{�Q7?5j�ئAwu�kҁ�T~u����f��0���{Ӽ��O8�W��<X$�{V��t̖�Gگ�3.��_A��I�ŬVzDsA����9��O/Emq7�W�y>1c��O�8�{�oq��{^u���L?VDv�\�(����$�E"n?��ν���0,"��#7ӏlz%�ex{t�����ͩU�h"�Z����9^�b�7�O�J<��;9O�p4IM�<x��e����aNaY�U���������	k����ʠ)KV�Ŕ��UH��pL�9
�ָ������FP#��gR�!��FV�*�cG�ǳ��`u�Qj��˷�Y��zȔ 1�f����=�2���z�1Re�v���L���zU�£w��v�YBz�O�Wcm~c&GbW�@kP�	��={#оֈEȚ��s�(\"*Ӣ���g�� ��6����s���X��+S��J�
��g�sFb3����~�t�50�6S�=�^Feﲂ?���͠7)���_�Z�xG������tY�us�dN�IdҘ�+���c�WQ2�~�GxElI�p�B��.��J=��ARp�G@M�?D�W����sn|"���|�D������l1C-���M�����o�>z6a]'�s0:,�|O����O���g��U=���-�@/�8|�K�m�^��iTQ��3837�>@_O����x4�\���<u����7��(-�r�|�uc�r��.��l�����ѧp���'Eg\#tc�j�I�E���R[g�~�F�I�7#����|�׈�|{��~]"{D}7͗�a<T*Q��8Խ��Z}]���R�d�@�ȣg��*o1w<>oa*�pTx�0*�~0D�~���^8��ȉ;Y��u���Ă!�/��H�DO���?�\�/W� �? ����^�@�cf��~�z�B�����Q���i��(h[Ί�T�j�o𤌪J�z��;�Y?���FSq�B/i�\V������o�.��)�?g��":8�W���=z�G	C8�`����g{�1�ܮ.�6]8������`�ծ��*�k�N�'��=?��(j��_Eҙ�����ޞ�b��T�|?zia��nWU��X���?�@��>o�HY�$��؀�g>{��j%��7S����o��,Lr�J�Y�¨�$��jh��0��(-s�MD���P`ŕ�$��+L(�
Z���,�6�8�T�Z8^o#�o!��o��j쇨 ��2:炖s�~d#~�`=��nG��}/�+ț)���	��u{��2]�����-9%��ꗔJE}$�],���:�0ŷ���|�
�/
m�4����i���7؂0�n.r�O����QZV���G�&� �ު%��i,i�c�39A2"���S�>���B���k��I���M�[q�Y@ȡ�Q��>@W8�V�sP��2B�3��Z�cv6�*q���Rh2������G%j=J�Q�W�-��П2�(W+Z�� �R��-�1a�h�cf�`����2u	�Nup��_�����u5{B@�L#� �;�J��w��>�\6�0������wjQ"��)�r�Ct��FM��w��U`��>2��{��R�(��F��&[�1&��<5.���ו��Pb�F�6?B�^9�
ب��p��J�?;��3G���>�o�?�b�ͣ��3�M�����dr�4��z ?�>�QPl���D�Mi_*}����mt�Ԙ�]�e2T����r0��eb�a����-|�;�Nlk}�Yx�
dGN�M��[s�3~'�� Ѽ���^\�􃱅��7G�5U�R~� b�R� 6_���G��6۳>�Z�}�fd��}�Cc�o�תBLQ�z˙��c���Eӊ�(������Y�o��к���5��A���_l^���>�j����/���N�4���<���������m����Ǹ^AAI~)]y�m��ƶK%ɝslێ*3R�:�A�:�-/xPx�R��h�Y*U7�]<��G>	�Q��n[��|IaJj]�\l�Si#"Z?��l�Y�G�e����n��K�1�'��B=�j��t��s
>����ʲ�e�!	�Y�Xކ���i�'���㔉qA�M��w��?|����'�卆$��D�J���T�{O+K[�"�iZq|a�H��V8Wж�,e4E���K{�]����èy��^:�����kY�u�\p�V~��"@��#Q����E��6�D�'1}�A?�PX�m���[z�����TE��E�(fj��C�dN�;b��؊)����d��`C�t�������?�>K��M|u�V�K���\�K�h�hx��2L�1w1]M��kH�F_�.�nVIp�C�"e�0RJ40WW��	��O��.B�QPuj��>��`4 wCj?�]}O^�Tt�H�@x!Z�x����w�Ō�9O(����*U	�{�� ����@H�Vf|[(1ŬCtt���`���Cy;�0 �u�����9A�|LB�
&�M]�n2.�9
e��q����� � �x-�����9�hl��]�P04�-bw(x}��R�g�����S�ο��������Z�"��b	tA6Q����H�ݗ�?��@�e�ڝT���Љ�oY���&k�4�du?mɊvK�I�	��[z�?����,�O���
֮�vZ8RK��5'���X��Ì:�O�Ȫ��]?b՗2���}F�8vZ	�[L�|�Ј��i�e��i��� ��#ׇkA};�O=2��Γ/��֧�Ō���Ej��Va��]ˇ��|V+g�{�Tޜ�j��A*a�*~q�+����捂>ܭMN������ϥ�M8tK�F��Q��x:!dd�t��"y�#Vs�.F2A�W�	�Ō�f�%��dKl�b=��}��3��
}�K�����nS�l��/� b����ZQ����d� �S�"�.Ԧ�� �Ql����/��a��3��H���ޅ%yz��k�F�)�N�%���8ޛ���O�99k�:9-Q�M�#��F�n-�Z�AǴ�LUC�K�WG�5A�z�}��t���օ�aӽ
�����m}���j��$�r����.ę܃���� �}�%|�S-�$) �Up�9��Y��9ǉ@n�~3��x���d&)}�8=},��C�Eqq�;ƈ� �L?e�K��Q������$�0`�������g�X�1����۾|ܩi���8k�0���+�GdBq|%o$��6�  �4�B^!-�$�%�����R���"�Fȿ̐G�=���¤d k!��q�)S��չ��t���&��c�+���~���7�l,��I�S����y.Kd~�� �cb�Fd+�%;W�N�Jx0S�E�l�lYR�����O�)Z.�|#��6�v��$�,�!�t�R��i��z�+�jT#��/�q8؅�_:��fq_Jl�Nפ���J�C�)�@� 徻u�n~o���.�A��\�ɲ��T�i��|��x9G1�w7�ߴVF�*ܴ�<�Ëֽ��q�sF�/�����h�IAY}�� Ѵ�&��o����t�^yP>�N�����,=0�~f��NRG���b��nB��Ym�/6q�[��Պ`_8h�&��\\�����]+�]xr�}�̆�emf�d4c�Ѕ9��@�-��}j.)��wah�JH� ��m2F�9*F�Q`��X��]��0/�PX1��rwE�Ҋ藁�^���[7,���O��N���-�~?z7�t��'����2���%�A||�]��V���(ZU=!.fh�-�N�����`�炎aN�}�m/� #��:{U,�e��*��]�e�Q����q�D#�V� �����r0��qͨюy���v�鵛��=.]j �����źjg�͆
qc�d��'a�A�xr�m�*QX�Eq%���j��C��7A�#F$���+w�VQ<��wVƅN`��B����X�ՀK���ŀ�+>i8s��v�Z3�;�-��ǌ�:���n�/���_��@�N�h}z"&�FO�[cg}X�f=��]�u��si	s���|e+mz2�Iw�N�xǨ���� H˟��;[��b�{!i���|dg"�� ���}�V_S�R�UC'(OC\=\��h`#!=E�à�L���[�B<�n�aPfO�?��T� ,��G�x����u>F�ύ��Ǘ�˚���$Д2#v��3k
̚�Ը�^N�}m]ܖ��o��x�����G���3s:_v�^so�n}�$��)7�M�}�U"��r��7@7���~��)3'.˵�Zz	p
V	$�~������N�?�3��f������n�y�x^��:锷�Y�ִ�v��+�F��n��Hr͜0���ɲS�T_CC���.R�.wWg�SjA�4����f�
܍���ot�5�*e���QSK����2^��t E�#/0��U�k�l%\B8pF3{���Y_���yOK��9��Ҏ����^��>מ�_rN1Ae�L�k�w`2�#Rni���Õ#��Bà?_0?�d��w���%t�YC��o-/�o��#�Ǚ�\u�|��U`��6��H	�9��g�{�Q=�7��k�dՌ�PɊad(��w@��=9�"�c
l�q��C	!6�U��� ��Z^%�^��]��/x���L���+t�_��r%����^Hrԛ�[w�']�R�O2:����U?�e"u_R�'WL�ʀ������k;)�l�����B�MS���r��� qF�S��$JC���-Ō��&Ab|�6�x{8hk����a�͛�v/��l��)?w��|�R�;Q)a�c�RM8��Q��ch�]-�D~���*m�����H���w98���u	
i}�aW�2�h>X���LQO@�������R9�V�?�r�-�&��r/����-�͘D��t���&�0���C�����G�/�jo�h�Pz��%����p��R��Qg���=�?��7�zHi�2�;ѝ�L�H��m��:��z?�dw^T��!��i[0�!�@yxDD��J[?�"z��vPўcRZ��w�>H�^�w��1(���^���ZL�)v���r@����R�3��D}Ro�/��:~v�SE\���U�T��������K���e���#��ل�	okO�����b�.�i�IU[=�B��]� d$�?a����Oe,�A5��!������2�!6,=u�� ��b�v.1,ʗ�E$�&95CIW�ъ�`}�'k���n�Y95Rη<NK�8>V<�ڞ!��(�Y}%P|�N�_�֧��.���+|�}g����F
N��u�D��J"W^�]���	|�d�s�\��9�`h#�K�Q����K�}���K�����8�Wq�/L� y1\\B@vƋ�J�T��(��i�d����� �J��Y��<T�6r
ӇM�Ey�d�n~79��boN����y��{,'b�:��dsޠt���ܔ����6�� ہ�ь�,#҈&��+�*��zUo��P�:�-��n��0<�*k��R��Wq��`l.��ȍ��i�zO�������n�	;��U�\[��O�QRmX�V��3�-C�D�CM����Tȱ&�����A!Ԍ/NX�#��l�ۜ��>�a͜�e-�!$�H�������Eۢkb����8���Q�7����[ah��E�)3�q���v?��3��ކ�&%��,���>L�t[� �����pG���z�SM�������[eK���U��I,G)��II�3؛��c(����T~��fm���_l��h"��dCV�s^�Dj�>/(�'%�Q8�_�VVI{x�ͩ���n�4GŪ�1���� 5�k\~`v��(�Z��K�S��zB�6v�V
�D�w50x�0��mW���A�ɎV8)�#��Y,� �RRo�]|�g� ���Jg��d���jm2R�fz����5�K5�ZԜxI�蝀����5`b�/��;�=��	���I�u}9�md�" ��I���B�O�����N[@^�@4%O}�ѧ��[����'g�_�o\�R!��g�ˏ��-Xp�ja>$C�A�[�&���a��ଳMe�@E(��͉<���(���X���W�5�H�$��L���W���մ��8�����
-�V��{nJ�>��O��5���sl�QIf�Fb�>u�{�+HC�y��5*�w[d�{L�ۿdE[��M�^� ����=]� ��BQGx?�<�9�D�` �=�L/�שּ-ߪ�H}Ny�~cd�L���ߪ�P1��7���|HL��Q���W"�&Z��p�,��F������I62?M�=}Pz�w��9�l������N�2_�ͅ���<���4���@�b�I�%�P�j.Ǘ)�/�+Ԍ�Dy�K�y��X�f�`���+47G����m��֓�����t>�Y@:xΙ�w,��~C�m�6%�� T����;C��VS[@�J܃���w�������P�������T����pll}Gi~^�#�[>��ӿ_��;i,t��Ǌ���qM(HhM����S��ݨm�!M�1j���ֿ�E�%�J�xL��@_��ʄ�*��|�f�?=\��a��S��
ή?eYџ#g���x8��M#�gw-�<Y~ف�>��Z���d�ޥΞ�P��8c���o�`�׍���<$ځX,% �"��%}�f��*XEDR�n*)^x��TS:i��k�>ʵ�.̫�&T�"Q�7&W�s\���_b������3������zѪ�����l{5I��r�1G�v[�5�E���7��˽�3eB!�	ib֪��Œ)��fUZ�����k��0UM ���u�U�,��os��u�U4���y?0�2Q��ⷉCQD��7�{�&�p�/m���s�+�	�Z��l�>A��(n_Q������(p4�Mr�PP��k���A���-#w'J���|�+���'������g]��3������\tu6L�K�(�����&�Uch��'�+�"*(��]����+�Y�zl��w!�Q�^��`�c�5M7GX����҆U�q?I���ũ�U�=�L��@�T������Y�/��>�2�xYT�iი޿�鸑oy�ke�+R_��$�9K�ۚ|�՛_�+�?�������0mg�+�QF�Di��+i�z{�g	�-�L᷋�5'�@��Q�
��A����˗�pW)�2���]T�?��������� ��[rW��V�����6����M�u��K15�wگ���	wg���qL��i�o*z�L���O���=����{�^Y��g����&TR�������;_K��1�g����ƽ�i�ؘT(�'�\�����D"<��m7G��)�(
��O�������7��KU����7��ve~�a�na���_ʻM���g^���!���K�]�t��\n��������C�EQ����H��W�XG�[�Y����q����QC���+�P���M5����vNV�i�iZ��S�}�G�Z�ɽh컧'��i���p�la��$,�l~U���eOp���P"w���R����A�3:�lu^Iln ��ggd��_1��N���?���RF�����K��qq>�����㳜�g�3����@i���5P�2[�B�o �N%w�+x�y��{:��\f����c�E�h�w���y|0�jn��(H��Q�������s��w��d�۞$��Ȭ���`R{t`��c�3T���I��C�~1�܃��19��/\�].�_y*��do�,�^��L�W ���J�[��\m�'3ԁ�C3L�*D�4���8u2יI�2��OZ�3����@�u��ߧ��q.��M�g�V}M�}[�8e�����y?��n�U���ۿ僟%eL.R�@%��#@S)$���AJAFF1+Cg� �CD�2�Pd��K�5���	�J�-�5���2�ihI�܌ħo)���%��~� kx�����][��'�I�n@�+P����f=��L���m]3ϥ�{3(<������*��E��sގ��2��0O�A5�Ӽ��EH4���%�K�$�z���[O%��>]"o"V�����Si�SMg�z����H�8<7�fT��F+��t`�y���u;�FmO�T���٠�8�����ӧ3۸�0jU����(����J���ڒ�r�j*���n#�._�j>�K��v�@w��}\j�������X�����n�[/�J��F�'{��16�"����C����Ժ�҇��PYvoG	\p�nG���C.r�{9d��@�R_��l"֣y)G��`�W�E��,/�����`	c�_+#�nm��G4ZA')t��@�LUJ�@��FE��4���}�+����Y1Kᒀ���<;��x�\��(+&�i���[�LI%D�M��̕˂�fI-�����y��gi_��������sm+]���{dI3���Jq��y�ߣ9:zޙ~+����"������r6D��hX�,����}�#��N��k�"c�LW�n����t�ܦD�H�g�`l3�����4��gkٮ���*(Q<�T��,��'0��0��8�y���U�ܞ7r��������a��l7��`��jC&���B�f�ׅ���u��̢�7bXQ����&[:�2���t?	��ڞ�W ��"ӕޣ*`�H���z��;�d�~�f�R�A�m	��
?����Q������^��m�>^���>�����P�Mݸ����DmD*�����pQO�l6�Kv����V)�u�1}�"�Wҩ��씽F:����U���7��q�Ks��7x<M΋R�i_��'ʱğ9Oe�bkX�C��UDc�?�z9�Mf|�J��	sk�u�
�ٝ�(�|ɦ+ٟ4MX��y�s�9m���C��_����` =������t)�_�K�h��O�N�|gb�,%���}�X!���N��<�"��<�+���Я+}W�H�����
o��H��T�ki�#f��HI��Y7��6�wx�C\a�T.�a���;�����3���x����R������l\t��Uң� v�.Wb���R�����@Qd�PH��E��|q�3*��)(���k��̡��S��h���<o�Ft���j�ί4Nлv����[�oA�n�_�o<_,�".���S�~�ؗ�E��	��x��Y��{亷����~��k�Z�'�"�������4S����e�CZ��k����j����?��U��A'�uP�ά�)�G}2��?�¨&Y�X#��~��=���Oy�ҪGs�)����i��׶N��uG1B���/t'
p	��]7dTa�.��ΌB�%����_��J���߷���q"�)�v�}օwL�B��O�e4|��{`%|H���N��5��+5�e��"n8F�F�>���/]��Xn+)b�����_����|��O*f�U��I��S���6�0�EXۃs��>0����Ż�nD�VW&1�=f���=���4��<D?}��ś][�����Ѕi���{FƝ
AxRs@Q���7k�o����_�:���Êz�X�2|��h.LZa�D��Wr�2��I��S�V!����2��QK�����)�vi��9T����N�(PT���*����`��FFU�/ٽ�	*k]�|�r�@�k6��	q A@�����p�5+��UE��G&w�"�2���=�y�������Ջ��Ж#�N�$�ϭ$b��D��4΅����󍮛3�k�$�ݢL�!�z��}˃�f�P����.�wkK	#5�Ђ/P-���?�tv���=�&s�Ǌ����k6H���?2�(E���>��fxY�|]���/�皽:�����'	Ԫ�Q?�7D<y������ o7�g�b�b�'ǿ'4���u�"/�B�i�w�@N�}�a���lyK@�I>Y��;��l�P��nm�p%;���g�=��*?b��F��/�OU^)��R���+�k��8/��� �G�2�ǆ����T8��bKZN3^��4n�g�̟<��܈��h���5�����c/�vBf2��+]�ׂ���5Xy�����t ���&������+�g!eDo�p�y�X�$��5E��B3������'���s�v�j���,�{4@��[e=ܬ����O��[��"���9jp�GV0G�B´q>x����̳߁;-,w�+�ײ t�aް�����3��ǲ@�W#6�+ �$���5��`��R, a�����z�Jln )��S4@%�"P6�)A�,�?�� W���t�s�U���l{ms�d|*h�i�S:���/(g�B8� �7���.]d|�vP��A�c�ǝ.�{Mu�����=˒��jIT���P,�L�N�W�ϒfn�IvP������髄�f��:b�I��S讅��atr5ٗ��8%�wґh¾n`L�Y�zZ���� I�j�S?0i�p7�)U~�,O��I�!��������
���_��Zw�qU�l}�L7NuZճ��)��R�<�5w�Xh��&���1"T�����ڥ��җ�Ǔ�Jz�4k��FHV0%mCTb>�No��)��Ė��N��ck��}>�O�,cÞ!����?�A�lX3jA8������#̑r裻�>�x���iF+��3|ij��-�R��JC/��>���������צ�!m:�`J�窊�q/�ƀ��H>����;l	ĵV�L��A:c� a�{��t�\wߘ0b�M9��4L�C��)*D3�t�s�(x�yh�Q6Dnآ��d6l&Q-��D6�	K2��@^����W,�
*9m��7O�*?�T�T#`sH�6	4g����3��1�-�z�\�^م���Q�:��w�KX���=�΂���9\�'��8�ל��G�E!ڙ����3R�V���赐�=��Oݙ�=5���l�R���zoG=e��<�i�ےK���Q�0�#�ޙn��m8؆'2� �m���ע� ϔ��?X=ރ<K�w��xI����g���b�p2sy� (8=I�<�C��>n_d�6Ս���4>J��.�@�q�	|��7D֩���''���`B�	�H���lw1��X+ ڮ�U�Y��)�N�C=����9���Z���O�z<لn��ID�Vg�����N!��.9�>��M��Hz[�k�w����ʿ_F�ON�m+�����q�x��Q��8�X0��	(\��������e?s@<*���ZO��i=DB��V$���.�M��Ӏ����*�� ��-v�x�@%@P����������e���V�~La���-��H��bF���7ao���o��K0)�����
�^%������[M�F���/ӾHZ���{H�,(M5p�A;�5�O����9�7f�H1vf6��5�r1�m���Y�$���]	��W6Na�t�Zǒp�pit��W�~Ӧ`����1���4�_w����������||��J]X���8(����M�z�����^��<�z���CK�^�WU"Fܤ�~N8-o���'��w�@E(M�+MJ�&���BE3�߉���p�}-�Y�r�}G��g��@����]5v'uJ�����C
q��{����Y|��!�/�?-����Vg�W��������%�T|,]m�o9F:=��6��*n�d���QH|��KD�b(w%���g��Q6.K$�c�$7�H��Q�>�=�Ҙ}HN(�]D!s�3���f�a���*PM8�h����*[kߟ�o��m�kfUnF�N�x�-]bo�m��A���Ϊ�oA�ps<cm8�M��N~7�H]�o'��9�
:�r��ș�ƧpC/�Cs�����-�ʄse������«�ߚh4���CN��t�3o{�˷]�6��5�C�jj�0%B@^2��_MU��c8J��6.�$��`Pj�Nrc���w��I�֨@Ë�T����$`6�dU^����L��>�>7"Z%ʆy	�BW&n�g��^<I@���l]���d�>���IL9s_��rP�l4�c�v;7����2�"�(�G����܋��)X��R���~w��`��3���$�慩��!��f�gnJ����[r��~��p���fn"1�~�CR�K�yD��aݩ��.͎y�/��N�V�����sƭ�]r0���X�5����%b��{�5A8�Z�m/��<K�U�Cb,�P�
\���r�^�[�x��-��)�~�
�5���\_�λ�0~_�;����v�������u]���9UoKF�e1ß��T8)���/@���(����d69.b���>�L��2�731B�''̟^c�1#��ض l���Q*b�nU�[-(ڝV��Th��a�EU��e�.�w�vdG Y�V�o��[�<��ͮ�O9���� ��! =��c�v&=���
��]�(k>���g�����]��PT��N��=��0�uB���Z����!��nj�s<2��:-�04���<�6�|x��Ƶ�$;k��:�JXf}�����(g�.o=f} 췶&g9�m~,��wQ<�A�q�s.����ai ����B�`ahoY�.:�S�.��x��V�' f�}(�lf� ��&3Dz�����O�e�og�ǁ	1���v9�?�+�u\��w_۲�A��Ț���<;�T���-��y�����q�lqK)=!!��{�U�L���R����E�u��d���H#�x�ք��H)����%���H�e�iǢg�v^�#���r�d�e��lAj�_�]ٲD����1+1 n4s�`.�Yg�<�%��I�ʻ�d3o\����7"�lf
�9��A�V�!u(P��Z�C:���@n��Dja���*����`�3��W�6��Կ���ذ���lO��U�rB�f�n�H���E.�fq�i�igD�yT{�F©�`>y�z��>��;��),U:��՞>v?�Z.��X֌<�0��dƎ����<Wގ��m6{#����z�b��VH����ǥϙ�����+ ��~�-φ��w�5�۲��ܷǎ�J��ҥ���-m~�i�gBΐP%ݳti��-5���1����zh��j��.�����v[�3@�)���$5��,�ث��h7K��ұw�/�D�@t���i�;���끱�18�	�x�tX8���Cr��@�8(���Q��
<
����RL ͋)�>�5$劣-���Q-�B']�����k`�P�%b�ũ)[?m����}���ߥ��Vv��l�,�~^Q(eԌu��>a LvW��x�,pX�cܢ��&�V]�"���A��2��ɟ��$5�;(�25ɕ�CH�� ��׶�d9~x-礰 ��V�e����Ϻ1$���8ޓ��()\
���,��\	��*�O�ȭ����=ݥH=�6�h蛢q؂�-�	���m8��w9�Z^`MWtvV)KX�_�6},X)��;p�a�c���B����.��|�B�0�SC�J��Կ��0x<wE1wFQ��[��W���G��6�.�n~�H��Y�Rf�ר�TR|t[��1.sB�z60�������ԳZ_y��2�`�| ����ɤ݂��
�Kj���+�Rh@����G�!1�.�b��ꮬ�D�?�p^|�U�)	I]MjHB���L�,P�Y�ބ9�au��U٣��=1�UF�p[8���E����4��4o�Ũ_��R2�z�I��7̴���Z���LamG�:y�f��%�������Oܠ���Qi�ҋ� E��O@#q���Sh��^��H`��_��?.����p#~/i��I���vq!U�5�wn��|�+�s[^V���e�gH�����4�y�L�B�ҭfq�`� L�Vب՞���(��BXҋ�G$�-���9'�$O�\	���a���՞�x'��L�9໒��d�Ĭ�׋���	}�1��]���۶��6��9�V��s=��l��������{���_400��K��`|2~�t8FVq�n��p�̉A z+��%ve����Q�RЀ$& B�������Ҹshj����Z�}���+���9]M=�'<۩@NQ9���'�r]%P6�����R?FAKߚtޝ���H
*����ѭr�5�gq�\��ľՇ=�H�K�������/Ê��Ϥ$��.�������y���Z8�m�q��p������(ăzBN!�_�{�wW���=�fs�v��5q3�
�Ԗ��.E���a��`Č�9�������;Z�b�`ǜ*�H�E�p�t ���7)y�|6�-G��W�5K2��� �1\E����(7�� Y�SZ�>l߸?�!�z��6FW���1��R$�T·�I�EԊ��Ix1��a�ʹb.����a*�~.W����JI().�o/�Q5w�l!�G ����HU��j���}kdk�������\�/z���]�Ŋ��G�� �������Q5g
�T��~��!�TזNc�}�Fu���W�x|�^.'�5������*���ȣ�w.��3i�ᕁT����2D�c�jm���܇�%���rNu}�@�b�Q̧>H����Z�t�:��A�ܱ#w����'���y�}�
�Ͽ���0	��k�V��������P��]T�QA@uf	f?"A-8dI��PF�]���B˗٦:@��:T�?3-w:��ڎ������n��2Q!ɂfq��m��o
k�[� ��}i�i�F�]��#f<D1��V�������[���0�;|��LvF�l�1��:���Ƶ�Q�Z(�F�Xt=M�i��=�mώOo���rrZUʉ}:oq��'�>NB��3z�V�ϏNշC_Y���	"Lz���U����W�<�{Z,�h���5��o��o�j$%@�ۯ��IN
Kv��zEY1XĘe��_�>��˪����׿�S���F��~{)1sc9'm�MO�i��x;k-�e�P��J�YKoӣ)�Qꭣ$����MY��o����SȚ��!�Ё`H@�p8�%���G4p��U�jh��E���;�(��0c�ɡ�u�dh��2[��Y�Z_�y���S�M����9�jB.v��*��ι�.%�[�'*/���ԞLCD9�i-]K�B�Q:V�tB9���X#�6��]=��ȼu)p��8i�o��4����,  >�����;>��M3je�:��e��k�/���΄�K1��;V�\��#�)e�8yyN��
�w cl�"?תE����ѝއ�*�NM��yp�\:�ra��sc�q��#�o�b�ۜ�,
A�褀�O�l���۲���<�o1E~u��Rq������a~���Z�&:���,��щn�fd�=F�م���z���%#`E�v������-�=�J�촭��{�%�����\#=d�yf���>����&�1|?�z2���a�B�'0�i�r=v���I���ܳ���^�V��c����X�of�v�66)V;��e�b#M�k��K�וE�/R�s+���2X-$�a��[��|����g=eCe��s�NpghI3�J�4�<M<�q���x9	�u�z�¡���q�P˙�:*UY\t�+.�{v�F�-���PVI�Z\�W��Y ��^�a�! �a��!BMd�$@�v1��dmj��D�Z
��O���@�"���k�p{=���y���@Vm6eo��_*y��?~NV�x�?DV���d�{nc��h�wM���6���@�$n��@bcؑ�E$%��
����w2��~�����r�ig>��L�8��Y�:R�2f���&���z����ejnB(]�k`h���$��ʔk�'�x�Oئ���ؔ���[S]1鴀���?x�E\mҷ}1_v/�v���.cf�b=I���c��ٶ�WV�y�C�0��K\|��$�0G�R��L����
H��2�E[���"D�Xc.�MO|;�%���+{x�������Fܞ@֖�V�e�.�u˃;ߑ�>M��Q��C�^���	�>��ED�H��/ɵ��d_�N�]�kc|�l!`�!�䗦���v�g��]ɚ绔�ǁ���ĕ��;.�c��ij��'$C�R%~Ǆ�!\��k{�Ϲ}eu_��i��$�>;�g�|�1�A�z*�2��f&l��_�*P�D��N��Y�Ы��X����Q��Ǣ�+�j&5���z��Ϻ�b�Q�� 4�r���`#�������K9��vRy�F��Y@VŇk�H����V<��W$�+px���o� ��9a��R�jo�d>��`}_���ɛ���f���i��z���Et*��e�)Tn����;W�p[����,�t^E�1��=�8(��.ge-���͌k�[cG�/~)�����}�/+AJ�Vd�$�9D5����loX�c�K���ށ����%�s��Z�Z;��M.�� Gk���=L*+����چ�J����Sm�<���?�A3J�E.�%1��^+ax6Z����_S�<��O�>��ı�W*�l�uL:�L��80���t@��n��\/�.n+��	��3}(M#�)jMl�����*Π�:�W$����W�6F(�X��M�rcBK�c����ۥ��$�� �3�}ݶB9��di��}PV��̾j�J�����b�DD�q��C�ꦔg�7N�r�W1q�M,�V&������`�|�ga�
֯�(/߀�QԜǪ�8�h���������a��ѥ�دԞ���=G}m	�3;�ƿ�g��GX��m�ˑ�D�-b�1��+�n��_�N�^��G(��+�s�zRk#R���ä�k݀��cm�*?jOb�������|�L�z��j :_���^q���h~��HjW �qwʧ�섿�.�A5Qi_j���|mz:���d�DBR����(��E�amȂ��Lu�bR_8%�*@J�#?:�į�\��,3͏�����0�e����� ��?�m��d�4���F���_*�|n5�9�k��/��q�[Fݶ���Q7E����oD�E�>��G��{OM%W��J-��X���䔷{�ft��f��׼I�u�˾�g�ÛL1FV�uy����O��D�>��W1w��]Us��	]̩O����ѲD8Nh�����6���gj�?,cE7m�1��[�DJ�yCf !�9neW�
l�;��n��� d��;:��5X�����\���"� A����q�H�qUmi��+�>IC�ZO"�i�vG�)v���=Z���yD���,�^������"�K^Z������`lG�n��D� �!�4����QD��g)t*^:��𸹹I���^v��6�;�<�n�CE�ךR����g!p;~��{�2��T��w�8BC:@^/�w�}\�Չ�.d�D"�j���k>"��hZ,H�j�A(�:�rBN"���1�����K�;ĬQ�)}���B�:v����#�y�fҔԙ�p"�O�"w��WSt�Q_�K����蘙�!��E;��њ�}���:�E��%Cgp�`�t9 !�X�[�1���Q]޴Fi�,�c�GHxp�fu.^�0r!�UJp�`R�AMFC-s9ǧ�5Cd6�V�����.�T�.'k��͏��*姅�ǒ#r�-a��tq�0(2�/��n2 ���M�E��I@j��w�r:0�����EgI���I{��st"{z�k��wK{g��&�p��ӕQ_*j4����X�^}�Q�ޅ�ϫ�zpwN�y���b���;�̃�ǍA�I=�\�8l.�$r����v~0��˞x�!m������;��E�弤��h�w��$��׭9�v���Wt��Bc�oD��]>l����}�ԋ��Β�8(d� ����q��}G
�K�-;s�C.ą:�Y��B����Α���w{��~��D�\��ڗ�E�B���	�����J�3���g!�6��<٬9��+i1'��[;^VL ��Ov�?��=��Y���'�}�ɺ����r���#�E�`=��\��)����z��]*[a����~�*2&O�JQ�.�K$����O^>���L�2�(�`jS�Z�+�h�+�7<�����\��p������Zu���$�9ʼ��6����>FvO�r��v�=�Z�0U��]�
�,��7x�4+��Mv!<\��A.��N�Y��PO����8uIٿ>�%{�X�����Τ�:Kú����b�L��	R��5�N�XꔳJ*ٻ�Z�R�tb�$4(S���gvB���+���j��'�8hq�Lhϼ7K(b�r�SK��,�V��$�=�}�-���E ä҇�bW?hA����,S#���"�8���M�{]��;�/ʔ��Nu�J_�nI�N�Z*�c`�iQ�jnw����G�m_�,��Y0�?�x�o7�_5!N�6�=ʈ3����LT��k��˖ܓ6pD�K&�n�dz7�̐��+�s�t���DsJ�9h��0�n��ٳ����Q�7j4tR`���=}I�^�$
��QҨ��l�{�]�}e����4�+�ax>�߾�ֲ�lm�p.##�.���;�h2f�Rbz����D�膴9w0Bir��/z7�MdQv�S�)ʺQ���'��˾��������\�v�~������1�|����Vt�s��Q7�_��8#B!O�����j��POO;qZeT����n^�ZSb[�tj&��@CL�b�R<������F����71�祁��w�,��}�V��.�-���kW[a,�ƣO/����:1��p:.��@}�j��Y�=s'��֘ȋ�\o?��t����{u5��F.�g��ZXL�z
����müX���O;���%%�ϩp�*�6/�@��1!2ؚ�0��e�����\���t&F�,��+�j��������M-�Dl�+WzK؏�f(�̳`�~k�d	�9�b�ű��yّ��
� ]�L�]x�[5�T��2&�Wr�"��cۿ�y1��,E����F��7�M�'(��{[7xήm4�ͦ`��rq���W˒_!RH�O�]�l�	���!]h� ���%ww3!X߁s8UVӮ��k�[�`#;Y��R�zv�15C0'�v���F�A�o6�$Sm���q�������K�,�f���}\��K)6a�f��m���Hh+��E��(�C����s�H\f >_U���8v��y���~o«���=�$Q�	͍�G /�q�$!:�a6�WUT��`1����	��B]*�VsjO3u�>Z��+���2����H*��g���c�I��id�a��vZ���T8���Ǚ�*�5��In��m���"k�5E%���<X|f�#���l
䝊vB�`7y��u��Y�Il��C9��8��W�TM�T�(��:�<��ol��뼤���*�*TCWs�F�-{:�����ML��������ɚʉ^OI����	(��][��`G�d /'��Q�����~�QFA�{�;3�m��#�sKuF�SQ��g!(�19&���kP䚟A�D�s�+r/$�n�҂���Z�^�H�3�٧J#��
T�u�eW�*�u���S����Y$:�ܾ���s5�@��k�TO�#���wܼ����{��Q]����#�9�Qe	�z�M��p�UgE���z�2�F������}X_�:��9��<{{Q|�c7JV�yd�,���+�����v��q�BY���nCw�X��?�0��q�D~ou�����tW�����i�6��eW�z53�N�\	���������ue�(.��yd���O�	Vq!�z���f56��4F*xd�4��N��4!��[B����I�m�O���D�B(���AQƺK3g�8C�����A�FO��}c[�:+�)�&FG�_)�0�����E�N�BT�o��$�3�P�h�sm��F��0C�w�D�3���٪G�K}��>�:����>��c*�H�nJ���\����C x�BV��zݪ�=�� A�|6�uj젙�b�v����O�S��K֧y���lT�y�lp��d�l�����}=C�Gf��k�����M��PP��)�T����u���/s�C
͸��J��k-h�W�k���-h��Јul0�]���bf]��"{L����2MґS� ��k	�(#��H�@�#��Q����p�UP��a�<���M.߈�;��{=WW��N�L���oT�E$z�ƮF5_E^? ~3�Ǔu ���+��~}ݼW1J�F!��Zp�mZ�(4��9Tg+��smn�p�H,�/
R_�=s�kJb�幂r�"���fT�H
�����(l��]�����R��˻ut�@�{t�]Z�ɡ_+n滛����k���A���� ���_����6>�R�uhi��rqV��#f�so�{��ij���#2::&�	�f�}W������:��S-��ۦ�L.$����Y���dY�����(��@�D�p���P�P����h���ʖz�0rq�h�d ���ɯ5��+���X�F�(�#Y��X�au>E\H#H8�4��1<g������T).y4���2C'���&u�o�	K�M�,DXj6�����;ԑ]�g5�L(�OF�qd�c�L���9����B⯾|m)-�ZW�%&d�^�ܴ�EX3�ޕh`�]�-yMvB9��M�M�� kCHx�_b/�	f��~ĭ��sGnZn�U��h_rO��^�@��s�Uw�mi	e*`y���|B}�q�l^����G�Z�����*��7�u��[>���3�xd.�=��/<�3�Ρ���Mx��7��;��η)#z���'��<��]��� �z۷�>��<�U�#�m��rl@im��b��>���;}������H��{X`% ߰<+m!&\���)c7ܢp�������^	���\N-�G�H���Xˏ�j1sK�VD������d��	gܨ�$j�Ke29-gx3�g�/��\�W� ���p��3�XN�|u�3g����V��=#D���}I�Ӻ��Q��� �J���e�qE�MBȺj�}Ӛ�%|��Rg��*đLj��&�</�~C@�ґi�y�/�@g""қU�#:�riY�P_.�y�c:�N���Ue���B�;�$*z�kȁ���g�����qW���bZI�ω fII��K���۪�N#�C���T�$目փa�g�<Lx=5,R����[����|�*��x~Υ�5&�*ȃ�I9������T����K��-�P?H�[{��$ky�D^�V����`�§9�m��,�}Sx M�	��[�=	Ӣ�{��P�\�w}7k���^k���޳�L�hO���E��r�h$�8��������߈E���v���p}�b#c8%i�_���� ��:����.�Ի��?���3P\�[��k���=�<X4Vf������3[��׉͞P��bT,�S	w-�E�<��#��-��W�]�^K�4>�X'ʕ�u��)��B�{�;/"s&��v�1y&*��2�U�a�
�w$�-�>�jK��ZѲ���Mi'����LhC�z$�3��?������6��O�"��3Z47��������xS�{O���M�8�*�A�����4�;`�d+&��T� 2��z�L���bY�~*����e�aգ�fD��?��)�`�DE�������t+F⡺�����n�8�?Q�D'�1��0��}�6d�n��u��� �EZ����]_�E�6��BdM�X�Y��Z���n6##��s��D�u�[Αԣ��I��>����7�.� tO�s'���|l�B�2&�(_�Pp@�	0�#�wA�V&A���o�#_ekRqf8g vOGy�۶J�����86f�F+�N[�c�^��Gʹ�z��3
���ԛ�����-N=u��Ҙ��$�]���9���xg4BSz^e���cH�G|�?!d��>,h�@�%����ޖBZ=hL�%����r\��Q\��ݐ)�}@�˗ߴ��JԱM�cY)@�X�kؐ��t[?�YZ�ƫ��|���p��s�7�T�q��ym�����xFbZ���|RQ'�_t@��.^��LKT����t�N�n��"��}4�U�|*A�ǔ�0(� �@����h��ߐ|�R�}5�I�+���h`�/��R>~��-�f%A_��SyH�IM���\ъU��R캲����!Y�T!��̚����_�ϱ��>�a�j�[��[�ŧ�ܛg�;l�:FcޅW�������Q}�gq>�7�¨�x�/��K�G�;l�_mX��N\l�e6�g��吨�BU��җi���ug�s0��[��!	�o{�g��rM��Gs*D��\ܚ�������\<�ֽ;�㿸qbd�E�L>j�U��N�<^̏�[�m�qb�:�+XҼ�=U�����[	��$�7WI�0�U�����<�m
ϵ�l�;����@���B�ĳ_�}��/?�WB���G��O.�����������-<d�C�vu��;��<�jC.v�"{�3he������s_��C�;C�s�䏞��Ұٰ¸��1�P�����D��?"�_����c�5 �t~�$�TG!�2Q�E>@��O0|�^P��fSd��0�A�'ţ�߈v�4	�,{�\��<�t��*-2���`���Ԙƾ#�m�[� /#yĻ�{6��ȳ�@sKʾ��/O�S��>�C�6�6]��e�^�/�L~��/��������}������l�O��S�"��F�(<�%�zM7EݗV�����ɐb���-r,����3wF����>��+dU�9(.'E>��y��R%Gܚ��P�F\�5-;X)m��k�?�Fmy��ڟwt���D0��!%����a0M�_X?Xv�\_ SF�d�l��&��z"��1�L�����/^Qv����ؤ������F[�ח�:�� z��b�IK����^�̸4��W�`��XܩO��Mq��
��SmPG{�1'6��I���Ӊ,E�%ܭ�(e����=�I�^_�n=Y��O�s@�ԫQ�W�P˔R��=
=ጐQ�� ���/�ݢw�b�^]S��X҆a��X�� $D/&�\�wU��r�S��ǽH{؃�R�/D��49�s��[��2��D�@f�� ��e�q9k���E�P$	Z*�S�3���!u�8;v@Yu��G�H?�7"�P�v8o��:S%!�����n�u8�ʕ�8�]�2�ӟ���V2;H5 �yN+j�G�@�f��?)"f-(�Y�{�pCRSyh�*�r�(8U8)�k��(V���A���ܭ#�[���X�a�c���8'7��S�|>Uo��W�D����r����(�hGr�)+����w���a��bR�B@�O-��򔉻w����Z�D�a�:cEG)�(�����uJ�QKLne��>J���n�Ȥz���wˀ*�c~�6�h
�U��Y�\�m�^��ƯL��h���p�Gdd���S8"��F�YA& [�J�=��^���V�2n���K	ە���G�+�Qo�����8W̵�)w&��?r�B}ڦ]�(j��Z�����W�6�p��f<�=��Cn��!Rit�\��$�/s�Z�î����u<��������N)���cѪ��5�ڂ�--@�g�%k�9΂6Tܼgкw�bi�Lú��,K����گ)��I;�ICp������Yd�G�᰻�T+ �4ݣ'WT��-͏P�D�`��9s�v���he���I��9d`�Iv`T�/簽��i���q��wLjáK�������Ի:�Z���Q6�S�)ۨ�;[���*Ǌ��|��2M%��Q0��\<��3^6�Sa�!�Y�D�Jȥ����?E�(9΍�B:�s��uJ��]���z�f��gUn�b���4͖�1�W7����1��VY��%֗��8����v�?;k����>/"vƻ���P��	C������pw8OTV����#����Zd�������j���������/d�~.$�`� �ƴ5��5�}�|� <�CR�e�Oot�a��ꉐ������:J��Ns^̄e�~���̐��j1��5�?J9X��0�]��BO]���Z��QƩ��j�� �5�?絶R8�Ʈ�$Or�����U:~%�B"����h��J8�шa��G��)�8�`�ci��u@O��{��p�p��:6=d��k�H��<��YIO���]�E]�,S@�s	��w'�V��7��κH��Y�^������=T���� �t2�A�^ƺ �ao
8�$�s�7f� �^�\`�k�n���o �]�D���<�-���P�i��v�������l���өLJ ��o<j3����v���R�;����I"��k��]k�{�{�{\>w�[�/����\-��	5Q
G�ef`�o?e��[C�� �IB�+=�MmNJ��O�0&���AOM0�Q�'��SV�[G�sq덏c��c�hb�*E�q��Q
~(���|�P���}� �S��e�z���uA:$$Va�\���0I(�۞����WMq�����:��M�������~�:Ċ�{�r�ט]��C} J��$Ip^�^3?�LPM��\y$NOы� �����CqL6���bN��e�~r����O������jZ���ā� ��,��G ?*E�,�$�F0���d9W�j�Z�?.�����S��W�{��d5�5���I"�{aҩs��=��}z�� ��L���#���_zYr���|���0�C&n�ϱ*����~'���4��ԅIBM���X>uč�鑶"Y���v�dy�nZ�jŜh����p�N^ �7�K� ���YM�,F�="VX�4f�>��e��K��Lg�[������qЩGa��O3�m1eC�`�z�w��;^ē#���'� D��o�7��U��ɚ������QM�n�p��S-ṟ�s[�Ax)!�g�{�	[�
��x9�~_Y�����U:�J�bb���?����ޛ��[P�S�&�=��^��!a�@8ڿB��N����S c�*Ye�wH��sX.�U���u��(X��WH��R�!p�"݈!5�ܹ	��u��H{O^ɳ�Vؔ)UAV������y`�a&��ɒ����x�R�&�l���C�葞z�)ֱf$4��ɤE�:�J�Y����FtR2=Ox��f|[�w��į��74�Ј�|Տ1�4@���wV>Գ�Y�L��o�
ks���Lמ�<\�R��b�H�i�#���t���w5��6�EO-���tgp):w��t�P~�M�o��D
F�5���X�A�of�5o���@�����)��ѫ��,�s���FN�y���׭�3�R�ڕO#q/&�bM�TK=f��.�,��H�  :m=rh���R�$ �u�E�����tuNu��Y�*�O�dOtz���F��Yn��%K�O�'R�vb�_�6GBH��F?oӴ$m����^�ᨉ�_g���Z�7�&�#^�Y'�.���)�������_��=V&� �I
[ߝ�;{n%�-�񔤊���y�ȍwB�NS�l3L���e����F՟`54߽��4���X�\^�Ð�=�&.�Մ���{'���v��� ���@10$;�Z����� LD��38At��ns�������$P�	����^� �_���񿉞�Oq[���e����C:X��1�*Hd ����xF$ k�gQ�l�!�V���G�Nw�D3^Jc9�0A�A�]�A����|��)�%��f�{�.܍��|�F�OR���^f�Q=`�w3%��m,c,ig6kzO7��.�pT
,d!Llf0�N09�Z�����(b���m������0�{�fl6\�YUG[Im#���B
�$�\Z��7��_��׸0��O�A7��ۃs*��dJ�����L�Fu�I�7ud��|�B���c=�b�G�
?���=�-R`�Ё�-��&�=��*ӑ���!O�Q�V�t�{�;�.�N(R�d�q�� %?�$�=�J|U[�*�b��J(eȮyQ�yM ��ǡ��
����J1�MdT3-~�}��a}�֍�\s�d��ﹶ����7`�8Z�{3�Z.�8с�걓<�
������Cxyv_]$;�����{� ?o{;�0��:�k���O�0"���k���:�V0�l��V��j�_,)S$~쨒�I`�p��Bst}�6E��*�f������j$� P*(W��:$��pm�72�x��Y�^.I����#\3��t���/0�����H�nfdQ\^r8�qqB!,�Y;�;�Lࡂ���ɥ���g��K�F���P��{ �ܺ������tP�-�{��^J���7�2	Ҽi�F��ŉp�5��8,��3��/d�ֶ�oi������9Go��A�^Ԯ����;.�����&�����Sj�b�E_�Q{�F�TO�d�N����ݚ�'�P�{]L�����o!�m��Љ��*Ѕi)2�!%Q�@A)�N��ɼ��e�ɐ�g�y�`�����ߛqi!�"���(c����C(�v񻳍�4;�0Ùi*́S^�J��Lż�b�W+ϣ(�R������f�P�������'Z��X��q�,އPޅ/��``8��rA�HWaQ�3Yi��M�˵�H��c�Z�]���M��H�6�v�*>Dza��\�L��ԩD:���`yDH����.e��z��+�ʣ�������R;��28����е�Н�b��KC��fc��,뱽���������7V�ۍ����h�q�t��ڄ�nB&Ow��Im6�����68���m���R��؉a�z\�n����٘�^�+RCXli����s�Gr ���"�	|�t�:�C�=cM�jǶn�/?�.����ڭ���T�4Kb��2/���\�q4�\wQ����B��jS�/X���ET�D�CEF��NԪ�[a�E�t�� ��C(i��Y�>q�����Z��jO%��W�<m�U!��5";���#�ч1s�2q�g�Q��,;sRi��UԿ���b�[ͻ���'�P_�b����T����muso����J��I�iUHi_$5&��SY�3S|Y��o���jn̄cf)~˥O���0i75�E��*[�l�X�}4o��wi�1b��0{��m�̩iN���5j�òv:D���c�I��ZGj������u�x{R]'U:���(��&z}M��%MI�L+{4)9��RvQ[B@m�T�[�o%��|�!��a��6���}�?�Ƥ�|0����.+\�_OJ���_gw��h#}3vpK�';��(�6�����I�&�~y^�42�~l���e��yu��2�33�^�~�:�E��!��H+��E 9bM���f�8�g�G�uccB u��r搕O�y�Ҵ_o�,��q���	3�lUM6w�|�x��;"�-]�2ڱ�v�lj5���=G;I7��i2v$S�� ���.Y=�[���Xm��^�����3��?��M���O��-�#9re�z������R�ʑ1�ҀM���{�i	:�%�F�OX����p�B�Kl������V�SE⮷�����YVިCCn���	4�`��S�����G��MI�:���-t�+��Y��\8X�+H��qC>C�z-��#��G55;p5����QD�QF>�}I
ڎfW�Kܴ״�0��7������J.�*�G�"'��JIʢ(v��	��E	�����*	-=���yYN:��s�P�^�n�������չ�%k�s�Ì��8Mp�jIj��� IG��otc��������}'{����C�%��<[���h2\	B(��Ƅ�+t���>Y.��3�>��|�[��4��@�j����K/�=���M|����ҹ�ђM��aͱC�-<��Q�ew��	�������D掇!1��c־�/Q#�t;䪃�8C?C�4X�+����=$f��Í1`<z�������p�����ˡ��/�\R�YWh��%?z%[�Q�;�3��X=���ː�3|��,Yх�b��*w�T
[�D�����P\5B��fZg���}�y]��N��o���FC�J�%E�pS�;m��Tė����J�{J��D8�P3C�<�(�p��| �)Yy.��V)�H
?���e6]J���#P�q��2`轼ve�Mf�~yZ<�s��6�g���{	Cr9N����Q�Y6"�5t,o��r���1}�
ʔZ&+��0i�x��S��C�xMYTu�d��`��(P+�b���?R�e�L���x�0Xr�d(��8P'�������{���j�I�y�Y+C��M�k7�9}XP2�t�G��e������B�i���-̭�\I�8M�	~�������&�i�f� �mE%VU�=�}Z**�#��q)H7����/~)�������}��#�XGA(*���k�G<�9F�T���x���x2�
mE{:��<D�%��Ȼ�Y�4.Q�Y�Pe�����7�/�5-����lG ��}���z��f�r�\F�'W����}[-�e�:�NS֩T9o3�����L#ux�:���-^�
 $��頜\�9-\р��ũȢ/����?�W��27�Bh��릴�"������?u�!R�"�!�"r���S�qZ�ضTm�p�.����\�r4B���B(�����#x��w����Ö\�z���Wq�%��`�t��~nbyB��!��)�AE�֮5��(@G��jqe�7_�;���)��`�y1�j�$WF������Ulձ'�}�Z���G�e�TJ��8%M���ۢ�G�a�=�yz%WAjIh�j|m��քT|��U�T����ˣ����9����b��JB%�Bͷ]sf�4��d�ɝKZYU�7�������fb�oi"�ٕ�Î�:�6)cd����K��<����@g��ȟ��1��á��YP�-я�ol�j{%�ha�M
��:l��/�̡R��:���F��B�k��:!@�+'k��=б��"��c�s��� + ��i ���W���
'? syr<������ykj:��r�n��3�&�:�rM<IV�uO)�3#�J���PygS���H<ݑ�&)fM.}�Z�|-E���h��u��P ޤ1 qA&��Ӹ�Cw�Uf@�ι1!4r9�:�hP�n��2=��M�e��Jfo�h�kߝ���j{��0Zh[@�ւHf�!���M�$I�'t{1��$J����m�_�gQ���4>�����}���_6�h��k�Ra��7�mlAr��Ջ.;�Tl����hv�L�~�\�Z����$���JfƔ�D5�,K�r<�#�E��?�<��N�Ւ4�,W��͌V�	���p�3m�y3!�H����_�`�F�:�Z��%R�I5-�7`g��V�q���?	Y�9[B� a��We�=4'�B͓���U�b���e)�޹|�C�FI��vHi�N�;��-4=ս��]I*>�f�v
���t|�=�ާ��V?�7l��7Ɣ���؏Tu���axaKP���:ʂ�l�ˌK���&eqӮ9%�,�:�C��u�,�)6R�tI�� �l��mf\��)���3���N'd���藿�����=-����gg�	����11�츠�w�>7׹����|���=lf�=F�k���t�0�|.x�8�[F����a�^�#w�%�OWfa��p:̗��'����g��!��:�-:}ͺ�mG�-=ĹS�z�^��%dt�h�*�s�����
�َ�4��Ӈ��.�x��^�$�P>�ysScq ơlϽ!02k#���ΚoڸY�3�����(����]@�V�d�'k��a�*�Hz��J��4)�����1@�rĻ z>An����#4��G�<���'�;Z�"SU�8���T����|Y����lf����"����ܲ�bȱZz=����\���B�����a8�+r��z]�᪊�Uee ͻ�ꇻ���k5r ��߄p������ �A���;����qJ��Z���D�y��ȆJ���߻k�jqLB�Z	;[q��U�߲|)i	�T%�h���C�r�Q��{�zӠ�P)�y���/1G��#���d�6M�j|9@��~�������Fc.W9Z��#�o	����K{��p�,_RYG[�)�v@NJ!�S���'U����G�;�%���)�/��:��
<�2T�D@)��+�N�p�̋�U����8@⨿?���)I������є�1�ǧ�������l����.���0�P�Rf�;Mh�5��T�������N/ A�>�҄�{���踌oi݀bW
mp�3�iq<U��X��Q����u�*r���A��K�=�*�?�eu�<�7���k�U$:h�/��8��#���n`} :�lO?fEZ5h�H�HO��d}i�-��'�����ɛ�~�C�[7��"�bdG��B�%���j�W�JM�� ��@���YB��^��Xe��gi�<����ˀ�떬��8�ikgT3���ռZ��u����e3 �2����<�n ��;���d��0�L���bMe@v���EږD��Z&�����	�ǩ����w�BXLItv�����7fX�G�*}���rg�B��[)Q'����/����g�kYT��w�N�+��yuw�e	����t��(<MbX��*e�xwVa屇��69�%�M����N+��� |K5���3T��Y����)�� 
XB�W<Oّ�Ƥ�Ѱ�\�CZ��w��1(�w�u�f��,�e���\Q����Os k�<�u�q%Lj*��!�! ���nJWs���وF԰4���;\?�����*~��a!���y�P�\��%8�"��.������ݗ_�بa�HX�\���~}^DH*��T�պ�فiPB
�
��V�U��������?>�Fs+�# ���C%U�6ي~|��I|���m�m�0�{�3����*�Y�"|~8�2	��Y��6��ﾕA#NN����$�љ{N�s�q������ ���m���: ߘg@�������9��2O��&����G�@1kFJ��M+j2�����aN�w[\�0�T�&[�Z%M�EEX�C�:��8��!��A#��Κ�kW|*�U|����ick���`����������[���Y߅0/䰍��K�o�
�+�����1*�:\��e��!��'��(RuXe�)kʇ¿Q hɥ��E�ㄡ/����n|\�� ���� >#�T�p�V�fb -y!��Ȭ��X�A�9�rIa×n>.���i��J�]bБ�轄߱b�>x���
a��<���UuH��/Ӷ cmR�؝�q�4����p~����܆������f��;y� K��lq�Â{,vC!�*Z�-�8?�e��ޥ��ϴ_�(�J��a���F��������2[�a�Av���� ��N��q1���b:��-�ʺS�x��