��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�xP89�f�`P>}�~���s��E~���6�OO��ih3bd�M�,?�='�~$>.�]t�����,�LZ����O���\�����p��M%c]�nuʏ]&�6�����lJR�]%�8�$)�?��b�5��{Cw(�D���R�H�ۻȃM����X�>���3�b�r��=�ng}�2�����vKFt�O�U� �@�EzH�4��fB���_w R�6O-D,���1�����������R%>$��&\=�{���@'Z��h�9+��1p�R����u��p��l�W��0����Z\�_�l��c�4?VU��L���vl0�^��7$~6�F�,~�%���ߘa��qƛ���Z�.8��@�-����?��BH"��bEi�)9-�̶Y���P\߅�IV)���h��98�W�C�j�Y
�y���&+BI��(���DUHA��>O�%�LA}�Lbe��=�����}x�ʖ�ɳ�,F�ri�{e�Q��>+�ly�����vN�����?�uU��9��k�{��?�p���s�����5��Q@?�m!L�
�a��A��x���ʳ�y�>ƟqXpD�Z�b��5�s�`B��7ƿ����<*�g',�=Ԏ`?������p�N库?�vi�'~�,~�"����(=mxp���j�ņ��WX�R=��9����h�}��OႴ���+CO�n���nL�`��yOtd3���l^��]�:qgBM��An�iϚ��gJ�ը�=K�>��u�1_��n�:1V�?�� ���$��x8���c�㬑#�6�91BV�1�`Ԕ�E��i���rś���e���S�H���v�w��N�d�>��>��.5�K���,{��/�,3^D�B�h�;lh*�
d(^/�߀$�`�-2��,�s�W�d��4��laP�a��JS���*����߹��4��m�������X<�]�~ ���-s�)��ES%Q`�[|oo���iZD��к�	���n�ň0G=ZM9m&��� ��PM[� '���V�U�CU��q�Y\���>(w��P�^k'"���*��Yn��3ҝn�A`��^��P��^��[3}�9��	��8���h˚��d'��r�;A���F%����Xly�v��5O��)��D���u�w�x�
��ܕ�gN)t����aE9bb���S����m�[�i3�|2ٓ7(N�z��D�GG�������n��#��'���F�_g32ƙt?뤍8'�%��Ry�yf&E�'a@J��m����`S�M�'+�4��A�����qb�b$�_�럻+��2�o~��3�Oxe�$߹�"�k�I�d�i��g1����e�����-�Ms�]#_+!	�U�6��ߪ��z�8
`x{FE߭
����[[�D�g>HM��+35;��բw�Q|�M�_4{z�E6>�ʁ��ѐ�,MX �N��x�C�ڙ��׫���ќ�~�+vז4L�d*M�pEv)�=b��>\���ڬu>/<�������%ߒ0 ̔LP�Α5�9��>�rXՙ ��s.RB�,�&5X�/n���u��/��f�qP� (�t֫��V~�٥i��ۓ�������eW3R�|L���z6�^�2���������S�pUȚ�5(�i�����K�n-��m����7K���5��Qi#�W��8�5z�ڞ�xq/��h2C�������;!�J�ĳ��^�z���h"q�/v������j��L�7]�:������$�;ЦR,M9����|��{>��}��k�h��発#��5����EEqۂ5]2h���>����`e頻�
�x���D��>iR"\15�p �џF(������yoZ���)&^�5�