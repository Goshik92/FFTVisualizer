��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]�{I�O%m#�9(�@5�g̼q����.��q��dN3S1F�j��%�Qs�H�:��f�w���>I[t���J4���iꃝ���E�ύ�J%u�1/�LqQ�Y"=��s.���u�k�M��'�⺓)��z{�)Ƭ|�L�P)@�~X���I}����h��t�*����4���d�2C0�Xn��vbF�	���,�[�a�Kd��/t�ĵ�E�i/nH׌ �nP���F�l�Y��h:����1K[o}ŧ���u��f��x��3h����	�~�ם����݌{��� �X�g|�G���c�$-�pI�ݿ�~��`��d��ß��iK`���g�⸋�P����ղ ���F|�<�3/{�;�L���u��~AKD�����)ng�����J=؂��(����@z2�q�s.�ـ��"�GE>J����tc�e��ىb�5�Zո�%�����aX&�J)�*Y��zg�y �~�l##�A�Y,�a
E~�5��T��2n���52���LH��!Q�#��t^��3���H��qZ��J5(޷);i�%���IP���gH���ɸ,4)�c��[���?��|T$A0!�j�b�v�u*0
E؅��ND#n-��i�b��p��*H�]`(�����V�*h�0�u�q�b�Ȣ��i�L�3��	�4�����o�P��;���w��� �G�;��R��Tc`Ȍ5��%�a�'t�񪬚��? �2�I�qas˽�l7�9��y�$��7�#CΓV]{l3M-���_���Vy{h��̼F��e����V(���"l���M�)�£�7/AA!{��r�n��MLT�
�|�7̭7�,P%ǅ���qp��s��#�+X2W�Pt�3
'V/t�`�i]^)�nWbS{���K!����:Κ�.X�Er~�~���&.��o!׍lbwV�!����m��"���b�����.�O(�J�%�HD��`��&:#�J��v3c�]7{Q��	�O����������8hDSVM�9���%�ooV;�#Yw���qEN�}-jBet`��oY_�{Ǫ^J�O�d��I�ã���d�db�/����8]��M��/ݏ,�7�k��*�C�`���k�@#��Tb)S�j6]U��A���i��F�K��F��������5if�ƛS��B�&qh;FA�^'�8��+:*�3�F(v��h!ބ2wڸoC��m��Z�*���*\�.ݺ�cc�J�.�*h��?U�1���H9@��R�f����M���I�4�M�sAV���8���W'@�7����r����s	ŭ��,YB��]�]�R��ҦZ��zF�R�2�U?��ō��.�q�T��,�rBm{��Ð��4'��KO}AIz���p�v��{��K҆&_-���;�����"���~f�I<�����\*T�^?>��2���쫏R��P-�2nn
�'_rڳ���ܘ�!Yg�?)���>)�w�]���;������(ĺ*�>�+�@�3�S�0h��`
�H�q�W�X��l�g\��p�O4=d��C��T<,M�?w��N�w��v$�rE7������9'^	�a�L�S�_:	;��`/�`TO�3��`���H"�*����Y'���:"(J�a	 �c!����a�;����?ī=�_�Ù���� ��Θ�9E�kWcē�?�#���r��j�s_��]r�_b1 9�;����?o1*L�>���
�T벢�����Mr�b�Y�IvM��w/S�n����ԟ��=g�rc����Ǜ|ۆ�t#U�x3z�.���d�>$��5�K C�>�~�~�:Y�V^�bq��J݆�w�{����)I�LEq�*�5����C���'H�qBa<ua��Sɶ�A��!�xllÙ���xo{ ��#�L�g��%9��\�3��(�:R����sL_�.�y�r���
�/�P>��B=��x m�53�th�5*�&�9�ڂ�v�f�H�6��ᗪ��g�@��x�x�X���qf2n�d����1�5v�>�7�!0�B��粬?L�y��ւS�z��E��b�����@�I�#��j� sD��Ў�w�ܶ�(<�����b��A��4B���t(�o�P[�g�5���.,��ZВ�DVڛ���F��>[нW�Qx�!P���iX؍��(�'�����c�u6��� ~[�=#��B2�e-YT?�ͭ)��j�D�T)�)V��S�IϏ3y�`�Ȯ��J�|n����pݗ~���ϣ��`���LK ��[��DB=Nj^3�����|5��|����_��}��ٔEe�O�]���߅��?��������=�爁E�f�M������s�-�����ڡ�wx{� 
0 ��h
�Tx�ɞ��9�����N���Ӵ*)"X����4�Z	q.D6���%Rc�q�J��N���_�ŵ�W��i�h%D�(s|z�Ewdˌ�S{�ǂ�a>yG�wU����:	��79���YX��{�ɸ����	N��Sh\��;�����j_�Ȋ^J�r!G�~�86!fr�yr#��շr���򒉿`|�$CZ��y�DP�϶�i���S,�D�37���zV��oT[��yt9=� 3ewx�M�fd��E��G�ܙ ��_��-g�X���%D��gݭ��Gٔ`9��j�0���uz�I���/��];Rl6C�����'^�e���K3H'xY��hc=	q�ʯY���Zߖ�"
v���e�S��z؇1�������o����VϚr�z����ֽ���g��x69�~�?�� ��� Lf��᭙�:��B?y�+�
 �I}�ip��]��K1�Oc���?�y* =�)y�m���:�zS��w"=�k��z���O}F��`��h����	��y7���Z�I����tR2,��V��$���`Q�dL)l���=	8J�a80c�8��q1�vT�*9+cQF�4�����\9���t#ƁV=w��V���D�E��*'�ΐRwߴ�`{^��������t�8aHA�*c����������Fs�j�'��#͢��9?$�O`~����Bƹ�_�jut�6ql����E��bO��}�T�F��k�M��0(�Vp��k&��E��u���R=�+:�:�ź ۷��1)CPC��`V�O�n =ѥ��{���E��Z5����� �L��̌�ia���ϕd����>��4�*򳙪�$�Ğ�#���A^1��%c����߇��
(45�D1���`p�Y����A�}d���p����f��L ���&�稞�n�����]�iHMC�m�B#r	�O���e�՝�ڕ�!��_^�0�v�Uk�d�'��]	�	�`k�X��]�KU8���ޓ�F�z����k�c4�{ݑ!`	���o�~��*�:ȔER�(��?-h�裄��|����ĸ��}�}���0 ���]0ׅ�5~���`�4C���dSM�SYv?�m-��F�c���N	�P[0Ns�\������h�`z_����L�Ȩ�w���=�I������S;Ա������1�KdS�4L��(�0s���=��7T��m�C�f������^H�j�i�ic��.���OXrDC��k�_|��ۣ��)0����b}���0��*ʀ}��S�t��t��e'l#r¤��Q�cJxT;V2���!g$�W%�@��Ƹ���'N0����,h���D�Q襙{T��g6y�,��аH��,otmO�L�2�`r+ւnvܺ�k���C����9�m�b���b�L��Kdw�Q��Z�����)�K�In�jG ?�
��qJ��������:������li�l�-~��j���Dl&��zI�U!wp�GfIܡv����6-�.�j�1�}��Q��4�8�E�s?c�����A=��%��o�]|��W L�\�{�1 x	R�O�Tz�s�p!�~	���M^1���up��٪�"��B�dɊ�-���݀��E�3[t���SW�T��EG}2�{T?�^�#��_��чp�*���ט��r��T�����+ӟ�i ��h&Qt;��X�Cq���C��̙�����19g!0��A[���Q�ug���;/[�7�$d����lD/<\&��8o��V����@�@jy�R3˝��e�8��V�d����)��Bǡ�����!_=2ܘ�T�n�&ZZ܄)�(Y��Ӥ+�� �u�/:��Iz{vX��M����k?I50D�
v˖�d��~���ִS�\ڊ���*��H��t�\3{���[��#T��p	c��H4:����~�S_YH�����^�L�mg����g^U��S��u5���/s��7��Ԫ7Է�B��y�����=�Fr�Z5M����},`+PGJ���$�{����|?K3'T�FN�/����Z�1�T����*��π֬����/H}1����t���4�ܷ=����wZ���o��E�SG] <[x8g��~�l;���zU3�c���^!���<U�����|0��o7��ڷ�0;BO/�Ԧ�L|	��B�98mjk�����s���y,���D��n'j9@4���&��"��UTK����qW�6��R�'�~BGC�����ٯ�h*,�lk��c�]�U�F�og�X~�����| $���(��r6+���[�R{�_y(>�W���I�"+��|}��7�+��8�@��a��y}l�eW�����č�N��uo��(��;������,�%J��c�Z�1kO}�˥���Ն�{�
W"6f�}�	Q̐?eY�c���%sD���j�D��܂g8W����3�^��NՕx�ګDc���2�9}M�q��	��X_P|e[2>0!�Y��c��FD����t~^i 3������?��̙'H)�Q*�:.CZ�겣����$�?��� <qN՘��=3V�{2���T�\����U��r��zd��/����HR�/���|
f�>�*?�LI�ٓ7F�S?��	=��U[����k��<�����N��0-?�u~�G�}��F�i���<�������}��h�y[����^Q,v1��_�0���Vc�?��K���]탈J�l�EHn��t�ɸd ������}�;�'^��RN��gKj�Cp�ѭ1A�ߏ��:�)o�@��[]��H�Ø�����b['+{�M�@����ml�A��\}@�!�~e��md�B�O���I�*��Vk�Ln*4|Xp�:&H!�r�:�A_P<��0nq�cXë<L�?���:'1v�)�6�%�S �=����}`0�E���a���͎t�$�I~U�2.�i���!;Y`�ا+�bˠ��4�6�y����=�j��|<��ah9�4J�֡a��)g���~�*�L.������&���	��;Z=��^p���
�ϋY(��x�^��/�=����\����l`%\��\�m���n�Q:b�<���:�>�~�KH��Mv�o�2��v[� ���P��U�m��.����
�����x�P���;S�ǒa�͎/�l�(j��1�(������3��ό�$)�f�w�+�@B���!���m͙�Ba��4�[�������Y����G�b��m���?�
�y������t��|����1�e������aPq��E�)�9C��e�J�ǀ>�R�a��QV���+����U�.�v�b��va���/gP���og�������O���Hԅ+�3ѽ��>�~6��ZKVԤ��k�cI��R8�^)c ٖϗ�5��$�K 3�h��R�4c���ڨ�$?����e56��@�}bܑ���ppɝ�I�����e��zC �ԑ�~���{Cp7@~ʚ紆>mH_�T"yׯ6`X����݉0qe**笆Y]=Z]�]:F�n^mZ��}�Z��ĝ����A����]>��
�" ��\L�B�/P����0q~
Gi9Z�>�?ߜȐ)C�`k_-{*�:��CF}hګ��tb�/�33��XE�&}���?kȪ��ʾ� N�/�	^����dyQT�G���j=[�Pf+���7qt�0�:���}�i=p(�{�^�NWX����0����奆�$�h���1	C�;��^���$���v�{�#��H`���=[��7nk5{D�<hw�A��h�����h�Y�z�g�_��� Y� �^I4�� h\5"Ea�nfm���`��!����G���Z�d�K�t�rZ ��d�-p0�5��E���%6�L�p}B��������I֏V��I�,s$A��Ś�"
��V�6͵ֱ��}:/�x{��E���|����F�C��uh����i���ˀp y�L�g�d�/���y��|�����\���H�tu-ț�=uqW�o�t���c�e�?ŰM���z���#%�m<;]E�Ij��lD/,=Z0�\Qh!p�Ro�_����RCh�1r-�sZ+j�	���-�+iY5�:s;G[�#�T�[\Xx��m�>���=���5���i( �K�ɥ�&�s>�!��I����}����"�d�ui`��c��X,���/��3�e"[�b�-�Ǎh���<H������� �.�qs��	��
�e"���(�. ����DJ���H�~�EF��V0��&��m��*�ON��mO���&��a �ψzX83m��<�U��x��{	�
�U,1�&�����@m'�9�}H���u%�3]<�WtNr��cC�ߦ�!h�lA+`v ���Yz���ކ� .�MH��>do�����[�8#�^��|]3
6��슿�iC�(��b'�Wسюi��[+���l�8��N.�����G�� ,��W[�#�v�e�=Y+�3qz��߶k��i�z���׮i��2��ÖH��"�ԏ��a9���שc~�Ӝ��e���[��u��Y��Z9�uY/x�V�T��\-����{1�v�3H�Q�n�J)a8�B�t}Ѿ�2;iJ�n���ȌpK�J�(bʡ�"�����@2�f��
������E�Jl� �yv7[5'$OZs-)A`��O+D�Q��X	���.{N������z�jms���������-�-Ҧ�$׉�&����@w�{��]�������vjð����`%���E��P-�y�� l�d�ũ�D�L��n�5b�-M]|�2̴݉WO���:��~Q�v�0�����&^]e�w�ׇ�G��)$LB�����`p��`�/���Tw�G�>'��q}��;@����{�)Sv�D���e�4�U�{8��&p�r����QzP�{
L�o:���d��ѵ��0�葮� n�c^��d�7廁8ݍ��a*��]H�a��z
�����Ja�,�X��窃d�i6X)JX3�e�h4�6�x��������poFl��Ү�iG|/���oz\o��3/�=�Q�A�ϡ�S'\&Q��!�	_qεHT�GZɠN�5&Z3~�ΦB"$�;���::R�����¥:(�{��2����̝*��Q4��qI��ZgL	��&��UI�w����~� �g5�}#�=O-C�4�o��nB��7��wҳY	ƺ�!�:�|4Y��n��C�+���_�bQ�7�!J����k�7�2�}�7Y�ܪ�ri���G�f������;�l�\Y�~oh�FbN<�Z�Q�Eg�����l��~����^�Wa,�Ē���[���F}n�ލ��8���+L%�_{�
~�j*�_*���P��N�m@�������ԁ�0�ёx1��	��8гth.��$f'S��H��]�����藜@�����~��]�Y��H�u_&�c�À�h�K`���E���ֺ ��Y���n�	J%D�O~�@�Q$o�ߨ�,�r��=[����c�n�����vEz�4i�#-�p����N$�/������/����~�]�dݻ�Pހ�)Mg�s����}vD��xl����|HjQl|��C�|&-߀Q\\k��s"I�:�Uo��زRo]~�.[��XͱϾ�Siq���|{kŏ���Y>�r�� tc��2.(�����WQE?��5�����Ƶ�8��[�¢�p�h]s�����g���.gܓ\�*�҆�h���(;����,��V5�E��'g��E��A#�(_���%�J0����y6� ���+���i��܍�Itu� ��g�@�`�tݨ���,wqW/(9r"n�,��˝?��6%�ڰ&#����l�S$�����x����B� �
[?�N�h��Z�%�!�
o������9.݀z�I�T5�rÚI��b�"TҪ8\/cl5dfְ��\�9�g�YxP��j��VI���W+��|T�̕��.I�A������y#�g�>�_,<f���B�8�C��[>^.��\�R�"�D��J�I��k����v�{�S뫸�{�#W�P��߯��^���y�K�s�y���L�:I5!�	n����sX��􄞶[ؠ5tc��J<;Y�Giy�CdB���TOr/�E��kkŘ�R�r7P���	���d=�˺$�=���m�=bG	��xU�V&��(�X�O��T�_��_���P�d�BU.�a�ZQ�P"ic��焵�)bO����R���"s��d����bj&J�2&�5I��Kuu�N�Sa��'mb_�5[�v1Y(�bJ�g(�ׄ��ۡ�Y$g!�ߦ���)/7�u�t�k��2c�G%nV{����TC�Bo���D2���c&���y����d|�.��R�>?C�Y���`x��D���32��	��"���m̅M�KK\f�l�����M��F�Vi@��yv[̸�4����JC���)�r11n�o�n�@�a����=A��,]��%7X�⤢��?u�Q������w{r)ʿ�8h�ܐ=]�r T�����&���?�iW��Hn�z]�l�~�)�qZ(�ְ�8��<���F�7W�ȷ'R�
Q<`M�v��6�#��"[@����P-�Ժ���a���X�u��N4�>R�]C0������,�:�`�Nd�W��s�x8{4��w���Cq�ZDۖ9Q��qn�-�-���n\�-j?E�j���s!j�ʀ��Π�J� �
M��T�+8}��=���&G���s:�|��:���xsnH�
��:�oy3��FlN�Z+D��n�	�L1 x�{2d8<�Y�& ��I��*�p���rf�%U@ʔ`B����Vq��_��#���tR���z����I�ҡ|�R���,�̛x|���¼$\��z����>]���x~�B+ΓbJ���C����S4\ݨ��kR�%$g	��J�v/0��yĵ��±�>��,��.��@��je��I�w����H_ӥ���ˍ�`��A|��J�]�]`N�=`�<�7���ila6Z� WU$��jt
���Q�UsIn������Tj�oK(�
�g:T	f^�L'ʇt�M��<�3����1ʔ��wZOe��sRS:_���<�k��(�������^jfh�~��v��%ۤ�m�y꣩�<�E�lu��L�S����h��O���ֳ�ÀP��/����(�`�scşA���c����v�����O��h��wH�����O�q�]|%taoE�J����Ԧ�y�Ж�c��
[���G��2Hn�M����a�I�[`��h�K��{�:�o�Q+R&~Kz��]H�ԡ���u���dAɺz�!Q���,e���I�G�M6��IV��ȓ��:�>���v�S�r������Lޟ*д`� 3,+=P?�������G!�
�ze��<��$F�h[y���Sǁ�Nki�Aڸ��ɹm��;��\Դ��9;@�4�ʴ�� ������Vb͒s;�s,z�>�9I�em�O��N�JVtĳË�*;�"�Wz���!F�>��,�D�����❸�!�ibO�x4�\o)clwZ�f}��Z͙&��<X��'{�ɢ㱄���!:?��4�����E訶�s�;b�F��=j<n)��!�T�)���lP�*�c
#��" �Q��3�Ǯ���Y�鄂�M�+�Κ����}?ő'����8�D4O��� ĥ�ee�HpIE��7��[�؁<�^EkH�[�k�Ý6N�䀯)v���+13�+�~��$���E����6!�s��`#D$���i��Ʀ欆f��d��/�6;�w8P<�x� ���k�:
:�SVm���(t�ش��׍5MJ�7��Z�(5d'#�✼�����.�&�,�k���` �[�B�,j'y�b�.����D���LOd
��#�4b�W̍�Nʖ�E�Po=>�U�'��ASTo%rxOl+;�%�*cp�z����*h!����@�����D��=^pOH�i�p�<�:&��i�djV[ާ���-�ȁ|L5�/�0
��o >Bݕ��y�CR�,¢�?���MCs��"���`�iּ"iѸ�o�R�ДvjcϺi�O<������*���q��׎�˶��� k�$�s�)-?EC:�=Lb󘔄)���ql]z�p1A���/mIo|�V��Q'�t�J�$�P��J�d���T�(*�a%_��p�Lcl�Ԛ�v]��UZ/	cи�r����3�a�Yb�\�5
X�J�3ǰ�^ ���Uc���(��"B��*���{\��!�!��$-�K,��p��?��|{=r\0�(�pԠ?� (%�'����m!�^A�r(��B�W+b�{#e3!�o��by�\�{Ð�h�UQP�io��##w�E3�i~����JЖ�i"��(-%�Iek��U�\z���j�,|^߱���=n�����[���MJ��%:��Un�m a���ơ��
�k$�ܑ3�s�������z���0�L�q�ǿO�����M�����*������_���\`7��ɀN	��ݵ�n�� �}��M��B�`��ru�9�m͜~�5��v����Q��o�+��.L�8���!0��#Sܝc�(����/C���1���u���.��xgI���PJ��9k���N�ˏ�j��N׮R�9�^����V^��=�-��T����d����t��'��x����
I�q�m�L��N��/���z9�$�i���?W�#k�o��8��ʑ+I��bS�X�C��+`�S�wa[�Hi/U�ۊ��N��Eb��G����[ۭ|$9��	�3�I�/��a���"���"F���Z��s����A����$�NΪ"�*/D�|�x��A07c���q�������˫|�햲E�9݆��)�(O>�)�l�ĕ�f��*�'Q
�}p�u_Y�>ާ	{���>�z�Y=�+g*�D�8��,��R7�;ȕ�'<�m,S�q�^��m���9Tt���3�֓5�ܬ��t���;1��2�^�U�J�R�����33�S���Vv{H����ֹ�Qr�=���T׆�Ⱙ�P�S�C�(w���t�i�v�&�GYJBﾪ���E0���.���'�,�rh�*�GlL"�Ёb�/q���,jbIݜ��� ���Yݿ�����ːvM_%Dg�{����W�d�u�r����+Wy̟!��/��!	n�L$s�����DU8�uE�a�t['^G(���'s�i)~{WR4&n�IXR%��M�.�R���@�f�z�|u��_��|��D��STX��:9/��t�}�{P8�4M@�I}�p����o@�i~r��"nA��-���.�nL.'e�g.-����}�:wƯ��;���Qϭ.�oU���6���{@��C
W#`���v���nV�}f�3��]���iXpC�#�K�ʗ��JF"��~����-��������Td4�p�5��	�K��+.�]�+�ġ�R�[� �)A	�.�F���r�w> 
�UW9><��h��BpZ��z��^k�Yl����
���w�nd�)
��A��7�\�}���z4Q���E$'���3)WS;P%�<,��j�1���Ď�&bYPZg���� �Ny+�(/F^׌QX�$����ɖْ�q�z)O���D38G\�a�稱1(��P�h�#C���4���P�>�Nq�S���ٮX!fAg��r&?v�^b��ƅ�E�8k}��b��n�)����wѦ�_B�����Ƨ��D�Ja6[R������+����oj��c#��^���Ov;5�+���b�Z�[�%c2'��E�gv��/Z�� �J�]'�i�|����s�{R0xN[ap��I"��b'�0��=7F�j��#U�v3|蘏z�U�DX�ݵ�d=JG���ƭ���� �LWi�}-����R8o�������x�Њ�nyƙ�ӭ�SA���@��[A����=/�Aڂ=�\�rY~�[�>*��)�ET����t��`\�\PkymH&n���)�t�d���%	�W��!��st�]P�4ٹ����K\Y��;J��P���f��4�����b�|U�fvL��y5��N�Ц<)=ś�{��Hw^� v����X���Ҩc�^;|P�����A��kS���g?�f�>�.=E`,p���;�k�b/�Α��i)�s>?�� j���g!�wy/��S�tdr*bVIq�9��Ek�2�8������XΑ�=>1)�)q~c�{Z�WZ�#�Ōx��y7�k���k�2pI����'ܮIk�M� hl]�q�r��F+̻r-R���)nl��#�v�(�%Q[yI���yFJǁ�Y�y�]aa���*�T�P�}�0g �8S��PS���&o�J���XHx�����V"�U�ЕX
�~C�Lt/wX��Дe"�>Ef��]�4���Y��K,P9M����C�Ǉ>=��?�D���AS@�z�E>�Sk�7e�[���\.�{@�$B�t�|O��r�d*�x78�_�_�ܒ܈<�f�J�SY����Ey�⡄�zEIR���8����;i	�wK�������ِ��96ϼBFc��<5ͫ������_� A�ia�G�h�}�^Wښ�����%��9����l��`��E~^m�/�(��ZX�,H�$sv��z7슧��`�b����$'� �̀�
@(./��{�}�!l����l;0���1r��Y3gf�w�S٢ �I��."G��f(���ݴI"�}_�aiisA��[5�ɥ��+qt��`*��}�T����g���#�$E����2?P�y���T���Y�Ŗ��!����9��9��N��k��_��Of�G��Gq�Ԙ?L̰�A4�m�ttw fy�	
�؆S�>��/�r|ps��aV[����ꚢ$�@CH��w�jI�'I'O4k�55�48�ĎIfjs��L���(�� ��I�~�[����9#�c�
Y�[��x��� �� ���4jWZ]�]o�	<�Mͤ�b��ZA�Q�q^=�zM�;��nZ�y@��ߵ��]�}�+k�E*G8$�%f	���I4Oԭ�ǉN�V�����3eSY;ĸV�U��ĭ-��͗��9�uFjC��"�0.*�1�I����\��=�q [���=ә��#c�˱1{𼭛G]f;�7��_���9�}p/Bs�����g�3|ǅ�k��a����\�hi����լ.��*��~od���Q��X��b� n����v�4k��~Ufp�̛E�?�@H�}/���Os�'4:�Ӎ��M�����O'�3�y�`�j����g��<�?�,m��L��0JK��������ז�K�cf�G�*[��2��=�wTs���3N7�ȯ�B�@ѻ� ��q�ּ^�6��?��HwT�G�w^_�����c�TY�[�:T�!�B&M�O�v�PᲞG��6�\�>�w��t����{�8�X�44��kl�!4t�uMZq"y����	)(XN��0�]>iԦ�(�����I�֛��m����+��,��H��aɟc�K��&���=������T�X�����x�B���*�M\O��qZ��;�۾����׶G�p:��H$���D�^[�?dg���G��<�lT���+q�l���@��L(�W��" �=N�)as�J�rJME?�PucC�d�!5�����K�e��7Q�&��<��$w�~$��1�V��$��^�a�n�B�G«�m..�$րEQ����s�9��6��^�#c�V�6y/Z)����|�ex��Xs1�Nؿ�9۫�=q���|{b>ȅkj	�nC�����g�q9�0�z"�n.y՚6;J�����0_Uo*�v^��Ov>ح/.ժJx��)u>Y8#`C|�s��R����B?�$z�����^�Q[�Aq�i�#(�͞��a!жb�#L��f�vX|�}8��
��@��S��y�J~�+�]��r���.�Cõg`V�0c9��Z�|3����4E���Ͽ;���)�QD
��3����m�W��YP�@%����{qK�ZBb߄^�W.��KNy�n����uf�P'Ӎ�!UG�M��r�O|���d�z�E����\Y,�Yk����aO�t�zK�E��X�W[��wq�7��/��X��~��G�����:y�8��;rN#�6G@	����$��|<|h�����{:��#��B;w��W��nO�ɕم��o�"i��7��hF9�g4����<%��L0aK���e��p{��c�>b�8�0��{��
aN@ρ�P>Ľw�~���D7�37rq .,8��1��n_�h�vL2���2B�dþ���k"��E*��^��+���3�&�x��� �r�^ٗ�sp,)Y6;~0����Ն��HhF�랄�MA?Q��[�Q�`�5�@�NO�b�=��Θ̬����`)�8�в|Q���C�M�����wL+i"z�X�:�=!r>/���if?�3f�P��w����y���ߘl+��>�*{���y��<�u����)�.��K{��������6Ql�`�����h;Ή2�Oē��4ET�n�">7P0z�VlLx�&�U���Oh}��b���ۑ��ZbM4;((��qO3��S�O�7����N@Kiׅ� �Bu�I��J**�'�<L1슖���GYv���9kEP7���P�����ʄ�凘�M��x�D,�r�fݘ;X����bV՗�ׯ�����؛m�B��n!W�Xq�+b��3(��M_i#��%��+��t�z[�@�p��A�)�X�g^ &������<���F�F�x=Q�M��1�>�g�B�޹�~�e]��P-�C��48���[�K1�0�@4r�xi�uB�	6�1VA����"8l������ �u���,:u�
��ƭ�t��.*�?Y�ε�011D������m?
ql$cG/��0$�;�:��.\Z�a��C���h�b�[C�8&��d�Z��pָ��3�k�֭��
�*�z�1�J7kWSXU� �H�|t�����	���t��V���=���OxEv� ��1lE��}x
�n�:��N1��1���+^��Է�qp��Dp�i� S��Y5=h�r2��Cp��	��⠄<��+�}Ү��f��vx*8�v87�&��Z��@��4�^퍬BL�WI�g�-�Ϝ���U���BU˕���8�(	=��7q�á�)�Fv�{�h9�@݂�(���1���7�9/-/�K��x�v�j��U��P��8�5VLoT~M
�i���M���{!4u�T�v�;:��u�;����e��޲q�(�^�p�6+���ts帞�,K�zx5Ks�IO��I��a��u/��G`�л"�F���u$zF��\��ϣ'��D"wN�.��(�|��o�VB����Sf���?y)	h�V���נ̓]�W�_['�8lCXt6��69\|އA5R�P[$L�@�Z?��)����F�z��omYs�X��5�I���o�w��` &P*�!�w{^1�1��m�g��N}�p�K����KJ2���&�/�(0u��@��`�K��!V��g���$�W8�P,Ƕ��?f< �c�2�����'d�帆�Q"el�P�V�-����=̯�����=�z;zov�;�D#�9�y�NV
�R� �Z�<��}��<�gʰ����Ŝ�WS�;]��%aJn��B�|_�k�2X�Wv�����1�lI�����Kxha�G^���F��Mː3�f'�7Y��Gy^t
(����>�"Gz�	�����༅ ��n��_�s�8C�|7tU��H$��<쇁oZ�+^u��:��=Y���g�=/)��=�����&��yԌTF�����Y�FpaV��Y�"��d�%l4����[ɡ 5��>'Ҩ��ǈ+��f}����K����i�h��dme���"�����!m7?�̳:��0Ӛل{n��G���� ����.Y2���Aؿ��%��rh9�������q*A7��E�2�S�>7��8�*2��lю��FM͓�}���
�eNf���(ә�n�0LL�cNG�5��v]5Ǖ��C3���lt���s��}��1����s=�S�7F�r�~Y=V���{mu|/�H8F���H=���DG��b �aE�eK����C1���Q�jcL�!NY��\�/��bPs���}��v��)Z3\��7��g����]��D�l�G[W��2�}�]�7S��E��U��}ʰ���b�>L�=m�������9!�&����ˊG)��J挘q�
pie0'��"a�"dJe�*�q�Jr���~�̶����	jR�ǱK����,����H5����M������=VP���*U�σ>�s�N=�1�v������W �ڗ�h�q�ڿ�*��)��1�y�����S&����C��_��^=Pv-����}ڝ|��S6{�Q�> ��g+���M��Z��{�`}Y�]M!�'1wHC�m��}c�)�<SX���-��.[}n�_�	ܤ���һ�U!�}���+�̿�}��~��^<w�U�x��k�O^���͈k�7^�+ti"l�T��b ��X�;�I�c�����j��^m��y_M�"���M7�|��Ѻ�7�ɋ��*=���:! [���ݽ���Y��'G����`���4Q�;쟼j<Pyd�e�ȑxΆUD��Qs	��qԵ��A�R�L�)�n����6�3��<h�je�<:V¬�h�G\�}����^�7a\�h ��:$|ٍ��6.�
L�.�A[9"��>��C�G�N�V�`G����Pȍ$VO@MNւ+\���O�wJ�PNn�	�O��[�%��H��>d��c�!36�?-��|���ߖ�l��%����b#1#�/_�<A$UX��:�>�o�}1�,c|��͒>�C������(0	 ��k���D���^�}�s����%./���@�S��A|����F�H���a0a-c����݉�"IvI���t�xTn�j`5hpi�Ƹ�o{�}B�)�w����]~p�uT�M}�!qh!�JT7>�g�P�v}��9��^��z/Ej��U�-�نA\�T�S^�We��l�Mky"j���q{�Cٙ2�W�����P*�%�uʽ��,j�;�#��=�ӞO�1�5����F﷩j���*�Ȍ<���O��gXK��2�v_@#���o�O���W��^�+5� רd���l�r�n�pG�]S����W"�I��K�)�"�j�{,U;�f�;��a�RWSz�n@K"Z��`���1.`ʏN��B��h�ѿ�eN�ƈ��MT�2ԯ�^�>+�g ����p���O��ӬiJ��s�
�|�J���S>���O�OQ�_���́!i��2J���eq���F]g�5�'�Px#1�9�uD�����,�R��M����։��!��,�i����pT���{�˕���L���W� @P�ce�+���t�vgh�pLꍟB+�)�ICX�7�4wˍ��1;QN��'�i����cCP��}�r�q5&����V�`W��l�6z���P?�Ԇ+�N����Zt�����`�gfgZ��}{�W��m��D8N���r�R9�y��㮥E:k5��� L[2�T��aW������b����H�;ya����k��3��7Wc*)O�j�!p�hC��&�>L|-F�[ׁ�z
X[?�	��W$�v9�3K���x���!�G8����
vC��|��:n�]�F��6:�P�� z̈́��1��j:��TwKØ�ԪA��jO�j�'b��^���n�h�F!)�1�c
��Z�[N�d��ÖH�ힷ�R�����PL|�f���y�[	r�u��2�|�s��/���EN��x��G)-��T�x ��N��|��{<����gD_
���!н�KeH�Q�� i�����@�.�=�Ouz@��5�_�����7>�IB�2�.D Ҿ�bWM��Dﮙ���R�"	|�Z������BMH��b�mJ�L�ف����o(�n�-Q&���ƀ
0��[a�+=Ѻ�IM��`��c8���/Y']ؚ�N\G��Ҡ��y��.�x6�4�J�U�X��h��e����#7J=
��=��f�>0��(����X��9��ڛ�f0z���|���/�+ɌM�~�F>bPO��x�.t���zzP-]҃<߿�%B\�������8,塨�'qz�a�k���D
}5%�%c`�8�
^��Gs<��U�_��Š'��&g&o+ bb�����;�b���đ���$zA�+��PĢ��x�0�g�����L@ʈc���^��c���.����$W+Id�yGH��J�w�����ŀA�W������������9+5]���h��������垡����J����ȸc[v�S�1�����Ǟk�)5cp`F��^q��Z瀐}��c^Wޖ5ҹ!$�v�]����c��K6w�:{�����w�J��(��`�GA�D�$��m>�d\���A"$���K*�0+�2�M�O�G@�oݱN�`Fg ��A��)v�wc��X#����
doS����4�`p6m����S��>r6XL�b`z�6���#�Lr9xĿ6C���Ǎ�׈�_3ǿ�p��@@�0�d�%1���y^�"�
�1Q-s�i���l�> � ��_��t��UW:�\u~�nX���L���q���N���LMt_��h��u'�-38bx� ��hŤ�^��~�
e����&��� T��'��ߋ�5����hU�9�a�F���:z�)JҼ�l��ji��������cq[��^#CH����]�o��Kj{B�/,b�.�Tm�J*�I�UB0�_���̟b~V]��w|�+]oϓ9�k{���ACwq��}a�*?$�WB�^:�"���wy}#�H1��U�2���~U�܍������뭜s!�J� J�A#^�l��l�3�x{K�k����N�~Xnǟ�eH�D����6�5�F���3�ߥ^a���M�����֏��.WrԆߜ�Ə����=y�Q���G���ȃ�א��KT�������l^���9��it}��'�gj7Rb�@|(�GE�4�Y��oI��0�$�2���ݛr��t��O]��=�8���C1D@�wHȢ��Md�����.*��H�iCr"\�^��F8-���y0�9�P�{��Ce���/]�8��su��S)��G�����Ç!ɍ�"y��dh&&ݯ�Z���U�!�!V�^����X�G������.�4����u_LQ�qΊ��#3:.��sv �?1(����/��ϝ��?5#6��(q�ݘ����Ub�\l�N)푺��T/��̡�ZyMM��Cr�P�w3]�a�E�]|3s�L�h��§��k��5`�7��E'��
;��2<)�qP��� �/t��Mu��*�g�$�`����ٯ-~. \�w��@�����s�@�͛`n�IA�\�II��t��T�����U�V�ț�A~I�Q5$4���ӍhS�ݠ�Ί�*'�bp�в���8RNs�ecy�����ĉ�Ěw���4�1H�q�>d��VmrC�d����D_��~���zl�+D^�w��� ���a�6/��-��/�ɘFK┽�#�i\���(V�W+�ߕw�h��±�(�Y�\�j��_�إ�.v޺�eʽȐT��z�1�r;�k,��Y᝸>c���J�E��«�8��E��!p��!�	I��+�"�����Kv��ɶl9Vo�z���k�)E�H�3�=t�nn�����ƾ�B�_�뫗�����	�����KI^u�
��ص��V���z{l�C�DV-�&P��쌪��k�	o�M���dbc�H����i�1M�n�.��a��٣� ƭ��<�8�b$*��{�A�BH�4���B�o��I�YE���2�W��K�~��(�y|L�� ��1F�-��\[E�F��%��+,���#������!���-2�U0:��&�hio�gO�)�ޞv�z"���̤�vx�8�i�N!=��57�<ѕ*m*�]8�/����OG�P�����Q+Ș�i= �9��k�TWo�0�����:}u�b����e6E��cSi��! M��慸����ĩ#|���Þ��Y��Ds���aW����<��tJ�ܹ�i@ޯ�;:�U��GGϫPM��e��s���<E����+]��E�V���2��Ѿ�l�/I�_-	�x�_|c��K�x+5�A}�_غ��������MQ
�sEָ�`��2Z�-V�?��G��Rd�. F�Q�0�tF����Q�����>��;܉���7VT��6�	��:�P�P��������i`t6�w���xԛ���}+n+�H/K�{���[�z-Pf,�NsЋM�$���3s����Y!? �YH��[f��7U���&&Tf�<��i�9���[���B���s��W�M�Mܰ���,[��_F�A�EI���+�u4����\�\`�v5@\�2x-I�˂őV!gc@��W/%6��˹22�9-��t�px�B�.�0ׅ�cF������p�v���l�l��q��0�;)�?���Lػ�L^'�{�1�T4��\i����Z��ә�y�e*������x�?&�|g:�k)
�=)+���D
ߌi���iqj��Y�h�"��<-��A��ګ��S��ojZ� l
-O�	N����5��+'�k]hcc���XUZ۞{"�.t��*j�Ou���l����(W:;�5�c�{Sz���0-�+е�z��r���f�o���>g��;Bo�w9�ܳ��zH��f|̓���-�1Ak>���=4�b�����&�FPitnvV���b�R�<���s���p���sY
�N��?��Y(�̺������|!�~^��ݿ�=Ʋ��<���=)-�|�W��X�3+��U�`�J�3ɖs��ʣ��jw~�L|;��1v����ӑ:� I����pU�A�}��"z^��6���x<C���`+��'.x2��Z�&Kn9����`�?�%�yz��a�MB9JГ�'����{&�����ec�X�rӽe�7�n�3+��)��B����wޒ�ﭻ�=w}����1�"�Մ�L��
S;���e���)J��q*l�@T�%r�Y
f��#�X��HqV>ۇ����c$��5 V��vjvq�0˗F燙l��F���c��*�A�7mHMJ��z�έN��%�:_U��2�R�|b^@����(1�<��qMt�I]_{�9�h`��oI=���0|Sx��z{a�O��Pۘh�ִ�+��0�*o���S���TL��R��6�y�:&�ij�Q�@�yD
��{���'8 �8v�����ܦ��~O�I����EߊI��� U:so�!B��.?���,_��\!8�bjS�]̦��ƤC�)�NI[�oi��<^ ���xe?���s��)X�$��a
2W ��Ըæ�}}�ߎ-P��[	�
=�<�wz�����e�6]V�A���$��X��zD�_�܉I�
��7�SJ�m+QL�� �̧�����)���f��F](�����X����YY0�3Ay�2���B�Ga��M���Y�/l�Y�%(�6��d_*C?�=�	09q�+��+W	2�g@n�4�`0��fTg?컳��N)}�RU�NU��U����:��2|A����X_�F�ZcGb&
Y�7o����x�D9��{���!V���M)˶��j{�� �\�%�I8	c7�2+��NnM$t�����c1�2Pm��
g�T/��2D�TSipę$X-�p}�1=�6�E��S�#|�ݨ��F#���L�й�x��$��Ч"'R�k�����0d�2�-�=�81N��&�x5$hg��M�k��3$�f$q�g����4M&$~���`P����Dג�G�⥨�DY��g'��EsZ���J���CR�Ď��tY��O��Ӌ��ӄ��4�����5���
1=ӞQ���Ԇ��Z�vp���&���{�ldpT�H� b>L	��v B�y7t��� ��F��I- �����^U�]ħÙ��8P:\W�t`
����UGS�,�r�!$��]@J�-V80�6u�tN�υ���Dh�������d��>���)���/^�!��K�@�O;8{"���
��NԸ�w��Zk�x�L���#~䌥�t��Gr�x��&�̦;K=�Z/� w��'��Y���>X��;\/�J�=V�eB�BfҜu�өJ��5�b�-�w<���as�P����Z���K(�Q���M�w�Q ?��/����?�r7���8��X�N�9����P� ����y�Xt~�>�G�KVԌ��T�6������^CH��+��H,��T���c��KV>���A��6C�2417��42�] ˢ{��&���м�Hx0�G�<qc¶�K.t��|n_������!y�NI���^�^l0�]�<i�����14Y�s�z5I�g�NY��G�0ρ����N�5F�fFFd�}���eߡG��!�+�J:���	 �B�P�"� ~�����ڨ@8 �����ޕ�тG�<�_y�1����8@Tx�rܸ;�:^c_�w�Q���yg�vrH��M��`�������V9s���_���|9�)�iT�yx��j�i�m{3K+/w6�X�|����?�@��?$Đ3�S�ƒ��	�T�A @��y�Y�k����OA���˴�zA9�+01%E��/Y
�|]�(�z�ۄ�B�R��ɕ��U�M��O�R�jd]^ݏϘE���JG̀� 2,>�EH�X�c��*Z'�Y#5�[*o��B�!Q�.�i���?#���}� 5�E�p�U�,3�+�uu�[1�)R�+��������[�Q���Yo�����\��5�?�!� �Uں�֘�rA���zC�r�;<�5g��5$���-:�9�?��*0�x rN~/�`77�nT0v�?�S��aK�*|6��(Cp� \�c0�Hh$cf�j*�q�tÃ�CsnT���$]N_Q�iA�,/�������~�[�}O'-UO�r�����}����E��n�'t]Q  �AmQNr�^�q�~�ʓ�*a���|g��+���ݘ��[���}$�"r���|
 �p����)bz!CI1f�ly�������C�9�����ްfOM�MRx��u(�@����nR��X�k݈w���:[�9��{���Bp�GQV9͎�L����e�b4,�h�1&(�5� �\�ס��qۡn��eq?p�
�}-���_=e�A�òZ:�����'�eA��~]T�Sޗ��~��H��^��/��Ӂdh��@����� ��	~m�A�_1�Ｕ�s�cd�ڰ�7�>Ȫ��^��&sǒv h��D�-gm��=,%���`�mQD��I�P�.��I�l*9�7s��x��3�%͠y���z=�G���R�UU�"���[��ׅ?$�1��}F�۶�g�N4�1t������s����~�Z�VYp#��Vj�מ�"�WvI�p-�d��&��ku�S[Q�G����x��ʖ7řN�e9�u_�|�82��朣��m�ָ{b�?�B��o�F�h��ջ
kR�y�u+�P��o�?i���ί;@� ��|t��Q��'���J)�[�?������KY��l���^)5�wQ"a�jR�lb�
��݄���ɒ�ܶ�jR	�,���� #�t%.�[rKmgEű��LӞƚh����>>�Iq%��b?ߋٚ��CU�X�'գƆ b�����[�YG�G�N�p碿�wzҭ0���K��K��pr9����5��,q��H:Zr�a [�q�"���E!4�u�k,�m�I�!��Xf_8��VG{�!v�_�N5x��i�ō��l�щ�3�H�<4�V�"`"�����:/�9\��6�?����T5rae�?/�6S�ձ-�@���j2ZX��R>�	�_���uh�����?�,��O�����}��v�����b�t�m�W;Wܳ���w�
on��k"�����TBcn���M�k��ʃ�A/jQ�껄���d^x��A1�쮾�1X��k�U��fF8�D�̨<��ِ���kM�yH��K���'�ݞ��~�M�ۣ�ՙ����j�g����;�A�k�E�7O}>������0s�Q����+M0	b7L����V���-�I��V���0�g		� x�sw0�"g��}�W��� �K.��ӭ�A��o'-�6���r٣�GZ���M*��[��n�~��^�O���Q��ں�_��|u-�x�d��bP֕���_'����ʮA��9cT�=mb�no��Xk�Ѿ�;�ϓ����{���j���!�v�D��l��M��k^��i2K��6���X2�s�����.P��	!�!4�Չ�Ls��V���T�9�u�[�=���7�m_�h��b���:���C�D��A�!�tp��k��!{������)��X��-��"��z F8҃��\�jD�9灇nupu��?�ee��XXh�(�
2�p��o�V$M�"@��;2k��J
��*jVt�'�N}v��q��ѽ}�ZЈ22�L���x�5-m~L��#%��hQ���S��ԫ&��^2���M#�K����.�o?Z�����Փ�Ҽ$�q3Y.N�>n��lV4�W��F���]��I�xL�Lƞ���;��{�X=��ծ���:e��ۻ���P����,�U&
l�U�ۈ'O�s��/<ZIF���}wI��=h���i���a�5���'�&��5y�
�۔/}��_���0��A�z��Z(x\���4�����$Vk���������9"(�x����]��p�#!\���C�h��2����C���8X����ֵ"n�uT	���5�W���&ݗ3�_��@����2�b|:��� e�6�5؂�����1mWo�TD��L!p���v�p�1O�?9��a�4Tk͎7xͲ�HA�E+�qb�6�@3	ZaE��k�n��n,�i�yx0�	nRh��;��хɰ]z`>�2#�y�0<�@�G*�A�x��'�Z���C��!�O���ۦb��k��o*�������t�Z�	�G��挌7V��D��uO�&'�8j{H��%xv����`�;��D3�} ��<��M�bn#s�.����6��`�߳��ʪ��fЇ�>��H�Σ�k�RM9hO*�-뤲DÐd��V�O1���F<3Bn;V�,'�e�9!^ۧ�>�%El}������h�-#�+#C��sroi|�,E<���
�{C���0KT�zY�B��^�Ti��&�y�V��-l.�0R���5R��Esj�=���]�C?�~���X�`Xj�N���ޑv$��9���Eh�/۩�0#u���o��י:�R��N؋�&�W����G���ڽ��0C)��G5�f���"p]�f��'G$�y��/C���M�+�L������ÊÏ�sp�܍v���Y{t�� �ی�w�g�)���G����k�ň�O�.Y6�k�f!�%֎��0�B�z�|�O]��ѫ��|[�q��SNQ�@�):`�R`�2�����ݟgⓢׁ���y���"�����l�t�Sj�o��}����(��T��[qg~�=��!��yݨ��%���&�_��������y$y��Т�Hs�E҆%0���B���|4�g�2�+f�wz�#���#���VI�N΋S�B�\���sx���6A42��Ѩ����#�Mu����_2nV���ɗ5۫;��W��*�\Rn�_�М.u�1	�"e��E�cb9=��~� 9������s�h��)d���*�"c��ۖ��&�)qs�s\��]N���	
E�)f���]!����݇q�/��Nx����]��z��8ߑ+P��A�u'��-��Ҥ�ظeQ`q�����\����;?��R�{J��k���^�&��(��PB�s�� Z���ج�8�]zn�-�v~+�aʑU�&jc��d�a�fi�_U��B$��$ѵ�=�{�i���/��QW1&�	��>��갾JD�/h�xo3��J�fd�-F�y���8�o:���rF����&zQ���P��Ĩ<�Nw��w��G6{�v�/�0@�J�����l�"�ɝ��6@��;��z=��q�~�A[w�ԏ��Hn�]����q���}��`7~�z`l�߄vu�!���pkg��TN����:w���#��1�f��2<��zv^O[t��?���u�U�z��n=B"�Q�¤�/Kз���1�:Te�L
��1C��!q۵���۲���Q�y?C���;���1���1u.1,�{�5ѶIOϲ:����QJ�t/%`x��?�]���M�1w����)�Jh%�"ǆafrM��]d�/t��Q�^�
�m��&P�#o{���`�)�U�_c8W���gŉ&�7�����H���B	q�:1���$r��Պs�Φ�Xo��M��~�g�m�S�b<,t�"�4�:���~$k�=�<~,}���� �c�k=�h"��v��p�A�@VC>/�c����"�i24/��)��5��H�5�QX�j��k>��f�X�ƎR����Ni���\�bN�a�E�"�/]�a޺?`șBv��YO�M[EH�ʜ��b`-�Ǯ����]6�/�<�?�4{�q:M�ܚe-5�j��� נT`0{v �c��c��`����Z���G�3i����x�.i��-E4�5D����J���8����J^��Lw�k/�	�D�v��K.���)�Ɍ�hFd��h�4ٿ��Z��m*��#=��C��]3Ӥ�!0�+Hm}���#D[�D��D�S��|�X��G6ѢԚ�n�ku�oL��5�����d�\���ȡ^��gt���x�M����L�@֧g����\��;.��ߗ5	[�ص@�P�-�(RlW7D���H#�:�)�q��po�L,�9p��N��'�<>z(K�Zÿ���ns�����c̺0o4����$��s�u�%�Jb.�DQ����)�KG��A�/S�{�9z�r�sd��-v�q��CH	+���<e���֒��C.��'qa�Qxt��(b�<�W�֖���GԵ�L�ge�O!`��D����J�}�Fz�����Ex�qm�S�Σl���)J�DYJp�1�������\
�=�HrI�e&�*�ˁ���`�{k��Y�*������P��b��O��;��"�~�ME�9?I#)��8 }c�i�Ä����� �����gR�R���Ye�T��͠n�	��q��˼����O���bX�KU�7��SW�$���e��͉���\�'�0��l��ս��(L�zxj�#�H|-�-�P0� ���~�����B#�����ò.J����Q�xB/�A|��_u���N��
��&_�p��;�{-�Җ+?�'a��"�y�*�k��`k��˅�����#�:Ȃ���A<Z���t�Ga��fe]�����u:C�bl.p����4Iћ�c�
#��9H?N��	 �K��޷��n2|zǜ�I������y�h���ɇ�����o�>���H��~i��.��CC'X���h��2�K+���$ Y����w�6?1c�N٩LM��:�'+m�NB��`A�nQS��T���v�O�OZU෭�O��ڼ*��$%�~�7�z��4lȪ�	{�o�>�Ⱥi���@�/�u���v2�tX��-���s̐�:��WAD�_��O�,�w�$�����ߋ�8�0z��⬼n|�G�dop-�G��e�<������˵1��Z�=�� �w�7/������W	���g��M���N�l�8�K(����/'�ɖa3o3=n�� -�����#k�/�pX��8��$��|�4�C�#������9W��������Gh�Y�5��D��ˌ5PX��Ԡ��H�e%"m���Xax�̣w�-��V�_+�E�^�e�P9V��G~�;���6�\d��X�F(;�$H��v�h�@Z&Vi��9.B�Vw�,���8�au>����òa1��6�y�ΐyE�@	ū�L���	4e+�<�w��zb�0�E� ��:y�d����Q�;�|�'�i�I��僴~�C"�W�*�����r7}rϾy�����������GV�����v֋d��輇�U���n����c鏑��W[a�$$�XNstd̰�&�"�~�pf���#C����v5owk�N���Ћ�
���⧺����Aw���Z㧒-^1߀�!�^��RU�0�X���QɴY��p�������#&/ưe�hr�nv�I��*Z�e=.���ɝ"Gko�>n�"��ߚ-��{t�������ʙ�((�t��.�a��V&WV~	�Sv�V��d�B)�X��OɈ>Otq�*}f���b^��pwn5��u�HhX+��U���=�C(�+m�]��E�:�l�:��"�L��B��
�^�cg�3��M��q+�����B�0�12�����j#H�{mW�Nso4�_4�v*�צ����<rtߙq�i���T���M�8��qG���!M�8'+{�g�Y����a��8�ϊgg�Q�Ƚ�N��6ks>����]�����ق��1�y�W�
��SL����-6߿�44�XG��4�PaZ8e&����:�GL���`x��+@4t�>�=W�wb�;Q<:����P�����w�ǵۼ��܌�D�+� �pa��`(wɢ[�k
KjU_s��x҆�ȅ͚���f�F�z3�9��=,7���rY�ѧ���3.[�t��}���#����šn58�әFX��ڍ���oM����	�d�h��QJ�v�6�T`�H��� �tA�;���j�%�
ۚ�Uꐝ� Njw�����O�O]V��^W~f��*Ú�co{I���� �����|�/i�~�R�Uo�`�j�Ry��D.L����~!ޟ���UV%{� ��6��'�Ͱ����L=�1��O6*V۟��]��M��V�����dg\z>F����k�X�:IlK�ˤ���M_�&�� �݁[� �Q慄��Ӱ!(�"<�J�g���Ŷ���g�v`��[]�=��T��)�{�,���A5Ҭ��e�^
2�y���S���F4�YW�&E�����p{� ���^ٿni��_d��;otzg����Qeo-��8��w�'�r�4!������
���͛g�.s"����Ҏ�V�	�Y�ͯ����934��=�ff�!���?�f��!�&��53�W�5�O����6���BۛE�E��am���>��h�2�f1���=a�1P�'���V�3θMr=����f`�����<�A��XG��\Y��?k�n�L�J�XU�ca��`�F��-��0<ZmH�@�؋�6/�~gvX���s%�n��;��%ҨP2�1|u�4�F0���im-��hl�IU����#Ȏ�O<kH�ޫ���/�`E��ۯD"��ē;��V������t��v�J�|{p��/sʹjL��ݩgd3�T�97�<:}����bo #鷥�l�0O$�8̂����kf�x�����׿�p�2���V�����)��s�8�J�,m�	XާuHq��~tNl������5]�gcS[s����uÃf�l%�a���}5�L���7�K�özn��qx�ڝ���9�0�pv�)���$�'��2�]�F}��V�@�Rʇ^�zӸ�GZ���Ib�.twD~� ��m���&����T
oL�~�[e_uKüH$�R�"s�-C���0���ue%��p��giF��u�1�/_H�5c�-��4�M�#����� ���8��olˊV���RB-�;�L�2Uώ=_�s����<DGf��D)盕pL���Hm����}	Ջ$aY������ժ o��߯Ob2�c�>1���;Z��a����V���ߚ��N�g�*�;ea�x�k�ª�G�{0ݺm�Q0G�&|��R�7-����1�'�� ��e��Ů��"F�㏨�.�C<��)a�"h�}hG���#A��Jα4ċ�O�,bu�8�(YqH�7>X��ڸq�r��Ľ�7�r � {d�O�\�8����S�L�@:I��3:��M�W�1�p�.:�
xox�@���'J�G��Y� Ԥ��$N��q���Ktx�F��eԘ��*Ȥ~��w�j�r+�{��\Y�xh����4��j^o�9*�f�.ۄ������X��s��;���)O�m�}��>f�Q�H^ �	��S����Z�� e�G8j3^u�B$���h�w�"/Y�>�<wW�m�Vb�ц���<L1��@<�����-.o��.����������W7fgP?f֒.Վ����#���Qe?;#�)@�[d�^&�P���b�aE{�flT����{:����)�
B��u�W�����k������	5JW��B��v�Dgt����o�WI�u�T�>�����6Պt�id���&"�.�|#�?X}�y�)�oY_�����@7[?։}�NS-���1�Hk������)��W9�e��j�7��m��+�v�+������8lx�[�?Φ4^�n��5�N�Kz�ũ�wM�k$��QTJz��*�\����K[�h+����3��� M�Q̨�@ ��ڜqE�*��N>Lhh��	�1!��ӂ�қ��-�wg�N�`�I��`�x��gK���m�l�%�/ǗP��O}�T���2�w�,@H��67�p����RN*�\����B&�)���?�-�� ����J��/�]�흤��Q�.\"��y�ͺ�XG��tp!�=��+[-����m�go��PN�^�Z��DW���^|_�F�mr.O��V:��_��������� �6Xk4�|6Y�L��*r�֞����L��3/��l��4���h�1~ե�5�!�d�_ܒr4��ł`�.�� �Lk���^���!�m��Ӄ�2q��3�d�/*� q"UH����!]Sk�B���^D��qO#�'�<@](�mO}D\�P�~,�&y�fݼ@[���³	rBl�)ZHȐ��L���rꍂ˭A�'��K��`8>ZʪW����ѓ)e��ׄ ����æ�\�J�S7g���y�U&.��	�.MV��@���]�`V�͸�]�1um�LS�8��H�xkh�7u(��3U?Ó[���l��Y-I��x��r�Ci3��_����4[�K��Y�A�+a��w�|K� ��vZ��!y)р9^��
�Y��ym�J!\�˥d(�S�f!������F]��j��p����7@������9ܫa�1qj!��jc���qɏ����k:NɅ^�������h䮇L�����1�!/�+��O��`�i���/��^����۰�G
���'��nPV���pf�M�n!�8��CN��/B�@�dl�\��.1A�Sp�W�(��p`u2�ݠ�"�=Q�!VJ����xlEh�����#`���_�R��3KTP��{j��)0	n_��P2�޾�[�C�-�Щs��P�6�������7�2e5��pZ[��bD�Q�ob�J�.�P �
�
}]�n
�<�d�	VjZ��~*d�y����q�2��Y���^w��1,1ch��B���k��PmU��u.ċ�M[WϠ�S�� =���)^��µ�QB���i���[I6ҹ}�8��v]l��ҚZ5�E��h�C�}*"h��{+����v�j�\��7z��b��n�Yk�����b�A�JC���1i��6�-ă&Y�(�U�����E��Y�#�)/�__�>��$E�U��qխYHk��R��xKUV衿�K\���d�_��G�@*@1�-E�(a%+{�H�\!�]���4L 1.q:��Q�KvK`�$֜+��+,�,=���׃�ۻ0i�g
���h�\��{&|��u4uل�**j;>LEݮJ���ܫ k�g��eZ�~�ʏ^�8/s&�e��Mm���Z����������j���/HI��ޤ�A� �����q��W��S���(�.�r��AZ�RjR
E���Tj��edd�"��(��a\�X���u����n�Ѹ9��c�`�L�]��,�F���O~�A���o�^k}�"�CB~�hM��8��0k��;׎�9?!�fw��X��n��m������M0�W�ᨐ$�?slW��7)�頽5�sal��X�fRW��Kl�.�C|ʈa�cG�^(`ƂF�����}#L�#)rԍ�����Pa*] �������vV���Lc~�/+t4m���4Ѝ�������]��֚�U�lK0��G6C�4=W�^N��m��Cэ�Q��{F3���P*	)� -�x�����O��ɫ4B��K�Fs��ݙ�fw{�5��*��S4;�?ڨU¢�=LZ����+���u�^����G����u�,�(#2 ��b�4�ե�s��@���R�����O"�K{���i	�q�K?���un@���Kv�U���/yx[�'���&�ӭ�  ��a;�_!I>f������e�1Lℶ��M�lz�K�����Ƹ�G�֧�W�� ����(��˽�Y�L �{��MZ¢mR9ɳ���*1� ���n�1��z-,�gæ���Kd9Li}�����x�	��0���Z,r�׎BTS�(�7nj-^�V�=��SN-[=�r²lN���#��Lu1��.w���L^�wt��X�c�Q�)�j�x�[�����[�"��N�u1 & :��h����(~w�W�9��4(+��M��|����j�k���97�K%��iJ�t�Y4��|��Z4�i����Q���ϱdI#�|b�S܁Q����F��z}�>��-�X��׊o(��%��}t���¾s���hnFS\(]s�_hU޲�e�֬�q��d�X/W�|��d �=�3._f�UO�.��Uw(��g�|"��)�h�O�Mm���i�v?�U.�C0 }�l��/��_�k��KQ�Nj^�˥�CHG̰�+KȀ���5̟����zN�+ЙA\,��淋����٠������g����`�H�����X�q�@u�t�pa��H�9k��������U]�ʷ84w��{�Ü�/4K6�� h&bN�\#�w�$t6;ڍe�F>�zb�.�UD"�Z@yd���}�GN���%��9+2��	��XF ��w�W:ھ��\.��Y/����<Ɠ�V>��0�����4�cNZ� �;� �̔R\)�a�t |XSJ��?��bt#�ǔ41v��~o1% Qy�xiC)�L��l�*aL�B�d�j�D /�1%2�sz�-��kߜ@��]��A�p���CS�����[U5����J��	U�Q��f/��P�R��}h+(���j{�;{#����(hX0f��X]���4�x3u^��\˔��9�8��>ɼ�G�2�6����F3�%E�vXb=�ݕ�����k;WI0.b O��LtK��˦����b �b���n��P��F�޴����j@�)�N�W���Sv���q��rޢ�"��u,�♧��-;n�^J�B�S��d{+�f�!��m
ğѰ�g$�����8�_�;嚉-���NH��v����@6U���1�� �H�wd���LH>��5[�tQ�a�X˧����;�K6�̐m�l���@\���|�� :�I������q�b%U�
���T�?��9_FI_�Qb���k٬��M�@�Θ;p0��cQ@�0Fܸ.Ԡ��;Ԕ-�V@������&���An��D.̦�@�{zQ��jq�����e������i��x/�<O�k_��1@�n�5������#�����@�������+�œbr,�]Q�T +_v�x2`-Alc�_�7�Or��?���]~܎,K.G��u�`�Zb�-@T��5И���� �ip�|��¾91!Y�qђ��Q���5~�!�F�����:��^Yw��+v�=I�'{@a��SI3(�+��(���&ʨ���ܣ�,g�y��r�h��O1��}w��#��Yz"+Wzm��+��5;X�7�U�ݎ35C��eL����Z��"�wh>�D�M�s=Ȗ0H�}Y�
��1�Tn�JJ恾 H��{WD�*��D�Ϧü)f6�g�ڜb1��tw���$`N�2�W�[8+���׊��h��lO�R�����s��}@NΚv�kwE�O[��l�6��V{d3.����D��[��ٹLC���g&���	����VS9��>�4���L�U{�͓��k��cg� ��GZ��c��";e�_��/��f���;DO�Y�������0ǅ�?)�8��E��&��yy�}%�d�7 �`�uV	����cLH���==h���U���>��P`�K'���x��铇�ǒ ���ԑl��ק܈:��#���ڸv��=q����~�����<��ȧ��̳�Tk��
�7R����i����� w��Ұ�%K>��J�c��%�ɡ��k\�["�� }p��	3�tiK2-À�Sc���4�+��J�!_���K�'���>��h��N�V^gV�,�����`�q�z�P�Z�#Jݞ���$=p=b��/e�d
�d9<�LJ��w�0�Y�����	X��Qh�㤊�c8��i�jBXx�)q0j	O�4�eP��;���o��Ĝ��4GW�s\ڨ����%�5�#���4@�q>��K�_1�G���ظ�=͇�[t�G��� �L�JO����I�yjٱd�m?�LXm���n��k1e�˽⎛co���j�d�n�-Dt����:MF=M�-K��l%�d�J�ݏ�|m�tN��䞞P��������ft�ϭ������X�� �g�̇�[�#�Yơ	�kw���,r*p�Y�9�y�)��T��5��D��������@3G��ׄ������%�yUx*(��9M�Q�U~{a�����R-��l�n}ӎL��<�u�|5��e��� �_��.�1�j������4f��һ�������6h��rR� V�IsaU[����Z���3KDЬ�R����so��K�A��տanz"�o����j4��5Q ����L��2��w�2i�SF5UU$�G.��zB ��t	]�(-�)���9Q+�Hc�i�����DƆsu0.x�����(6x�w��~8/�.�Si&�@z}p�~6�$��c�[8a��:�/c��D?w� K�#S%��jo"W*0���D��@�������<˗碃�9v<s�.�]�� ��/5�yǨ��$���q��<3	Oy������+0e&WQC�̵Nuj&j��埄e�o��G<�W3>�HwT��"	x��PӻD^|�� �hHZɦ~4����9�̎�ju�v�Ϟ�h�_`uB�C�a��)m�N#O#�}}�6��V"��<�䗡��O-�:~�m��>1�-:k̀�n�� 6�Õ�xC�-f�&�K�����g�Z��rY��/P~�~Dķ��<Z����%�R�	��%y,/�=�Ȍw��mv%�'o4�F�h����u�ͪ���N��trA����Eϭ�f�(��W�ޗ�eߍ�7�r��da/Ȥڱؚ��k���v��h�y�\kM���6�3,������<��[:�<)�T�����]���l�<Wb����F�79��y��d�64�M��-���Mh@�B��9;˽�g������^-�Y�ߎ� �m�)`W^�(qI�VdP��A��V��u>EL�막�5c���Z�ّ���2۪
S�A�]�|�^�������^]j�����ahc����0rql;M�>�s��qM��c��.�AݎǦ���)�JlKO�L}�k�}�q�~��0XQ��8֠������d����D�:�B_�ڃ��`c�X7nKϚz�Ҍ��������:UM�;�aM�oe�d
�oT��B�^����p�w���W��/-���^��{�Sw��Pe��"PZ�\Uk_����FM����k��;>d:��B�v�,��f�5r�g҃��a���CсlA^ׅ�=��eaS�lcp�v�c<y��(JU8*P�fGR���o��^�w�+y����+���L��O���SZ,����wi3:?+�m��	k��.2&�N;J*�?�j�K��F�p��� ���rgRm����H��H �& ��.�/&4b�D���S��	<L��l�J1�{) V�W�	�����G$(e� ��
0&�)a.D�Aa�t��F��kf����
Xrx��M�$)�Cp��>�����Q��_+�KbWԄ���2��S��Kxv��r~��}`�s�S�쟾~�Y\e[6���+��D�v$��8&�)��:�Pm9�l���m6���W����˪J�p��a��~U�K[ƌL��i�9Z�^3��i���]2���	^�ے�T����'w�A�~ `�Db�6�m�G��V�0��W�-��,!񩹧"tٵ.6���H���P�޸�eƯF;���1�y|6π�U�rQ�����;xKY|�����b=U��r0/&{���[^��"&<��l�&A��j���`!T�?47%]���r\Y�Pj��R�;g��Y\i�f��5t���hj)��v�Hb�����e6�]ڋ�(���{K!�WzΥ[i�Xmp⏮N7^K�147/O��ؙ���6�>�)��lMK<M�lXvTV��՞L�,����R���'��Y'�V:�N?V$z�l�E���?2zX��&r�\=��#G�{jM9��N����ձ^�CP�3���sh�]4�#�}}T��@�>.MI�F���O~�Ґo���T���1����0��@:m#Ϯy,�@�k�1��	�Xʵ��Ig�眨���q_��_����m�ѼL�>�GAM$a���#w�ǛBpb����a4Y
a�a°�Cj9�
�OF(Da�����`JX+��W���{��GXt]�%��f�,��>�%�X�(�Jt�"THmC�haLl���{�y�Խv31)�`X$b�h�����+�F�����c}���}�x�mo_����S/z���x���G�ۂ���>�b�K��:��٭�o ��u��KA�^���v*�a���T���7��ɱ�jY)c|hƣ����Ax%��hp��s��2��@���1Ah��OR�Џ�F2S/i��	���[�M<��Au*����$�u�*�O.b�&{x�����2���e��n�?�ۗHfC��E�����VW�= Y��`�惞��OO���wt�6��2E��EI-k3q��R> �C�N�����մi�?�"i¡��Y��{�W�a���On���V��u��@��j(�~�f����:��'��WI����"���>�|i��Lj�iR�V��%�����n����Tf�댸�:P�J���-wh�+�dv�i}h�fӪ�˩�/�5n��2" l��9�)�(�'Z��Vo�]������=!�վ|U/��u����wxC���f�� �M�aa �gaV���'�n�~��KQ=(�&ޗL�'��Q��]�b���7��9Q<ca�jqz$�@��¨��*��T�9�@�7�~J�˱�Sܧ��^�,��������;�]~��1h�ss� L��js���������$m�
:�أ�m�NC+ ��jb=	�i3���8[�q�
F���+�-���ip���?�����J�Dw�����UDv�2����O�s�sx��L����[��{���^��/=Y�Ghl�%vs�l�7�|��%��L!SLˁ�twы�K�H�]�CP�h��S7�3Xc$K���A�ˮb4�R������s�/�3yY��b:�	죂P��
*|Ƙ\����`�ܹ��Ť:f+>�ȱ�
�yu��gWb�'h��p�L������c\j�Ɨ<F��7"|Ŝ�Nn݌���s8��
� �f7���-�0U0&��7�t�k���n%-��	lL!GD0�i�j�{?Á����W�����׵IS\�Ʌ������"H�V&(����a��\Q<��fd���SD�E���6��nŲ֍8���A�؈�ncsx8����-p��r�A��[�R���c��l�ˤ%�X�W��	��N����'����
��^�}���+�(�7���X��G�O�)��:"�Ŀ�(A�m�`|Tu�t���۔��%ح�ZdֲF���M51�<"6yp�T���(谴XU^f�8�ǽ8���X��� av*økL�9�Lq�)�����^ύ��t+�q�B���TMQ�NX���3�P9�C�A�H�1g�VNDo�N\�)�߲ _{�+��^�X�PK�k�ٕA�
��UT��^Aȧ��Ժ~Җ��9��fMg�TH��i�1*�/�$����d� �����u����ʿ�=V��ۥ��Wn�����5��M�	����9$�b�͜l��0���� �δ`�3�$Y��v��;q�� �5qq��9@�F��|�;���}��a���&�|�4�c�(J�)��O����;� ��./��O�|{��o�&WX]�Y�@,��u�qM��=��'qr9͐���KlgAJ�Ƀ3-EOu+Ds$���)�������w(�kS�%����OI�0:���o��q���7ԭZ�Tǒ{����zSu��P`�9s�q�Y�3����$�t[9����$�O�^��6�p�D�'�T��c�ז�rѺ&�:c}ѩ���k{��JѸ�_�>鴓I
���US���}�����q�1C'{>�8N�Sf=�	�S^���O�,K�/��ɓ���Q��@�o��2�؄P�����E=�ާ��ϒ��:�A��c��+O�['۶�#:w
#����T�x\1|V=�o{�
X_6��l-х�(��{�x��k�=!������GƷQ~�kY�s�P�L�*��
'%�A���)���(Fh�m	)e���g�׼h�ȵ��Hc Vh�|i���yT'#Y<��S]�|-L{���#}oi�!,��Ap��k�ܞNާ��L�@wQ����v�/��1;"� D�u�(�x�K��Y��լ�U��'�zTQ�zM�Ĥ��0�J7����"^ۂ������r_�p����ϟ�Z^�NN��T�_���	 �X��K����[��<W^\3��P�  ��i�@%9 L�n ?�@���娪�`@V� ��l�8��霗/�j�j��+D��(�R��lɶ�?b��Z���i_�+���gE,�}RR	N!%dqKI�{?��7/��?�ro��j&�b�蜐�Y���Y!g.���D��M0d�6�>5�4�O@ʆ���3�T�1��ut��	�pB���)g�~�K�RN�˹}�=�o����%� �k�a�� A�:�����Ʊ�@!M�j���I�OS���P���+%2��;U����>@����n��r�yq��)��F^XX����فT�����szw����yZ��Q��|�﬷����)�^�!} f�"�J)ّn`֢��C8w~	|"5��db'�~^��-��a+���x
��{�U�!�"�s��p���ي(z<�u��C �W vl楴#����Q9�x�W����rS��d'~�ml��p,���l�:(�X�$I�E�Ͻ�U{P��W�W_^T/�A�܌Ot,�a����^P��Nv�ћl~����^f���0ut��n��HcV��L��q!a2x[����Zhf�6�)�y�:�����f'�/���a���F�L���a�� �,��������h�~���0�^�����_�]���ZF�	��l�uBQ܁�GR�qS�Vi���DiQ��`.����?��1�C}�<�ۼ��j�3�T�s���/4n)��i@��")H>�`���s<Bp�T��s�sda~+����orf����4�8VT�TL��iͲK�8eL��`�%rk��!�s�Tg|{�Q^S��v	�ާ�;���a�=�ʴO����ioI"}4�in\H�
����O����Ύ�m�e�E�e�5�x���%2���wHw{�i���DK�"}O���#�l7S�
Pd�}���%!�Q�z���Q�Em������_Ca��v])j��@����$	���Ĵ3&-uۃ.�V������z��'3j�W?��b;^�7���}�E�1�`����qu�G�Sda7�<�]����~H�M��@��[�����_���o���lŚ�Qp^8Ͼ�.�.�o{C�?/��NN��Ѩ��M)�wBT��9�:�Ðs�[�}���ɱc�6�����9�H��e��㑻�q�����!r�����kn�e���1����Z,��=���֛�Zk�ҁP�	�C�q��C�{})��a�4�&��Lބ87܁F@�\��Y*w�+�j�S��m�ʲ�W�<����[Y�Oe4�yB��{N5J�������!��A���j�i�)!tJj7e��gN���X,#��ǯˈw,� ��3�!F���\�B|�N㲫�����w���hBuU��07�����pekd��b�󐟤9���)b��}O�!\|�������e#q=��B��봀%!�p%nG�gqk����n+��bOZNi�N��-B)U�����'1;]��8髍�cav��&1cc1v���{�g���@�c30���AZ��$f ��T�6��ch�����y�ڤ�F�3��&��;�v�q�_�2k8f��v?�"�:A�x3�և�Դ_��
�B�M��b�jO��:�֚��
��U��r����)�:�:���G:-~��݀ �����Y ڀ���b�hؽ*zH���-I�ػ�����A�Ý����d�}�O�r<@�fE�'��>yR�[$����/|�k�C��ĥ=�!�;w�|�cC��=K��	�Ue����w�US�t�q��3��W�	�  ��H�>u�t:8��CR�n[��ٔއ���˓-ݏ2Q9]��F���Mv��s<�沒��|���KDM�(�B���8ݡ��^l��P�J��M�;>Ǭ ����R([�G˫�_Rz�X<���p&J�\��=�_�� Y�8��X����R����,Νv���2��_ ���[^�\���� � �	:)?�
�|������B��Os��;.G���&�8.|����fX΋�saMh.������E�,�Wr��Tm��d��DQ<2���@J��=d:4��PY̹h(
k����̸I�.�S�@��m��{���-�փL��XI��N���Z.�(E�	��%S�Lb�6�	�:�L���I_�1�w^Dm�?���@4�C��{ju)S��s}=��;?�}	2%8��!4�[�0�w~k��f	�v�[{;�����̏_�ڲ1R(-���5���B�-��!�50`�o^�(jp�����N�ZK�sDL��
x�]�g�y�G��k�C�@_	�Q
j�w�L@��e�W\\��+[c�E�,J�!%�39	�}���O8Cv�&��e�u����ѱ5���l�Z��}#��<�7;>�D)c]�E^�
Q��N?�V�z2�u'��� �m��$���mT�C���&:��cEp��1U$�"����d3�c4���D��KMʏ`�v��`�����gVbg=�W�8�r8���k�C$�G��O3�ҋh��V�i���X��g���ʉ����
n_U�p(�۔�$�p{���]Hw���Qʄ�-	6�"gUR[(�=ِ���)�F�š!����n��1���X�ĆN���f>�w�/ �ľ<׌'Y������� ,�
�����=6;���b�K�\�R���Z�Š7��G6���#w�Y$H�k������`VA�;��/�/;����)�95��G�����
!|N�.̫��C#Qk�ި��7P��ͦ+R��-��]{��G-4�Ҧ�YW
wocb!'��meAѡ)`�E���P&<ƅ��PPu��E��H7g��������A�d�Gʏ]�<3D�ؚsU�m� d�Y/����Ñ�x�ɋ�L��e����7��v7���?�$)^ҋH�Ӛ�,z�ޕHjr	��G�?�Ё�j��=�K}��>�h�b�X7������Wx���x���em���q�[V=���#��J��u�Fvi�p�[_9��e�\[�o��*]��C��)eڣ�|�=сq����KQ}|�瀙R�4/����ZId��R�M�f������2|�U��D��+bUys��̼ ��M�P~���I�,��O��dd>�
�f��M�v�[C��LB�ŷ�J����hPLP�M~F��������Ϙ�:�(|��T�_&�3���`�(?�D��b�	jrzL����W�@�?�T���2�2�݅Nl�� �	1HE�"�}�㑿��W�̜��/_�2�����H�����d5}P8�eRc���*٭��?x�\锹���4q�F){�_ZR?+�v��7��x��;:�ybd�� �4*�|���pM��U��f�� ��^U�s�k���4�3�lC~�5;�(�'���ߜ�]3�r���_ܥO����8i�p(f�;%y5`���>e��C+w�v��G����LQQ��� #ܯ ��s Ǽ������Q�cLft|�a�}�w����ǻG&�<R�{:��ck�Փx0��tAO������Q�`s�5ǟ$E�q�`��y'������zBcڡXw[���f��
H��P'&�x����n�.0"kk�),+��-|��D�aE	`Roh.�#�*ʆ.wU���0nRQȪ��<{�eHO{ ���Z��_?�s��"!��J�����V�7m�z�Ŀ��'C��Ɔ��J�ԯI1��O����5|f���u*����q��U�g#�ݗ\ʚ"�P��z�.����( ���h&1)9_���Y����OO���&�Vr%��e����U=��한&�� ���y��K��S�YS���Ȱ���] ��n���;Aݧ�.�ty��)�����)�=p��#�|U(�=�/��S�:1���w�E؋j�Ei����.�@5����U�(����W]��4)\I���������ӄZ5��0���6�k�kc=��{G[3����<�%!���Pn�H$�������n��/c �V-`��۪%6����yݙ�Ե6q%��Wn����X��w=e���i �k:��Y��E���d���E8Wcs�(I=x�$їS~NП�i�sl��h��I��|�����h؞�״|�~�#"��=L"s���Hw>�X(��J��jF�O+�����@�}d��lG�� �1>.�����Ti!o�I��� Ek>A�Lb�%S����s��\���@#Q��4��������Ct,�V�[�r/ҫ%&��_zg
/n��kK8rM�FW����9\�b{�����M���b�8�&�QӮ]$�i�g[��h����"���9����N7�m%H���"YGP�8�-M5U�ƀӞ=��0ȴbo9���+�r��	]#.S]���[�����IʹU��17�y��1�6����`�"`��
�8�ߊیPI�9>C8���-��ˠ6��U2[K&F���4�֙�n���Jzꞡ5�1	�i���C�Ȋ��z��c��Y�Hӣ���T!y
�I23ō�i�9c9ҽ k��2Y�p�Y��O�3y��j	E�^ �m���ñ������'z�7��O�7��f][��զR�?&����kם��gq�y�`;3���';�IC�NO"]Hf4�XѺ[u+�۩��#� �7uˆl�| �=.�ȋ��0{���tPE�)WX�s����_�#��V�v���8�-h��|��B�'�q_�����a�`�Yj$7��ۇ�hc�;<�H*O��o���]d�o9���ps-��/��+f{�O���F������3��(�����B
eW>�	����b	����z&�i����C�M�2�@�6�]�cbe��S R�Q�#�4��bGq�&3t�@�i�z���e�r^q|�ל]C�����<���?T�D5�FaPMIb�����b�0����L!��:?�(�fV�Z-�A�Y�K�x�YB��t��	�)�Y73���2`�=�^o��;�|bH���d:l�P��`)j����N0�\|qP
��4����`��d2�;��r����*���f��}�i)?��jɺ�"�3Hk?�#J��S��v.Ҹy��훳��H{�|�_���O�(�S�G`������d��������f��R`�8h��a??F�H��j�ys���Y���;�]����hm�_$�V'y7Y�����=̄�~x�]Չ�\���������#)�.	4ʩ���G
PEA��#�}��8P]h�pY��e!�;��XrC>�DU�HL�J!ظ�^|��x�eR���'7�[�<r�Sʢm�/�)����53��u�H�����~���D�]����z�1Yg��rļ{�͍�R]����O6H�q�����T���-G��U�K�:��U�J �/�����O��ʾ�'�0ѹA�I���s�֬�<6(c$Ne�mM�>����0n��7�ĝKI#����d�h�fX�~���,C$܉7����̾�У�M3�������='OKk�5�GDΓ��M l����x.uii�7���"X�����1�)�x�}���Y�#���H"]P��߯z�m�ELM����(TP	���{&�����	,�#����]������c�f��m�s�s+��m{�(�XN)�ǭ�:���0G�Dt�Q�q����T[�?�`�+쌶�q�5���7�Ͽ={>�葖�jw,r����G�����[�Cj�V���B����Ż���zf���,	aF9HPj���,)|d����$��)k�/�����ޤ^�'����v����/��D�W�G\v�C�L��mB� ��/�I8�H~�eZ"?�������p����"�:�u@S#عS��5+���Ɩ=�@	�I_R��ɤ��
<-E��u�9o2��B[�9U�0�ŅOYf�VDf�c�����o�#c>K��Vdޚ+<����5�K�|%>��ެ_`ྜ�=�R1�r��X�Ӑw�8k�:��A����S�B����*��)���Q�� P�]����N�����s�	��VU*�3��_��+p�ը��9qJ��n�%�#&�
`$g����	e��IIJ��C����-s&[U��8c�����1�I��ٟ;=~�����N_�����M�d�ӛ!臠�f3��yH?����;�gw�$�C�r��I�hD�@��V�*em���j�}~��Z$%��!�	C�
ӟ7�$k�՜R��z�Cqy̯%��y��Еr���y��rp5��e 0J�N�$O����0D�,U��b����U�U���e�ǚZ�<��W�A���u��4��/R\�TF�'iG�H-���ik��A.#�
\Jo6d�����`��j1	���LO+d�ΡQzvRnn4�;<��+�ɢ�4.�,X��D�50
�gԦ��bd�2s)���� %���@/�W2��KJ5�o��u:&X�ǋ�x����M4?��@sr��C�*\PD3�����;[o��i]wL^r�Gԫ#�t �
�Ը�-4H���S��<�S�����/K��Z P6@�9����C�� ����j�6,����.�f.�\����o� ����Ew�^F(�ͦs��ѽ`%�3Q��kݽ;l��o����ͺ��ay҇)�%���Q62{ʺPw�;Y)��d���<��7��X�G�]Ix[�?B�����*��爚En�=��ݘ��5�Ʀ=_����"�9�2���H2�T�*�J�Ѻp(�O��kᜃ��s:�U���X'���~�H�v
x�
?�$��~͊��6�A#���@�9�F2F �)�)�%6C��kG|5��-�}��~ ��t��	`R��z�{L��QgV&�%�7�p�}J����ߕ#[����6	�,��:�$�D+�j��l����x��xn�W�=�΅Q- �G�?�>o�ut��V��K��l?��@=
��"mɳ�|'�Q'���j3�����bizn��bS;ƥ$)���&�`��wj�SY������k����m��j��w(��M��n���-����Ds/e����Y�ɱ���(>k@aaa���`��n����rޥ�[�=�g2�J�A��L�-��Czl\]��A�2�� �H��u��ZRP1ř+��8}ؘ�i̞�¾0�9�o���Б���pMc���a��#�^,��>���t�8*�4�߉K$���M!j�JK�!�����Q�gCC �|@�����-���^Q��=¤�swh<7F��8l�x�N��b
���ce>�8�:�h�靵!I2<*�1���E�5�d@*�X]*	��1�l�u����)�08��$r�)�'�_��E��ÁY���Yd
��Y��n�v�����rf� o��߀c:.���KV��T�Q09b]q/<N-Q�yGy�<�?1�i�¢}��y,uY�)\����ڔ��'˾��p[��N��sF� �Y�{][�JWe��L�)� �8˝��x��a�=V$W/�BK�T��O'�ѕ�ۆ�ae����r��� A�q?clH���+Bg��彳�;��&T&�i_�D6�����ĶTg~�#*�+��ALZ)��������`b�Sm�j;�m����*m���	n+�n�4�  H�ÁH/F���ЗaN	P����M�fH���߇�Ec�7L��6�L^���A{�B��"<uo�ǃ�#�7�ނw?W��͝xͰ"�i�� w���2���^�0ǁ<g�T'�sլfGhzC��j�o����9� S��A�(����8̈�$�?�]���輑��ѣ�.LkR�c�~�r���+��rH5P
�4��d��X�3'��w�T��	àt�e��+B�]T
���#�Xٕ+�,
�%�ŏ>�A��p�w��a�2
J�Bרj(:Cik�~2Z�ԈL� h����7)�7����K��2WM��0�ڧ귉���"�n�cZ�eG-80����4�C�1s$$���80���f�X�IU�������YE�+��7c�1�,�
N*��)�Th�;�6�!v[��|�8��a]e�`!�d��WH��G���d����u��%.q���fWb��X��~��K�� �����!i�vz��XL���~��F ($f�rO�b��!���-@��?	��;�Ge�/5w�7���	�de�D�j�H�r~U?;F||�k��?��_JZ��Z��cP4)�V�	k��`���que ��&�œPHH��*�г n�^~�d:#�dE|C��㻁$f(���������F�3;LF�������36a�X�h���+�ݲ'����y�APZQ�64��8+�TP%����]�e?-Ǹ�
����5ю H5�#�3�/Z�o������|5�ܯvZ� <P�#��+|u��������1�� ���n��O��c�[�dw����,��0��BO�G}�?��_-�` 8���3U�aރ2j�3'��M���BK#)_¡�4(fD�Th�p�68�嬎m;zL��_���l��:]I��0�x&�C�������Sف%�
��(��E�v�\ػ���M8�x��5ԧ��8/�%v���bE.��y�t����P�Iu{H/�OC�ۓД#��J��HQE�S@-��kl�ɮi�Q_ؔW�h|��K� �j��eǤ��%*w�ܩ���������i& ��D��+�EI��� �^ǥئI$N�l�E���'`��#�1�tG�h��.i^���u�}b:F�5Ɲ�F����,�~m�d梌�÷r���'��~�#��])����J@����G�>k��b�i�١1�t8�{ I[Q}�����qX�X`�;V�&��tVP�f:��d�F�.hI/���BC�^�t�"�����
���6`�����[}Ha[g���W@ʾ�_m|K&�fח�����2�l=��h���m����vf�O��
��h&�^{�@d�m�=��UI!�k� ��Sgb�x�&q�dӲ,���M͓��>,�|����{^Ðg�l�Uޗ[A�=/�|]B��-<�~?8i�7@$g�$9�ƒ��19#�z���*�>Ol�j_��W|�<�k-R�Y.���_�}��c���x�%�Kǡ�=���BGy�"�*U����X�
:=�Κ�n�ϖZ��v���Fl��W;{��LlhK5r0VT��0ss��@"(�1�7�i��u�?��M����[�u;5�\�A��y��;�t��e�Ϊ��uG��:@6g����S��Ν�hA�}KB����Kby�Ć�1Fc��7��$��m:g���dI��L��
�ˊ�
>��nI/���_7�ܝw�L��ɾ��r�5KF��<}��[]B(��F������Is�쮿'�e��}�4U'��?]�+���Q|A�7ɻ�E#h8��d�5K�y3�� (G�ozC�
�.�>��1���A�b*B`g�����/~M��t)��Bz;��9�E�g�n�C�Xմ� ��^�� ��D�;;z�FZ�4� Ɛ2#)�|���5�BA�h��R�R@�/{�l��c�G����94���Ďy�����7���[��&�%,D�B��Aj�B$��I��]�����s7X��E���p:!Z9�6��ud ��2�49�.G��4$_H��ft1L�����<���&D�~ n����X#`?&\�vWAN¹���#��h͢u0A\
����l�ǽw�g��bg?��Y��_^L�B���������������b��m���xOP�au�\�a���r.Thl��Y8ծcvE��t9E$�������͜��33�e�.�`��p9Y�*�1�V\�j{�|z_܏{�����A�����=�e=��\j�����b��;d���Ӛ&����"�hi�C��
����ڟ�Ie��h1E�&��8���:�-��d<�Ά�r+�`���O�m-�:â��mq�Ch]�.R�"�2N,\��g�jhS]�@�� ���F
�Od�bH��s\�Yy?��8����ۡ#�e�u�[_x/�%���_Qd ��̻���W�{K���Pj��K���H`�#g8�g�N}�˷}q%΄���O֨�l-�W :ku*�k֚�-�k��J�N,o������ ��T����p�� �<°V6�s���z|�T�f�Iں�H؎��4Ò�Γ+��1H4�m�a�Z�Y�YA�3d�C}�e�Fÿ�s���T�H��h����ܲ{�,�g�.BOJ0ф�����؂��#$���~��zX��ڣ�K=6? �F��9��$uSz�:r�tM9�����ケ����Cp�������>���b5e�Yϓ����8�a6�l�T#A�p�Z�l'�`+�55��!�>@3.ˁ�ŗR ,��ՠ�d9��0m��?=��`�����9 F��,}/�
��D�G���1�q-��Gc��KO�:���h;|rF�G,މe��Z.�F`η�Vr}�1�L�z��Ek9��&Td��#Nzr̊���*`s��/׆���]�X���}+������=�%@���8���f���$���r��w���I>=�
�	������x�߿���<H�ul��ͤ�Џ�
�T���=̖�l��q,��4�J$������HU�b��4d�Sg�h4Om�أ
��\ �e\�ށ�6f��)j>��Zq�'{��$�Y�)L|X%�\V�}�U)5A��ҪM.I�Y�K�f�>��v/:�I^��>����\u���n:�SZ��%��2c߂b�'�MN�&�{R��;�Z������[��$��`�YO<2��kdy��,�xɞ����p���H��\fT��{���*\��C:?�8��̃��np�5�K>��5`͹⥡��ِ9}���ߣ�~<��7��&+�ߗM=��~g|��sd}y���˔�'�Ô=�8?T/>���o�N���1��9W�D!v
5�@��]~�RBt�y�㴎��V��ٴ3�+Z�b'�y��<E�|l�u:��]�o_�_�a�[��&~�a�6'i�(�2|%u��|/����R#^|�_�YD���˞BN!�]p{��x�yrD�E�k�T�N���|�-O��m�9�4�Z�	�Zb�0��`�d�]�گ,vs��4���ϣ0���W@�U��u�.Uj��ά`;v���G��aЫ�@vx�@��(U�<�˳y����XgcV��o�0��1����h��%�����R�8�<�?��N��� �a[jދp�0׈�In�Wu��I�,r}D����+���#���7[3����<Uꂭ|�! � ���ߔ�摤9�"�H�OܴU1��H��=v�=ϒ ��1��B^�]�5���J_Ja߬ş*���ͫk��-���n@"I4޽N��	Ɓ_���ԭ�Et�|~'P���i�6ѫJ��U�;���[����x��^���?�<��@�k�;�%�!��w��!��7���y�/�O��͙Q�%�R/�A��^�Ρ�-0'w�4j3:Q��[��#� �=��H��CӨ@�n^�5El�ȅ�`�:I	$6[0�ᦫ��B[��'h�uRt��V�
���w�r6'�P9�Ф8����K1�{"*��GXa<��)0���ry8BJ_԰�R_S9�"t��UƠ��;11���
�R�
�'X�a��: ��7�Pef��;�������9����~�m���\��&�
)E^6��C�_5����Y��S-�Ūݟ �q��C��%�!�D!�O:��o)|�?�|bS�H
��[|obw�G�+�v�N���<�ќ�I�B��E^ i sv��.�9�b»���:���	g*ga�,Է�m�,[ۣ#"^9%����"JU2�W�ف�20�1P�]�݊7�6���ȧs�J��΁6)��U^.4a�נ��%�:?����~Zs�E��h5�SnX67ajus�D�9<���hֲ=�����g�7tG�f�d��X��i��)n��5���Ӌ5�#��lȡi�Z5<�%T7>����p���r���Yt�M�GL����D^��P��d�N�?�'���˝ь�7��E���Md�MÓ"_�������#x�Z�2#:饼����}؏�s)�9?���0�un�;H�
�!��/��	2�`�|'~롽�/���&5��u}�
�*�ǹKwȹ�S�tkYQ5�h�v��3�֫-��I�+�����/�ߧT�fa7� ���/I/��s��,M�]3�}G��Q�w�E8��� �3���@"L��m#�&{�Aj��<�m��l�W�!�.����Љ�!x�l�G]��9�_���i��[�	%�T�s�����4-��JE��uۧS��$e�0�t45?�5� ��*�G�S�uV�Ą?
�Sd��걆��s҈�&��j����v�c)�N0P�H���~~�L������@hẐ�ݘȥ��r��<�[\~�!�<��^�P�pF6kuq�`V���#_����2ՂhP�dp���A�x�5/�c�ˣ������D�������Od��M�дq��;?��Ҙ�
H�Hݟ�r�|_%I�{�;�g�z�)Ϲ��=�7dNc	��ϕ#��#sUh21i�Y>ڇ]?;B>ߗ �ʓm�ɓ~6^�j��G�h��6�[�&��~��QS��/8��;��f�=Ѽ���w�Oy���`o�\S�#t��M��l����ϐ��^n%Q���_'���p�!�^d.�6
#�BՊ˵���5��Dڍ�{hh
�|ϣ�������T�%b� =��a�#DIS�J�Q�b�i�N��znr_M����7��������W�E��K[��sַ3t&�M�8W龃����۩h�t��$��
�wR�.���yT�3X���*���P� ���6 ��ސ�N-	��Y�)��_�Խ���-�߮l�n�h2W8���3P=����^	�
O��B$����PJ���;(n��������O9r��H�6[[�:� ���Ú}I�8vnfZi���í��
��Q"U v"ev7=�z#G`���#�M&��*<�+Hq�[]��,A	��q�s>����^��Ҟ&�t��%oض�J�KrY�x�e��mP���"�|���d)oLM�L#|�&+�ֳ�ְ��̯�'�Ҏy ۓRI�,̕���m����q�4�t��
��tl;�-���D/ߗ�Um�*�B;�K�q��ݯ;��R0m��H��-f���2�+���9�����N�#�T�̩�E��#�m/�WjYc��9(�,N�<�(��dsLO9^��Nvg����W�̌tt_8J���Pɤ��	UWJ8�����I`� �����	5=
+�u���g�jA��.��YG��[3XD��u�Ū�0$u�<�+�g�-��琥�==B;�)G�F�B�U���z�s�r����6;v�$iaޠ��4Scw�w5�Ȯ)���5�A d�ȑ��X�O���m���=���ϊX�������P�*�#��yG� �ًY8h�cћ�j5�U�;4�U˻Q��쪌Ed����ge!6s�W��=��W�c�{�-#���E(��~ 㙅����;���udx
�; ������H���l�q���ep�#M�[T���H�n;($t�8��bD$�A3��/WБ
c0��8�}7���4��2k"db�qc��6vB�uѨ�6c�z+�Mκ���ynE��"ⓒ�X|����/-MC%QF �<�LXz�0+Vr)�s�:Y���J����%�.�h�η\�b�A�v���G[��9�}�!P�B�®�ס�-!�#1��s٬�Vs�v G���!�	��r�gwq�d��d�N�a0J�-b��[�^h���M�4G�-n�_6rG�)RL��L�b�lKhc'\�+ݘ�1�����\�,���<L�W]�x3ʳ��eGNS�ݺ��ElR��r<�����g���O������A��E��ЛD_<[�3��J	v�X.+I�/��p�}�vӓ��s�՟V�ҷ`s��@+6pYӮ�J���ȗh\j&��ͷ!�J�K����n�5V �˧������i��3��Q��M~�(��s`�c���+� ���!�9� ���W�
`y��\���P�j�J���a7��r�X\4�+��*a�#�v�E{I�ۈ�l;JaL�'6�)~�F4ص�Yr#�&��ىb����ZV���W�t:tD�Ncq5��;������ק����2����w~�xX��T��1]�ҏ����.���ط�TRk��]�h���f����f��۟^:�J���ʗS�^������8���R�Q��%F7.7>�ke1��U�o��,H1y��*Z*+U#0ª:�����P)!��v�o�V6o���xؿ=6�>X��^{r ��O��&~������ȃ#��3�:Z�25
v��Ғ0��Ԃu���/�X�r����9mH�?t��;��8��c�@�#� b,�>��0��
�Î)�G�*"XLt ��8�8]������L*2+e�n2�k?~�5���M�-�=]�js��a1�'yt���F9�%K~rr��3#>"�O����g�:0�ec������5\�3H�����Izk�Y���� E8�X4q,�ޮ��K���
|C�Lm�h\�9��b��k� �S�-'��_���BE����i��ʉ���
�v0L�ta)=
��ܾ��O���Y]Xdڣ�[9H��O�Cn���py�Es@����F o���h���F� �Sw��eY@u��d\!�1�\^K�#��% ��M��u��Hq7ѥ�o`O�+�Q�������f{A�I
ZH���@��L���{�̆�Ӄ��}'��OT8gq����Cgv�>�3�� z�m5�B���,�|���~Q�O�7��\3=��7
�{��/#s
ˎ-]a�����P2%�f��Uj���7���0F�ۇ۵�O6G/ۿ�ᢼ'/��ǒ�j3�Wj5zO/�|���S�(m��^0��\l�3eo����\4����DM3q�!��"�fS�1+
�RO��Z��g}d�翇�Xoi�Rj�_L���C�;w��J�4[4�t'!1�Yv?~>��b�����^*��n�wgX|�p5,*Lu��t�=VT��w�` ��}����5�z���v��i�H��%_
�,6eT�T{٦(4�x�5P�p^���j�P4vL����=��
q�_>Ulߤ�J�Tߑ"� s}�(�&p;*�� C��T���TK��W����aG��F��]����z���D��t�IW��n9-1��eM�2�O��㋏�/�[2b�h����y)��Gc��:ʌ��\���+�;��ᓍ�i����E[X�	|�Fb�p1��ȲJJx�T]Ō����yV ^4��L_�Ռka.��..�U�J!(���OflL31�Ä�g
tB<%���n�L��O�G�o��A��8��;~Z�]K蔶����a�
0�>�D�1�+i�|Rp���]�����NtW��p�>r���\��d������I��"��`�okek���.Vt;��b�qϣ!@�:|����	vq
��s����RCK(i</T�fme ��`��W�����|��` ��1'%Y�Dq��l��>ހ�-Z��q�PI�U�>�Q����Gc�7N�S���S�@�ſ�7mc�WI�C4s �iS�1G���J`Xw	W��O�Ӛ@χ�!���f���a�#d��%7t�������!�c�sQշ�Ja���+��Y	�<�������V��"�28#V��	�Ͷ��
�����+���������t�����DS2�O����>�Oqi&��� 3C6}�`6*��v�c~y��xfK2z���.? ���J�$���s�c<[F���*�[�D�9ݎ�F��+/�
K�tS�2L�o/'G ��k嚬����=�엪Í��ǐ��-�j�R>���#2�N���`O�A���>g;���s��>Q|�[���H]:���-�6<�+A�7"M�U��2��>[��q��AfӷԮe*��+iPMy ��!�@�$lM�N��d�]L<��:��C��%0�ۘ)�^L�[@����:?Mۗ�c��Ȯ��H��l�Q�Ľr1��	�jfpVJS�����T
�� l��J����E��̸oAq����.�f���J3<�2����2'i�k���+HT���'��v��0�ty˙��L�ކ�v'n��Zoڑ�����9�<?k�5fêA�@?��C���D|.tS�p�$&�pZ��F����zȷ/�`Ex�3j��Ņ>w0�)v�%�R>�z��6]�����p,�3��+s$�2��������GDӖ�݅�����^�;��8%���;�n���Z+Iü���5��9��|l�NR��ZtТ�sJJo?\�Uk⧐['��f��-�`Pp)��/+qwh*u��{�J�Sԏ�׺���ə~�w÷ׄڄ�d������}���7�Q�o�2��g�!�_��$R#G��p��qjg�sA�������gG����Wrā�A��XW�p^u�*�6�Y���KuXL�����\*o~�e�2ü�NӆO�9�ߟT�߳�R�*E �6�� �B�����Hȝ:A/I�ĥ�2a.��
I�m(�Be�@��%Zu��<���6(%bhI�_����G�MJITTG4�)Y�T=2�cJ�B"���+_ac���OK��^{���j]D���zO��x���>���#�
\�=�!G	�7|��|��-����������rY��Ȑ��);�{�zɆ�	��TG��S*�Tе �L�6P�t��e�y�R�~2w�`v}u���n5r���I'�ȣ"����|��.�0�����?�����ǗA+%�x�4�ľjs�,���-�[%�|�v��u���a��HJ���cCo A�.�G�Ň��u1�(;����H������(�U�߯$x�L+l����}~����A�&߹xGT�u+><%�t�/.	{v����c�[��h�K�-86$΃���Ɗ^Hɹ�YXQ��w~�dM1+��ňI%Γ�����pa�f�"q� �!cD����-�@X �g�*{_��-$�d$S�$�
��gR��P?�	P>���s0��wQX<����KwC���=ۛ��KUH ;@��� H�-b��	��HU� o�o,����r��έ�+�Us�� b~���\���VOen6NPI�A���ϰ~�/^�:@kʚ~M���'���h�ȝ�څ���!u�����!˘�_ ��,B����^��6�|�J�E!�Xѐ��w�D%!t*�7�c�/�ӥ���N�|��~.�W�|S�i��`�j�w�;�r_1��`Ӝw.�A_TȮX�����+\Tggq�tW �E�8���A�a|A�uB$OK�?�-�7���>!��7�����)n����h�<�o��Pi@�2��:A!e�*mC��P{`����w�P^M���5|�t~5�Fx���r��|{�u���d��ǰgʜ�Lvь�oe������A8n�Md�]]PYf���eZ������n�&[�n='�/����|�l����k�1��'P>+X|�R���vꘁ!?۴�}!�\��N�eG����*�xm���]3n��3�j���}�Z6��������}�!z��MqN����(����e�h��:����~	(5��+3�lc�IH(;.�����[�d�BGI�D���dmht+�ؘ��m��u4���0X3�M������)�?/���Ž���kP
��򆈪i�=z�L㡍m{���9@��q#-'.�k���B�Z�3O��C�H�|������HW@�� �/�u��1ETQ�ȹ!D��}v.6+�yh�����-i������������,5��/����	s:�zv4�d��>�6�P�}�U�A� �e�8�(�#d9�KPK䭀����3��e7�����u�NQ��1sU~-҂��6R�oӵ3�����\$P�g�*.;�Fq>y�$�Y~�+.���Й���#}��U�ے+oh�A�w��[Ŧ�%���Z1���t�z���̲�}���A��3bB��_}9-=�	��Kj<UYu���#�0��7@�k5�����:�H.9�=�-~ʤO!%|Ѩ��y��Aج�u��;13��ia8| u
���o��R%Rf��g	��$O�+�/���ߦ˄�ͥlL��ć�@�
� M��9�bu)�6|���~$\d���R��6TK{��ڀ#��뙦D*^�\������#��������ļ� ���PZe�ɪ��-N��l!�='j�Ls�ܖ
�1fːX���������ܦ;뺥)�U�L+�,ڍ��SA��ҏ�cMb,c�u�.^]]��'Է��.@ʞ��N��P�A,1�8O��u�`[�	iA��lZ�P��,��o��$�����l�x������Ӑ�\�P4ˡ�#^�z�=:��T���cR�KqW�T8h��a�)4�U�>��/�L����磹��#xƬ"��lL�nd��H�������U�w�s��&a�<��>�eq��s@7GM+�t(�=i-޸u�:V)�y�GegQ�p喎� =L��.?:Wz�Q��̨�r|JWjۮ:�X��}�$����1�^�w��[��S�o���J^��RU���%f��4E�����]�[*R�h� E���[���g�d�9�Pq9�:���R쩌�,p��fy��o�^�>Q1��<$~�(�.�X;���=0��ް��Z��N	V��F#YZ�z��D��p���*O؄�=���{/H���Pp3y��%��|��:>ܧ��t)*5�D�P:�I4q�, ���/������^��R�f[
0P��'�\�Jΰޭ�V'�ޓ0�xS#e��>p|�6����"c���
�ҏ2�|I�.�P� �Ѝ��E�YwY;�q�	�+��iM��%Yd
<1�|�R�{��і%�*@u2LGr�?��s����r��lF�L����a����v�坭\�^���7Q�Y�.�u���¥�`<q��#5�(�*�@�obx}�2�C�J��<�Q�N���(�T���|!���2�����@��nA�D~l1��|�4��kB���s�e��ON07�A9B�P�e��;tD�գ�u�l�����X ]��{%�\���h`�50�XJ����#�h�ϋm��>��\<�/_�����&�b:뻄��?�M�Zf�ܝ1�e��}�N�$u�zv�LM\?�7q��6x�q;�
����l:�㜛���ض6��K��� (�_M<�� ::P��"��K ��n�t������Z�b:d�de���~/VjH��}��&-sq<�+���v�v��A�����Ŷ�R���wm���C G�$�q��w/a��+8�^C���$��w�T��'�� ���c
��|��l��}iO�ON ��W1ɯ����4<���Ǻx�dD%~�8Z}f�5�]�as��L@���F����J���,b�i|�L���Id���DJ��#!��{E���� w9��+{��V�*���[��΋�y��1��6�H^�簢]V�h;�ن ����f�_�q�%���h��k��,!ϥ9���R�|M�v&m/���>d�#��Xn��S�1��&� -K��?��K��.�2���ʚ��O�=���kK�����?�����8��C�1�ГM��������=�*�g�nAv=��CБ��j�6����4]�����_>��*R���A3����ų��� �����'J�͸� K���~˼h�BQDbY8�a�g	��a .B�0SE�HM��WA�l�nsO��;�d�4����(\�E��V󹘾�c���8����z��$m���Y���̻:.xzDI�*o�Vo���^�O��Df�UqGP�b45/�HC�wq�Y�Ws�]�<�#�Ҧ�LA�W ����R���)�@(�N��q�v\�E�}]J)�չ��Hc\l���i!�N�n2�ַ�5&7��	�ʸ,�����"��^�)�#����;��m�o�tʊ�wf�93�(vM�2���/��ۮ���;�<N���߉9�����6R��R��JX�c-����̄����>���O�?��&���ٺE�ݍ�2�^{59�d<� �'�N�7f&��)R��+��8��1JY/C�E=��r�"��pF�������澖�BmK�%&݆�ֵK��Ջo�kv�̶��@H�A�ǡxcy���~����m�ߊ�����/�X���b�e�''��~�W� ^�^ڳE3���N��mG���x]�|�%��H7���FhY��H��c��s`q��HW�K�c''�4p�Xx�[\�i�W�4�����a|E5���_��a�B�wV��h�(�}�e]��scf�ʃ���Tt_f�,A82��Y�X?��|d�� G �v/�j�P�d(7XkNQ_�;�]��8�&���.���D;n����_��	:(f@�V9��9I;��v���]_u�����Y����R�O���)��K|S��W��\պGձ����d���r(����TՓ��8�Ӓx3PL�`�}�		��U���110k�Vo1�SM��c�D-�LM&+X��OY<T�f�9S�[C���տ�8�J[q4	��W���9��A�%m�#�0�2QV���j�'_*a��k�J�ʗ�mCGD{��6��o�S�j����.�sa�Y�8v�&пoS��0��p�e?�!����ݮ̭��R�lJ5���?�6t�[n��g����(=�B���bmJ��'�% ��ϖ�uS�rA��ա7<�\aM:U-�bo�����{����u@��p����;�.�K4m�U�<�t@B-J7����P��@1�8��e�)���H%k��e���+�����QH�y�wŭ��f����a����9�b����W��ݥ�fo�@�,��w��i�yy���ʶ�Y�U%¸���Gs̑i`)�S�|OQ�*��vOqŝ���8��ч�T,���C�q�;��ї�8��y|PW<����%x�k|�5��\��*`p*L���jߍ�X���4W4����(%�s�MW��Wp�s�����|���+�)1�o����ud�Q��w������h����
g����
:��a��/��vb	�!I��I��h����C��ݠ@:΃�}�^_�Z�;ʇ��[ϊŨ���:��f�:�����9*#��t�D���^��1|�`>��S��F�UՔ9.O@|Ȍrj@q�Bnv��-�^=����u����7ʘO��}|F�s�X��qv��&����i� ��B��4�����, �-U��R��O
���1��fX�vT�"�#,�oYĥ�������ܚ<88-gy��A�	�׌����%������d(��	��,��4�5w��`�t����s^��2τu�©��a�0g�����I�����o��p�M>F������J3���X:r������{����+�����mm�nL(��J]�PP��<���:�{i'-'I�͙c�I�3��6����?3wW��;��d�3�esj2�|���Kb`�p����K���1�����>���P��]����!��sU�"�=��4͇�^�s����Tn��K�Ã����l*�O��"�	B�VRD�߹��'jgJ�k0�n���y��h��� �hh�}�វƦ��u8D�;\�y��n5��e���8O���a��$��$K8���F2�cW-���j}����>(�HP�QEn��^?;��J�������E�w	�������+�n������L��ҵK]����۠����\�]Kp��^7�䟪�  ����P:%k����k֡�D�R�����0b2՝}!�Z5z�,�_��gݭ�Q8�$'S��_ w�=��F��u�l�'r�!Ns����"�ԥ���R������x������Ϧ�#�C�H������K�ڔ^���½�R��?��|vfĊ�@��	#�#��3dI܎t~�hn��L�W�Ow|H�y4s���Y�v��
�c�U�Z���Aq��	/qQ7D�h7�jsR�ɫjj��SA\�����Fd�Z����/\����^W�C���_*�_���5�1�Vo-S	D�!{�7���*��\�~����)�0��lιQ��ӝ4O�Ӄ���T��:��۬�������R.���j-��6S���c���LڑR�s=�j lBÙ��}i������F�KƉ��.&��ay+2\}����P/5�����
u���[�>�ߖE7�2�h{���e��	�D��N+/V�������삛hk{W�!���� ��햙�gve���j��>��<؃#�b]���Z��q�Y�q�j�]��c3@%�&/o_�ڥm�Ɲ��}8
�*�hb'�?�2�Lm@K4��4�ZL�0Xڦξ�w&Q"XwB�[�\
�#��%u��c�%M&q�w�������F)����l�ʙs�a���:��
~�{���-�n��yq%p��>E���"ѭDѣ���P_��d���l�JSV�*,e��s8]�C"X���G��۱sND�O�Ӽj�ȓ�v�����=k�K�=�b�$���_�A���*���g���-1��Y^ɇ!�)��� -_�v�g�z��)NI_ C��w��QZ�,�N����p��^k���	
�'�Q���ⅥpH	�n״X�O�ńj�m�;ye�l��𮐸'z�r���!���7tn�e�#�q�ֶ?,�1H��}S�5�E��w3��X�̍�o0#"�,*u��먼��E;T�C�g�а�7}i�y=3Z

��y�;�����ON�G%ұ�=�ö%k�?���0�^�$n+�R(�t]�7�`���Al�%��/�h����8+�e�nE(b�(�3�ǳ:��`/Y*�U�m'�.{hLd��Ke��o��no ���Z��I�������;�;�G0ykױ�J� ��M�(q6��9��uI��	��:+xA���wi�(�ˉ����Wr�`߱�`/�UKf�Q=U扈<k`�Q�G��������8̥��rK��N��8��(��|����NO�5�oܿ5��Tc�mh�L-X�
��_Y����:��zh�FOLU<���s�����ó�ҬW���'�������VJ�gX~�Ɛ��a�{����2x���t9�
�Cl/�x�"k�RBni`L���l�����TP�8l�7
�����T%A�������4L�f�o&D����ˠ{d1�	�m[.�!5��7��F�4�=Q�*���{���8R+k-Pd�t�̒q���(�4�a5�%��J]e��L���y̰d�\�QQ�ߙd$3g�sn}������/��#���6��5+Yv�K���C��}{L�.<��&pY8J��/H3w���ǡK�=c�E��2f)~�]S��IxT����9�9�z�aS{{k��t^4��i9iS̪F� ��1g�3��� ���~�Xq�󹭩V�(!�[�u�]%N!�ֵ��E�7�1�F�[�W:��9H���ݡ�}S僇/�h�m�)!]b]`)�'���UX�*n:ڄ�"�V#�J.<$`�؟d
(�L#�X��qފ��9��MQ��$$�F���a0ro��o�h�_��xA�~���Ei�$���p]�_C�ꃟ��v�O�L)��E�i��������Z��oIG�}#�:��7F~j��ܚ�K�T`��B_%WT��|��s�˲�Q��;�̆�"#���ڮ��QK$��s����,d^�W����(q�n���(BT�Ye�~)�z��Gd�Y!̅%0��!�*ki�띤�'�'t>H���C��P0?��~��R�ɦ�?HV�Z$v5%�?�8�V�}ٳ�-0v+/66 ��a����5QR�8�Ęm��W�lѭB a��-��%d�J�j��C���A�1��E��*1h!�1�=�G?��HP�7�0�_�?��F���o��ۡu/9K����L��(�kp@�'�F�	
s�o`�M�+rr�Q�󡒲�w���F�T)�P9�������T��G�@����NF�Z��n�D���	��sp]���[g�AC�B	J�f�3�m2xY��9P#p��b���~�4-�@E��娖5���c���)�[D#߲-�T��<���Ki�Y�c!��;S�-@�/�� Y��n�ǩ>��JfB{2IL8���a&�~!�����l]̔E����I��|��қ��/%�ܓ왍���"R
�Mq�zh�ݱ��R,p���:J����������0����s�ϿOS�����u��(�J��V
�ӳ����Vlt�T�����tW@Թz�L�����[�
nK7����1�#���T��ǬaY�z�z+e/W����f��vgi�O�,U!jC�8��7_WGA�	�,�s�d�Iv,��<�7���������͈;�#$4�o����Y�!E��F���ii����K������]qd�C�����(<E��36A}�p��Zu��Uj��.h���/�<�p�0O���L�SX!%=6��~i���<�E��j���$�Ђ�[�����(��� H�!�ˍ;�EY�H�k�l�B�|6��lm�Rv�E��#R���{�_�	)�f�J�VM&������|P13!)�r�=#��.���jH>�(W�\'>l�ɒK;����R]<g������b'g�^�ג򔧕�	dE+�����'5�
a�A5鰌θ��I]���Z��zB�����/-����]�󗹀\Ɇn�W7!�k�;�H��-� �pm����8�9
i�T;��|����A�}{�/�`e��NA��?n�j�i!���T}�r��\Z���ܺ+vP�8"s�L��Am���[t�^���X�c���1�H?���=��X҈qi�U��5J"��fF@�a�-�'Ș�8fٲH�t�ogN���wd'�.{~�9@����!*�:��qT���Wf���O�y�<:��������R��/���Zw�|�0OU����K����e�\VT����[�$�!�b�9�N���މȜ��z�����������z����ǝ"���3��o@�sp=�2� b�#*x�F�>>:��!e0�,�����8���X��Zn��}�5
��'�6�h]��B�٣�0��M�A�����)]����h�/ZI!���+���Ȉ����<.�D{m�9ΦA[���m �8�H�p���{��w�|��)��z�G�
\ ��`[;�u���^�bt��*����ʦ���cX��NC���;�]$,i]\��ú�%C��c��Z˴��Cm#/�Aۡw���XM`�dB��Y�E�(!�3�V�+젔�C�Q�����~'w-�D�z��j��%ظ�����'2��݀55C﹅ �k\Tc����b:Qߪt�����2gCi��'��Ҏ���T�±3����~	���LC���,v����^�E\Ȓ�Bmm��u�C��'�FBTKEi=�K�C-��DCT���}�
4���Ჹ��f���_IR�������I��mc*�o���s��N�7?����@�H�g��ԄC	�ٛѧ��A�w�sx�n'��w��p��N!S��$c�!EVY�×>E�V�VSP�������)�� k&p���g�ˆ�b����\��a����� �af*O!��9��˽䋭��q-�ټ��g/.�-.%�KZcv��<���

�q�KMe"c 7�d�B�#OV+���B[�<E8 :|\����5t�נu�!�M�D�I��!�K)W�NM%�s�*�]y뮆^ ������=�w\M�n�0��G<�����.�N�p�KzF��8��ٚ�6*}!������NL��Cb.�e=�Ț��㔕�,Z50H��H���RY�8���Au2�R>Of�獍�.9R�hEZѵa��S��O���=�h	MB��R}2�,Pٗ�m^|wg����5�'�����o(�/<��=Dt�O���6�F���z";"�E[��	��y���+�����syN >����{8͏x*8>m��y�8ڪ
�?D����<�%9'��%Î��[����$ˊw������k:�t�s|0�Q��C�_)��_�}�M�n�\(%<�K���?'v1���A�=�EF[��}��1Չm9
��1xyZ���m�I�#4_��L �+��� �
���bٚ������d�˶v��N`����Y]��h����'K��+C|�߲�+QV:O�+|���g���kk�	����T�]��1�5LE���!��M�,�0u���R����\݆�����t���!����*���=
�f��*ۇ�1}<�"S�_���L�gޡ_u����A�����ı#v��]��m�r�������]!��;�q+ӗ9��A�vc��H\&�%�(L.��X�qjf��ŵ~!2R�=KnL~82Hp/%p��`U;o��� Rb�5�T��>�v�{żѳ�ڶO�:�o��p��D8@����3�fK��i��"Z�eY0g�-j~���o���|�����'����E&i~��Zn�8;P��#5�whX}������P�����ᄺ����I6�\��i��j���wNo��d��$�D�:R}�:�6ҵ��sVd���CP�!kG�t�%z�Ƃ=���:��P��zSQǷ��.�7���B"�ƿ��mJ���!e����\V�t�"�m#@���,I�Z�� �%V�S����&d��&�:D��Z�T")q�:�t�O�^��0�׵�~�(_y8|ֻ0!��ˆ|�߾�M�]�ױ�b�Ό=�s+y�I|�����i��̻e��)�T6�X�n'��6����2ݗ�;���-q�C�S���[Nbɀ^�Lh�ń�~��8�Oz�M-����w�������L��h�Ӓ&M���A�.�<�%�~���:9aCj���o��>P��zU74�:����ݗ1/�o�ɮ7i֒'���C�W�z�)�S�7�)����Pr�!8q~�_2�,I����8��j"��۬	��3�~�o{6P$Ė���;�Oi���� ����㪬�a��,��L��]������ގ�x2 `���
bwX�߅� ޲2�bP�M9:�u�?���컸0\i����?�0Ń�i����t���@D�d�_� �.뤤b���j��{z?<3JV��h��%��U���+H
��M��,�oY��v9.���'��4 L�v��o�����{:��n��X�L����͊�M[�����h�������;�{:�w�!����/�?�}�$����79��N�pu�E�a�tFma�6:1S