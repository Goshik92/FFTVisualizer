��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,����j!/K���k�w˘��rV��d����`p�kv|^��h�����d/���@>]��bi�� f�<zx3TN\���^&�`3�w��}����S�w#J���RM`��N=��v�*��˸��?�X�t���9;�B-͜����#�/0M/'Z�xC�aUN�i�|��*51t�DԠ!!��I+���s�������5
$�g=a��Lf�l�j�{/���ݫ����F�BM��D 4�BUr^��>��}*���j&t{h�H]�[�f���B�U?Y��<�)`�:���P��1�=�_,/�eK�+i��1�#%�����j[�{�\5x;�ph8�V�jc@F�i���XHn[B(/@H�r8�,��m�8'z_,���I����~�.���&����b���B	Lq�(�NMUG
M]��m��l�Li[h���b|uy@m^��v�heШ�Ƀ�.�/�湾0k�y~-3e�z���S��Y��;F&.϶|�z-<3&b!�2����C�T9�Q��H�ɤ���VsF�q���$f�T��G�l���=�
x�E�,�C��I��M1{+m�՞��.�*���:>�,	QM��G&@��a�W��%n���2@�_�uTb�!�s�z��>�xO��\����)e�%���<�5����찰��_�w4f'ո+��� Z�����]���
ӛM���*�dC\64��ڱ�.�曾�dF�iBq]�*��:�U����� ^�+*�($d�9�(����Ve�s����uh�C�3�'�� :����L�M-՛���@�]�`Xǀ��u.Ŕ�V�a0����7�=��-��w�����ܽKWk��k1lXs��"�������ġ9
Bd��<C�&�̃DҐ�ْy�k3�k0�/�����g�߲
��>"HT.�e�N�D��	��s4�[��y�W�Vy$l#�UWr\�����Ǧ��٦o�U5̢3�3�����G�eǙ6� �L5_�o�vY%	��s�����W�p��V?�h)�nP~>��*�H��\�]{�,��x}��D��11�{nX"���E5Z��@D�W����v���X�Ut��U̷�f��~Gh��x�YK��0XU�	ώZ�&l��Ҧ{�����fxz��tVh���Y�H�����'�Հ7Ɉ�#����ו྿��z{#S�)���`�G����O�u�6�l� �9Dޡ���&���.�#��?���j�8xȇ!��ż�$��A6\xL�G�G�����w��/�vA�4�(*�Ӿƈ�5 yPnF�O%zL�:a��V�����D�)��������K�}�����	!��9����[pAм�_�� ��nr_�?\pR�Q���,<�j�2��J���S���1w��ǵ@i4\�rQ=���K�k�����p��U��|^|6�������G�V���L��q�k8_�P�gv�Ï�7)��Z�054L|��^�JO󾎽^[���6>��D�nm���=Ԃ��mF�=���0A��'W.��Z��˄���޸�T������H��I��0c�L�(�&�KѤ�vgqx���g �ūj��^k�t��a)��S��c���1�s�9I"��
WT���6Z��J��|@�vQ5����k8��>ώo⃨SNk�Vc�M����8��>�о�;����ܙY[O��C�R���+�)9��p�(����7��q�&?4�|PD�7�P�nr�d��dC?�k�eTp�!xE�R����GD��.$�i?�  Yc��a������:+nd;?�Ƭ�c��%h$Jg���p��#�������6m�~�d
e�7�˖�9C��,���9�6o��r�`ŉ�� q��P'h�/�o�|B$�Ǯ��^Q�������:���XOQ�o�E%�r��nѲ�f��)�Ͻ�§.�T�2����n������_���f>~B�5�}	ǟ��eZ��b�?Lhg�������e�'�<��}wgƞ����tR
�qٙ����k�Ψrh�L��84�C�^^�K���{uW�ɽ�s3XI�渋�
��:��l�+�4Eڂ]mܨ��L����K��e_�A��p�|ǂ
Fξ�x��o���)v||E���pbZ,�NNI�,n|}`K� w�N9p~B$\N�V�@�'�s���0�����cS�64o��'fOn�U�����R�������ЯŨęc�m��6���q�97
���9V�7$��lRY�V&W�ZFb�9mE���e��~�*Q8vS�g�'��6���:��WZ��x��|�CB���{��|N�!��o cOQ�V@�\m�H���I���:mN�z7����/�	�)"q;�Pb�q�
-(�i)��m���}��D�@�+嬗�k��,��B���D�w��h�4�<�B��pDS����T|e#�!�_��l�/�k,^��f�ݼ��L@&*�̇��VO�f��I=?�5!ڼ�㲍��'���b�.��\�	Z�Cp�ÁS��k��-\�l?��ɈJI�r����3B�5��l�̐&|�a7��'y���@�iR]�7�t��%O�l�'/+��8(�{�':ŵ�"D��)����8�<��O��w��� �\Dȫor�Y��p͠�R�(K3�,Ir��*B���e����Q����'7��{７@h)l#کh��|�҃ �;S�S �
����X`��Z�lP-�S)�?�ʝ�ٝ쨒+�mih����ߍ(bZ���Ҝ�����f���=��:kt��LӃ��z�����6��I�o�A�ȃ�c�78m�`�#��)���Lw�QǠ�6S��~�\i,0��Q�S���T[�`c�u��zɏ�e���%�d;��	ګ���jpQN5�Oo�A?�����Wް��m�]�����ro_�^-�>��сz*�nY����t�~�W�F�ڟ�?�/��+-�`�x�7w�CMy\�É9#DS�us�>���Ve�[�����kW��t�x&2���������;�B�����ɳt~�����I]�:�PN���O�K��`���Sv]}9�

���\��0e!6h�'s	)z(v��]8_���^���e=*�!>`�Z�$p��F�~J�������M�_¿ 7�r�F�FF%�r��v�3��z�f�jG�eT�f�8����H��WI�慔�mHփ�m��{ݕ%����i./���&�����-���;2�?0��!�=3���j��}T1i�ԩ6&��~�({�v��3��-s�{��W�s=O.��$���j��7����ᘨ_6J��'�����7������>uc��rܶӳA���L��Y�$���⛠��rLd^��{cLT+4d�o�܂3�Gt�eL�x�p3p�Q��bBx���{��{8Im�FB���v��Q�Fk!%���	��h �%��`�I0�Kw��؊e&.u�$o�c�=^�c	�u�����j0b��V�0�5t�D�1��(��V��~�a�t�L�g�!���{m	�Xv����c��y���UK)P
��Tu��0�����#�7������;gB�ϓ�S��$����u8ml��^Z���]4B
md��	RoZ��j)D½6.!oʍ�Tk|rK[�;���ouCjo7��n�0Od���9���l^0�	�4���P����Y���iɥ5�(`6�
�K�M�������i/�w��t���!�;���e�`e��=l���W��X6̺���� 	����0�1���D�7L����Y�v��@��)t��! ��]�ر���)��8�������9yT��fվ��|^T���}����B�u"��}`O%��:��i���J���)�����9#��+���?sV}S��Z���ǸӴ��p�T�LTğ�6� ��j��~}�µr`��"M4Z��J������v(�)U��lmiV��ȁ��Y�q%[
e�IvJ���+Uw�TĦ:�|�<$�$�T�`2�C���O���1E5��AY�ܵ�mL���!��OP��3P�<����F.Q���}���~�~�g�\F?]����T���
D�V���\cr��ߏ2��Yd�f����'D�Hmxy=�h�ă�}ț��*-�3�N&���*cf�ţ"��Le���Rl%5���6>+Θ(E��iB|'�8ptZ�
;�H��K��Ѡ/�TYt���W|L��}�jHB��j�٣����ȧM��jY5����[�=��?W�'�­-I�W�(�u������U����ūr���مB���5(���˛�m��A�CԪӒ���C{w�o���0������Л�t>�>����F�!Cŀ��&�'������RQ���I��^�&�\�2�87��1#����_}tq�G�oS�`|�?9Oe�xƣgf><�OӰǫ�dU��}M��j���T\!�5H�G��7l�e�T�?�������Q��
�qg���8�������T�XۍB*_�?�a��&Ӽ�ݺ]\9���f�f��ZnX!���NWy�`�o�{p��߳��.b#�r�ǄG��l�z2d�f��%��"�cwˤ���ZRT�{u6�Jp�~�YU+s���	ycu@���`�DR�f�}ӏE���y~�M�~�})���r�f�C	�����!kQ#�mc�L���2*�J�8��^,x��-�Vk6�YU\��@V�
{o}$��<{P���Ot�l;"�ζ��^
����K�A�?�����Yj��3t�L2��U�.���|0A*��[�����&dw4��Y@~uM�&"�yyE�F��&��v�2�����{�r^�&q�h�ك揽�L{�kd.�C�cR�_�l^�*�`����ß�|t#�"�;��S���}5���3���<��"�QD|Y2�^ �&��#Ā֢��1� �$@\��aޛ,d���)��)����}�ت��f5��/���Vl2^� �X��R�D x
_���U�����R4�շ�@艽�{Z��<�v	�k�����- ,�o����V�?p#]>��&X�>�xJ����d[�J��_��7Sh�l 
ɹ"�:#�>��%�)_y|�s�
�ܐ�tS�������U�\r�H�Q�'�ǐ>V�s�xu,I0�k
i�o��x.$U���ϰ��#�f7%���
t���E�j:;HnÀ�׸�Q*�gՂ�P��A05zl�㳵�;�x�0�v��Ōx�D��I�5�N��X
��PY<���D���$@��j��.c"����ۘ���kj.�/�1��+T����P�,z#���{;�?p���㪪��{_͟��B�,{���ݮ7:�lD�B���MdhI���lP���)ғ�7����FiR�iK�ln�PD �g'"�Ȱ�cB��ջ�5�0�{�Aú%��x�#a��@��(u+q1���y��j��|ݝ�5Ā	�3����Q�/��S�S��������0 ��;fM�t��V��$��Hb ��*
"�{�Z3VmżLԸ;Eaj��k\��6�3Ӛf0�!v�;��9`<P"�O�Hbe��d<�첸�LE��� ¥�dF���>�S�̋�ԫ�U��Y�M�g�K�BC1`�#@�E����e���}�D�4pcM~�{����wlI�-��rFsJ�^��� Ѽ�5��� hL��m/�R`�$�S/�P���2�8 ���Fz�&�������^��W#�xǘ�F"����CV9��Ǜ��ިU�\�Aς���e���.�l�zx�ɺ'����ٽ�)�FC�ߎ�Ji�Wt\�s(I�O�j���~�A���htE�!0��buPDh9q�������+�9C5�d�/�{V���:nJ��A\Z�����s��mY��epJ�AX�{��-%�L�J��q(玆��+X-��?!C�!�ۅ�Ǒ�Ak���.3����
<,Y�73��L��Ѵؕc���&��@^w���D�L����D,���qg.�%���^Cy�E����O{Q<`��I�Ye�*�ih0�>��d�L�K
�֕\{��1�y;�B{�`�^ �}�,�B�)K�A8���ۆӜ��;��SQ5���9�C!�"f{�s`A���K
=[�f���͘�M�(#HO��
��,ő�0�QsIO=��~g���ʰ+�]74�$�1}�!D�MQ� 6�� D]!���5PJ��ች+�|ፗI��������r'��h*�%G������J������ŁZ���w_,eIZ�����a`��u&�������{��Eh��+�&B���m����T�Hv��=s�Y�;���.�J��d� ����È�t�ޭq$�����ڝ3����ʌ��}��2�3�<tUB��J�c2����n���Aã�|^+�{��yA+Q3|�w��Q�'����^� �ӧ�K�<p���T*gL�m�VA0b���|��[�/�� �`U�G�_��~r��JE�N�瘡��`�VR��S3fA5,n��������j�Hb���"tz!m�ܙ$0��C���'\]�xH�&]����Leۆ�j�^o��dJ�����HO~��@ܰ���d�aƲDq��G�
)���%��YDї$�3�.>��A�h��������R�{A�nB�z3|�+;)�D���gH�|�����P��v/��ݹ\�Ŕ`�y;2�/%��^��"����$��JR��&8���n��u0����T>��n����|lh���mk��t?M�5��I�׈+��뛝iy����L���/M7k�Ù��G?���M&�[��3�n��Ǒ��ky�Ɉ)(�'L�=�G.'ޔ!��g;X�Ӡ�\���>������M��Z��xJ�S�j�9�����-�h��/�O6��pP\�;��'���沀�P�4����D��GK��R�0���Vi��(?�yYM'k�i �r���S����-�2��J[�j9[1iq��8��Uk�&���u�F�Ž�mR���Ԫ�����*���������K�ױ��)w}�?�hI���.�+o-#:|��ۏܘ:(?֬��;k��3�s���r_p�yEX�L#�`����)�1ؿH�ir����s,�m"� Wz����6F�j��*��4;�����)�8�"c)zQ�BQB�{�q�T�֎�Uh�U�l��jL�I$�]wi��ۢ���H��U�����7IR(V���ӂ��1Vy�ߟ^�@��9c1�αHj�X���YE�&�vYi����A^��Rf��Z�LYL�����s�=���3��>ĳis+>p�MX
I@���'dg��0C8{|p�R��]���봎�+Ta����nY�C}��~�K�����r�s�����$
�\��a>q%��Fn�h)Q�������� �r�3=Oж����:ek���8��?�"H~�C����Y��&��+��#=�(���S5�'�S���K ������Fǀ�G��R�o���DCD~s�+���Y����N��A���q�t�$dͨ/:�+*,����"�C�݅Ixpj��~:&C|���+�F�6�K����zg��,�3a?
2������5��H92��޼�����M��"�]��t��4[6��VF����vw,=3Ԧ��j�+�5z?�F�0{@w�\�(�S�;^;ܐT���������EJ�9;�{�Bfʑ�\z,��r^o���ĚiF}3Yy?${QJ���x����O|T˽kL��|�y!(3}�������qy�.�a9���-5c�Kz_b�RiMe�~�A�e)�7��&�T�UМ�)�P�08T��"%����*N��s��ݗ[�o�O�
_��k�B�ǿ
��fx[�a5�T�d��hՈ�Z�|�͓�&$��2i
6��Ӎ�bL	�� �gԜ|᥉���������M%yFLBe�0�9�C��0�����g�(����j<t��F�M�Z�&*���4������]�,�3W���D*�_�'�"��h����w���iރ�8w��S�Iu�-�X2��W7���(�Y��p�'Z��m̄P�/��G�������q �"�]�@�z`�+T�~r�g��C�V��X(Rl+���L�%ӱ
`Cr�/���3@�'V֛�31���z�t0�4�6j`�6�f��ܝ�*a!��c��x�D����� ބ^ݮ���΢x�Kԕh�T�S����֞wj6]�I��ʀ�!i4�UYuϯ�s��qjK�"�}��P�|sE_�}BDb��O�ʫ>�k��p�n�X�,(j?��0%&ts������W��~�q��-��_�r9�h��vP����R2lp�5���Ι ��<H	�X�8�ʃ���Q6�k�d�Ů�B�]DP��Ah�0u�я�<]�"�H"��(�a��� y�HY���/�5ܔw_���c9�?�9�a�Yx W�C�z�����!�X&��I�t��BpG�ԯ�!���"T~��7���������:�b�n1-�U��"jh����6�yZ�!�I@*THe�q�[0���i�°����ZA������J$XlF%�E��YF�,/�8�����an�x�9��u=�"6�+�Y��֏�!�':NS�c'i>JO�]%m��t!��ڞ�cq.���-�yIT������˱ƾC3�'����y	���$��
��ʴ��{UJ@]@H��l-�$��˂#9q[�k�{�pj��
l���<�%��A��AJ�9��w�M����5����'��8Ww�l�b�I2�a,�U�.�����gUC';��^����,n�Ѳ`����tmT-��az|d9�c�>�p�|ۡv����M�Rc2 ��'9C�Sv�mV��ۦ����O:H�y=��_����پ�q���d�<�OK�Q|BL���LC|���7�=�\v9.g�Bi^7?�m��I�G���G�S��[���N^��7�����oɠ @,��jDk���>�/qa�D����X~�~p�uCs�Z6��=5v�T;��l�g��N�񓝙y���m��������&)$t���%*V�y*��LWձ��찬c���[q:�sf��6��r��$%���i�wi�ul	��V3'�ȃ��>���NP,t[�� v�"�$#�d)�+�� Ɩw��>�U�p���-~Q���
�C���;F��9K:.���KV�hy����a���kؼ�85�c���b,�<�I��p�z��exGg�����K_�s�i&[�5��4x���|`:�t���Y;�%�( }���������L��w%R˝)����}F/�����7��i�(#�c�p�/L���<Z ��������'�b�wJ�ٛq������7��;��)���Fpz,�#�8��p�����m�['q�Ұ l~,�v�,z��R��t�%��Z4�|��k��5{3�~�C#��K[�ѻ̉(����֟�����}�VHI��dϋc	���r�U�R^�y�;��0(��� ��H���"�vտ�h���@�vI=�K[�'ӧz%:�i�3*��;0�㺧�0�I� �,S�	�.1���UGd���x+Y����_Уι�.�܋�\�������|��Mq
��E=�C�����!ߠ��$~~d�!V����d����d�a����B.S,DZ�h������2Y�M��c�/�r���ؚ�z���H���V7?�UF��z.7C0Z�7�^��/�/�M���!����j��#�lx�I�������#�E?��z¦�_8~%a��ގx��«wZ�.>��RX�<3�>f
��8�J"�']�h�G�+�������RG�md}����z�	�%Y��E${v��և�x�CF������VVcK��?=�P��G�	6��o稓9��uÊ�1}m;#S9`�����O����W��L��M���2��b�����4W�M��V�p�T_��%U+M�i0S���DM�m�zb���&m���9�3xt�[�_)�:Ǫ٬�t���R��)9�{����sqՈ).�j�G)��V�bx\Ocs����&/r|�u�4h�Ds�2�?�`���.eb��M� 9*����!ώ����Z���������<)�� �ī��[����/x�{Nϲr<Zoey�1�oJ����V{y"v�3 �@CڪU~(w>|�"#P@�!\ @�O<R�"�-e�/��'����-�5���f��ùh!I�#��i�Uv����y�4���4<��*J[�%�v���w$����_5Vo���w'J*��w��KE�~/e�{v��0>_Z��{V���%x��� b��>�@��m�*������?wN�Ec4��sՐZJ�"o��l��kn&� �^����7�ި�Ȱ�p'g�N���6�I�?�;-��[͉��.i��	��A�TkbQ�t��{��}�r!n&0UʼI9Z�xh�����O�Ȧ��w<�W���!7���Lq5�S.���\J(�?��!��v���=��\�>�x��`r�Ǝ�.�����r���M�@i�v��֗��YH�M��UE��K>~��`�l�5FGi8E�v�h�um�w;����v��6O�r�B��W@��m�A�����7��Z�'N�Q�����V�.�A�D�vϬ�?�1R�`,ն|(OI"�V�lSz"�%�[�?(5��W}O�_���,&?���u~���2�GT�V��s7d�&i�m1F���q��%�������ϳ�ֳ���> _��&HKF��?�[�����Q���4�0�]�8�V�R�|z �tC4k�p��r���.=VEʩ�x|�+���_�y7��)�D�Z6����:�Z�C�?�e���
���E=�����YÎ>�D`�mm֌����m��t���]K�HLs8"��D��|uu���;�?,H�a����4d�:��+�*�a������(ǰʬ��C�# =a7xSP#_��r����-���l������yB[�K�}]�kh�8F3���aÍ����`�N����`�H����O��g�"�B������I�~R՗c���8:�MHA�_8�+���݇9�@����	ff����^��-��?�E��_`�5v.��CS�3���o�{�(�)9#~�s�h&���1��{!�[��6۶�08Qke�֗M�S��;6���9O&n��g]�֍�7�����A�M(g_�C���*�"���:��Y)!E�1�K`��v�2�9��]aD���	��h�y� �p��aC�h�FBH41���x%|�V#�'�&q�Y�ύC6�Z@'
]d"MHGI��)\O)8������d���@W��/QFWqS���ҳ|eEP�|��U��������w�Y�5�^=��,G!��hB�7����� F���x\H/�h��'K��zN�B!E���2��(���?j[��9��b��5rP��\�q�D֠QF�!E��Ʌ�������������_�����'P����(|�3��h8UJ��H�����RT�8!�k�f��m���Vj;B�k�ZQ2����bwjX���^�o.��?�.�8���Ŝs���8A&p�ug7^+� ��\��"�9��m޶W~����ӹ��S�܇&�y^h�Ҩ~�.�8�� �Y[n���;:N!�$s� ٗ 4�U����4 �� }�Ϧ~�����;�����N����K�O�{��'�ߏ�I�4��rE �MP��Ei?z�����w7;��@U}�h�@\�v�H�uNw�sV�|U�#1�mD\�D� c��=8;&6�M0�_�-�*������:��VG�c4
�$k��eSpah�Y�	_:Ln#\������~ם1��4n22͸g�c�G�5�z$H��ٻٳ.��A�L��$����_7�B�p2�Rl�p���hV�8T�^��g� <$�2�ڱ�u��e~�Pn5����Վ`z�i�+eñ�`�n�'�i#y�=��ު�Ѐ�g)$1��*g�B��o����E��#NB(��������N�*s�N�����������������d���̞FиŖ�x�OM�Ҭ��"�QLq�B��LU6^a;��J�\(��`A��b���R���!s,���C��Ym|��*J�k]^ϣ�'#V/"�mFb�iL�u0�<�d��
���j[�y�M"���
!ѫB25�$J�a��Q�w�}\JB�>���6�d-�yϿ����*�%Xz{���n*x5F�[^"Vxb=�ܺ��m�e�	�]�"s��[��GM�Ӄm�O������F��"߬xⰿŧ�N�>���+�*z�]f�/p��U���Q��Wq����ڂJ�� -�����L j~m��sC�FW�=� �d��U!�20Uc�����4����G�1I��D���"Tt�R2��;&���6�9�'��7�@�F ��1��lrO�)8?L�{��ד	 I�~5w�H�	Vߍ��l�'*�^:�<�3��\�e��{�YjR,L�<�y
d)_!�1-��՝OɁ�[w�C佊��O�-X�ѵFz�����wu)�k���K�<}�?T���~[���	����M��>5����u�:��:�������T��]��C�Bn�<�|w��~� �5�V��j�o����I�\q����_;��64(� �%�a�Cm��jY?d=+�a5j�"�X6ZI��8�-Q�1�[�4�LB��V�^���?�-yiHT�u�K���F�otL9c���$EL���U�n�3YT3��e��.�A;�XL��cjc�����<�t<��t�s>?���hp�\l�2��=U�NL��[!�|_�U�t�I�v�>���J�o��x2t�W �H�aK��Z���j2�M����n��vO��fP�6���4vQ�7��@섳��k��3�Y��T��C�e�Hב���9"�U*���^��LI�~p�tb��k|�\��?��	��,zY-x��<Rw�>��p Nz�hd�%�ℬ�8��/�L۶j�ֆ{�%,�"y�1:��f�w!AJ>DeIX�����@�l�;o�������k�G��3{B i�h��gۉ��U!$`�1�H��e���J��j~�E����U��� ���ZۺS޼��x�;%�/�Q��XJh���]$p0��WYg��_�G%���Z���4��iѠ1��hp�Qm�-�2���y�ZR���ݒt���B���"��h3KL�	V�P=0u�����1
��"�-c�qj�y�Чi�M�o�����55(`�E4T7S�i� 4XL�i�j)R���ʐ�yF��#+ <2-���Y�%�V��{�|^��� �uқ�E�2&�����Z���(bM�+>���V��>�o�!a҉�$:�f@K�d�Q�@/���p'���ETB��b󂏯m�e5�uf��":����w�挥��nX?�Dݽ��`�+�yu�C̠i%9��a�h���>��H��]���c��~" ��Ixšf�����<E&<$�����q�i�(��(��-��Q]�6e��&�0�.
��_a��!������1xJ�K3R�����<�|bׁ:gM�I�E�)?�,h/L�x�Q�P�ҧ�E��]fw[<$ح����e��='$G�|��R*1�/�4��j����R�JER6�)��&HEB��ܑ����{ǳ+��.��V*�%�Sh�W���J�Wė��jUՊ�F�C@ɴ,���Wl�~K�4����ϩb�c��0w,��l^uF.J�/h�P��,g��Q�!����!��ߞm�R���ԍ��G	�s��tY����r�)���c�l:$5�.m���^C�>�ی;I��f���t.�M����*u`I���5��N-�xI���\v�D�l+@[�A�lՋG��15}i���.S�\3)x���8mqd�\�}'+���Qz�}�;�����C�/�7�ߒ�l/cy�0����U���Pf��'��D��o�p�*N`d���f=���ggJq�F�\�s���^D�-�d�5���_&�\;�$T�?���̥z��D��7�(���Ŷ��U)�����'�jq�3w}>ǲ`"�;I��z���-��y�z��[�}��*+�} m����e^��O�{��u�����~�Y��)u�9<E9��V�b�K�Z���FP��gp�Jxe��A���l*��\��������K-��w+�%��pwB-��ס�Q�M���:�]�WK�&����a�d\�8����q�C�� ������	CD@ץY<�(U��3�S�� ���]���gN8����M����L�a���(���;�\���s����	�4�QE����;��bl%�9�|�_O��ͰU��dmqD?{�k���|�y����.vL&���̎��q\�K�R��1��d1�j�c��,��;f��?�-�tE)M����Z�u@}��+�����Ic���Yj�n:�҄����	��l��ұhC���$7�#j��|�29��M�6RxtGJuƨK��W��ʏy��k-5>��?�mCq�kY��a���55���<�$#��%�2�,Sq���0��0�$]}��� 2HV�3���d���Bؿ"&�G����B�]w���d�ӓ��.��
��X�*���+03���#%&dz��e.�D{�q�u�4�YA�9�	"���Ǡ6ė���"���F:�����.T������q7���Lv�3�P�}��9�_�c�?v�āc
�A������"?8^��QH����U�`PV��W�z<��Rl���\W����;Υn��Fi�J����xM T*-�ك+a�/�6�;��F$p���z�g��s)�~����4 k�K�GY�z����,8���i�p�'�f߉�D"*/Ad٦���2��Yi���j�i܂U��r���F����zo�DjF�~S�L����7{�� %�ck�*7�ƫ75�U��3R�ݞ>D0Oӎ��\�Z�UȐ�-��(Zk`��2LO�3&ث����!ls���ft������b���)lz���h���v��6�N����"~��z�i�yG(�����*���i�{�zʸI��os )�Մد�����0�)�=C�"�l��K�E6E��@;�(��!�=�GƑ�	.�Xɰyq��|�4	y�v���<mn�uݩ4^{"�,spu�!6،?t����
+������۽�A�Ȗ%��t�{��c�~���dk�6�\�zM�Hv���dm�-���yX݀�����bnB3�8�T�dYd6�]'8�app����*8�}}�bഠ�]Bo�?�Ȫ�Y��fUD��4�5i��/I�z�U�nT�5?�m�3���Qg#ҁS�8`/!v��=�����6{ڨ�o��Zn8�\�ꌀI��MYo�u���%c�b�j� h"�OI�0pb��	�vg��m�ؙ�:ڈfGxs
����E^h)�V�	Nx-y��2Q�U���'%z�@�6�Jmy��Q��ˤ=� �Hbm�/�kX���9N�D'Ǔ^���Ƽp����L�W\��Lڼ����'��/9רГ��et��J}X�,Xq�j��H#V���T�K�!9%Tv������c�V3g����e!v��Sm��u��{���F�m���/�k�+15�y�i8�$:*�����-Ny���-3�i���dP�?��q]��|[73���}��S�Ќ�w���v�`�Hz������#f�����#萆��Z��e�<M�k����*���z�J����G��O�׃ѱ�f���T_;�K�.}+%�I��7�����m�9��>�p�t��ƅ��A_n����Y����~2�8�m��/M�he�5�	��6��������k+o�F���@�U��;i��7UO�w��	 #%�ۨ�_F
�^>5�hS���V�ۀC���ԡ0�U3�^Mc��n=��l�l��8�5j\s#6�W\���6܍� -FY�\h�J�ޓ���f A�Y8�*�_��8q��w7�O)C�nz��Q%Y��R@B��|���W��	�AysQ0��f�[r�1��Q���.���Y���%(��ܫ�=Ƌ/�[��wcz&
�Al�9*bq�d�:��G�
���i�PD�r��M�g!"|-�C��*�p��M���x��Α�;��ǥ�^-+�ںr��/ʈ�.����>�,�b�.	F���IKf��6Z���uv��M#�f�pۺ�/,#�����^f���k"M{S+y�+ݑiP'��KԼ�v婢�;�����}}�IntI�LI��(a7$k��]`�I��|O�
ͼj��kT/.��0}$t�2ȯ�'5@�$����Q/��<E:/4�]4����i��WC%���][�ש�?K�8��a�ZE�h~�	�ʰ�B�R٭nb;���v��uVB�o4����c�tӧ�O�@���$|(�R/������H�첋Nmkؗ�z�O��P*;O��t�MwEP笉K�R)Sg��z�����e;`��߄'\4������r��`�!�V�hs�-���಄(v�v1���$iY�+p�	ř�^��>�=C���r� �L��Qb�Q�eg��j�]|Ֆ��9Y`*�x ���e:Z=��DC
[P{�����S���O�g�U�,�fh2nm�t�S�~�w���~֢$��oL��s���:#H��DՏuI�bJ�DQ�t��Y��b�p��A#LÙN6Z�P�u;�"�.)U��!<�]			�n'h�:HVr�ѩѰ� $�y\6}��l��m���6�[z�L�)��J�f߃Zi:�F����x�I���i�����pb�e=��������o�f+�:���+��	�:��y�fA	�o;ZU��T�9[���E��e-�󸟱]&�Gf�K�D�L�Ε����s�R)if'��2�o*Y2����fy�%�|�0u9h8��,/�*�N������!�"sOt��Ԣ>�$m/hAc�,&�DM��
���	�u�? �^Q�����[��1��lq�4j}Fܿr���|S��-ƥW�vY��p�	Q������y�{����%Hu!;<�.<=�+໼[�*���o�m�bF�N�*MĒ��2��Z�,O��J�]ⵐñq��[����8i%r�9�M4*���)V��i,h����l٦}sh.@�#Q�W�����?�̿0j1x��ե�ϻE�����' �6V���AI���*8}��Щ�fB5zu��Ǜ��*�Š@Y��,� -�S��5i>|������f�P������r��kv�$x�C[�B�wĉOa��W����s �O*��c�1 /�[6�Z(�<�|�ո����"̂V���uA�U�c0p�(��w�-�	UzS�ŕ��n�����J��O>�i�o����JI	0B�V��,�vwWo7C<cy)V��T$ɖ|7�)�y��y�9��K,O���`$1�޾��Ah^�>aZ|j��Y�k%��Ub�>+Zf^�_!�������q!O�3�1���>����oQ}BA�3�/�-m����l�Spމ�����	�9���+�Z�����yv���D�%��w��vc@O`��EF%o�,9#�"��m'c	���ޱ�4Li����d-�!�K��p�?B"��M"�!�`7��qRK�)�k�⋝�Ze7W���Z
�<Ί�f��Q�,�MC�!u���1�B'o�I3$Ԃ��a�$��^9������#��a@�����UBȷ�YJʵ��Ⱥ�ʝ����35�p�d1>x�t��`���Y�ڠ	���}k\'����0���]�ex`�L��Y N5����M�Y(�C��#�=���B��[J �9hy��v�֟� �Li��E�1ȍ�{'�O�l T�S3G�ejL��K.1A%��S[C�(J�)��+�w�7����6�l�S��G��w|)�
�nǔy��ߥ~$P4`��3�_��M�P�����@(-Dz����n�-3���ђ���{�!?�p�{�$oeb�
O%#��I�P�+�7y�H2�*Bo"����` X��m�v�:��<�G_ʚ5�]y�ܿ�F���,p��������a����8V�F�6J�	����)Ǌ�t�s������k��x�(�[�} �z�DF�n�6h�����^X��u�`�!�j�)�xZp-�?���=��h�O�����(�cT6#C��vU�u���oJ��Y?��e��t�[7�E�`�b�ngf$c@�@
�_�?�
�c��	����ߦg�\�מY�n�jز}R�B�]!���= -�\��!Uw��#�F�V�AW+��$���5���k���{��%�z����X�ʜ?F��k� ��8�~������	Z9��Q��:�_�*4� �;{�m2�A�e!����;NUyb����Y��������efb+���c�=6���y�`�a�o��q]�%���D.���B.���ʚj[$IW��2s����Nyg��_<���e�3��nrş��t���Gޤ@[�_�(�g4��a͈��5�	2�/x�NfD�2`�`��b��Y��T^�C�j�ʪI6��֨@Dc����H����h;����H#�-7�H�:�w�:"Le�[ꕶ�чFUUW���g��OT-��=��X�ܛ��9.8��f��!A��sG�̝�Jݲ#�m�k�	s�V�.�A�����VY:�Ba�Pf�E�V��h����@��/�%�|Dn�-$�
��=-q�yS�)M  9��WE��b
��l~Jm�T ��������^Ĉy�61�J�W�g��h�^�Wc�]�?,'�����I��D0-�e�b�a3�0Lƙ�>vwf	�
v?ͲQ�L�����#%��Ȕ�uN�h[�p�	�2��d���6� �|'Vk����+���k�,�C�;�Ƿ@!