��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��/��Q�w���a5P��B�~�/�'̙���S{���^�qѝz��'�hřD~dVr�F�!5�=��[�\�bYzy��d�(5���*������j M����J����Cw&�u����Dg��>_�,��o��3�9=]�sn��5���A<�-��Y�,���AU�G���̻N�	�Ϩ�g�ϵ�w�Ω�k���R�9HO�o�u�(v�W�T�yVL �q^�Q�0/�����)1�cڵ�E
�W�D�t/�Ș���~x��R�X7�]0|��?ͭ�m׭��e��%\rN���H�i��8A(_�P��0];�ű
�0��F{��SUD����ª6��q�͓C��c�qֲ���L��I��7t8<t���8�Zݼ6�Y�$ ���
{ˉ��\�<rl��@Ƹ�(�m�)(q^���j�B�8pN��@mȮ���0�������[�N���s�!��L��u��q:B	  ���i)��a�E2q�v�j���GE�h*L�5~O���"9E-<f�� ����`m�d0>/�T�IE
�V��cp����&��$���R Y���O�}�������nA���n���on}>��o
��[Oō�H"*U���q<�%�;���B�m/�����t8?%䞘�V�6h���֚eU����T�R!�zFI���� =P�'yVrV�G�����a�&�|�)҄��PK��s�\��|{���⃿T6$��`Ee.$ͷ�A��CV�&b�"�q!�p�ፇ>�jp�9�v+��`-�H�Rc&�e�i~���c�Jq���'��`�q���.�����D喲��\�V�*Y��bM	D�H7�:w�:ς�|a���~Icך �E�a���(�Y`F�������r�n�+�hg��f�.��i��f�G�@�}��CT�4���,?`�g{V.T�c��'aF
:췧�G��Z��?�ӽ������#�ysa
n��x�2�4�mve�x��ͤ~���A	c��l2�F��ͫ+�Zޖ��Tff��iZ�D��7FeUY\�N�x�������%�u�^:d��gd�O�B�|��2�ul�8�d	s�.`7�X�C��\h�d����lG�%k&��O)��W�)��5�TH���K�@�F:,��׳q��h���Q/lϬ&�Wa(b%}�B��s�&L�(�m�`Y�
G�!R��zPV�"�
ҘZU'$gt��.��Kx	a�!{'Y��$����u �L���iR���jV.��Ɩ f,:��@�jQ�yi����U�\�^��'Z��÷nmv��j���H��e3R�4КZm�m���L�s����,!=:��q�T���iDu���+3��8n�?]5�G��Ϸ�h�<7��0�.zř��-�ydh�D�qs�gjȯ�$ZkU��/��%�/��7�ז�&xL������@�b<�!�,���~WTh3Śaԭ�� �P��XY5&a~��y��T^u�8��	;����W5ܚl1P���
J��Y�ؑg�70r��NK��<'B(bL���K�(ܗ��8�z	�^^ }>X�n,�����9��z�Z8�g����;B?���+t���Fc��+ۥp���}Z��e�G�#�k��Z&4r�� �{�>-�$�?^��
�_A�[{�+Bd�~�)<�gi��/~�o�����KZ�����82X�4VpY�$�]D}�+$]5ջ�p)���o�B{�r�j����2����K������J��v��kSl+��,��H�G;��	<��űN�_6��]�VX���k����[�̜MS��R���o���{��EY�u~�h����?�
��*-�r���*�C�1���K>�U�(y�D���!>��6\Ն}�3I��
"+}�'>�Z~;�߭��Eob�8��0�蟎����^��DK�VՌ���: ����u�ci��X����POt� Pi��[m2�,�����;�א��V��_H:����7�f.�w��-;*][�j�@�tҌ$����:5ƌJ�6�y7��W3Ł�nR�p�(�-a�ǇM"4#ڇ������z�W���I��^�����j��J?k-��B�	f�+ʡ ����5�<��I;[�S��-J���;f�|0��۳{7_*�[BX������]I:����ydhM',�6)\����Jm3�6���ARa���FK�����۫۝B��|Ժ���]�@9>q!ŧ� k`Ɇ��)@�+~��ͥ���F<3n!1�3篻�,Kq%�?=��q?uT�r qe��c�\����'�Vͺ��>�Cf^$t��b�C�����������/����Y]L��K��R�� �v�zG�T���q蠎�z}qr�X�j@�wI:���Ɋ��1��
x.���?$Ü�p�8^@�~�^h��V�\�g�D]���h�2�����X��D��>w���`x����q��#ٿ�%9i����&��9#~��.�n��7=(L�e�x�N��]_��R]r�@�Nl�Oy�:̥BCj>�WhTz�?k�2���R�W����Sk)���E������.n��R�|�Jctd�I��vR*�)N��.K�t�#�A�P
)��RD�m���
��|���9K~�;Q^H���9T�퉡<�����5|à0�-�<�!O�M붃n4P��
�pJ����B�����'��!�Ly`�#"��8}x�.Ȕ�)U�-0����j^�2�z �B��צ��U��te�����]�?-,�+�[�6�(��C.���}/J�j����6�/�,m�1h��/iQD�{�&�����nГ �ǧ���%�D�%닗�ƍ�*�l�(�w|�f�קp����W��^1���"y�>�V�ui���5�25過��n!)�X���83��2ú�r �l�jSI/�����p5�%`�ͦ��]Ҝ�f�0�~Мus/S�g�#CCi�2�-(���X�L�����%���#[j������{�\��4�t�[�@2�$�����,��e{TT�0�B�<�Ө�&y7ޝ��hLs�*]��V���,�}}O�p�lT�jya�
}�K��c�p��S��ղ�>��9� y��$�8�2���K� >Z9��<���18�Dv�x�#PL���(�:%#�?�{�G��#�����6ecm�TsK���NHST�k^�nID\�~��t�Vɩ��� k� �#�1ngec��4s�Aɷ�����{%`�!�

1����L�`_yʇ4�u1ɩ!)�8�}�lu��͢������v�Ŷ�*���~�ƞ2��jK�U:���X���uі�~�⓻�F�3j	խ)�A���v����܋m�v�b�������[
�4�bά.�#�c��a>�ܬ�ǧ��4��rps'''���Zs�B����F��$����m��juMfcW��FS-(G[���� Bs�Y
ճ��N�,o�I��E��t��k�13������[H� !oL���H���ltD�=�\�~�s��������n��S�
vZ���ޜ^ƚ��?vap�����b���d�u�D=� X��� _�<C9H�������Y��у�P��`7�H��9������i9��/�	%"�u��ޜ!��������Q��|�'ς�K�~�����N͞��_�N3���ї�H	�M�Yi����D=HSi֘��
�� �	'D�ܬ������m�]�H��qذ0a�#��bK��	�\�KY�L`O����#��9L% f�E�<1�JA
�J�&��ա
ujeI��G�W�18߀�l�%�q�f ���kR��ǫ�툁�S1��OM��]b��0PCw�7G�����&�؞�UiW��NC�
e������D��SnJ���MA���)���X�,�b�,�[��>^�ϩ�#�<2�Mfj�f��(�*���Dh\ r�>�t�qP��,���
��F�t�8�4@)���\n�]?�:?vO��z4!����$�����s�x]�u|���G=VKɟFQpvY��SS�p� 6ѯ�g^h�<yt���
�p������p�f,�*X�$AO���!��舶ʩ{�x��.�<��t�d��O�ۨVR��z�$ham:�dȻ~�=f����Snfǣ3�%/��'p�����A~�}H���].L��.w?p�����W�^��v"�n�J�i��ە�$[�祝�M�3O�6��>^�M
�6Y���]d}ڀ��W95��H����ѽ@u'z����E��y��6it��G/'�z���*vU,wj� ��:3�!�1S��˓¯�"�"�-=�%���s ���*9��q�)�Zy]@­(\PYi���M���If�g��\�_�r��'3Q ���#�l������*���ĥXA`T�A�A�lPX\�7`%?8�!_V<��~AU�*�ce�������F�Vk*�nj�q����|8�ģG�.*�sB���}4'%��t����_��BVN��۞6��]}`[$�b	��D�۶D+E�WE���[]�/%.�����|�@��.2d܎΍k~v��EW�ޚ�;/Q����fsr���CQ[�7��@��A�6���O��7hYsn%�\�1p��~[��]���L@�l4@����}�
֡l-�ږ7���f�U"7-�m�O��2�~@�m9��U��z�ܘg�.x n	���*
a�
K�)C��c�Jf��J��f����0N��$aA�9'���m8�%�T��,�'DWSr�hЅ���;�,�'�Hi���a�[�.؃�޻��NY^�����Q��e�&`���r��Jc�T��x�mb[�4�'Ū�ꃀ�JMp�����kKM��M�A9\t2re2�*�仦��ɟf�R��S��f	���pb�%��E2��u�d���!T��.�=2�B�COb88U��KH��>�o� ҂|#�[(e1(c� �U*����Ҳ��� )��^cײ�r:�������L����[��
j|� Ms����K)��)���4F�!	���Z+	���7-@�>ђ:�{�7���h���.v�A���d���V}䔛��TF܅$t8� 4E��ܽV ||������!
E"h*|�nϩT�����ݶ.|�����%|T3~h�f0����e]a�*���+�uqv�����Ӆ�v��4ch�b	J�������QFeT�^�y�;	�?��`�	5��M��m�$��	W$q����t2'��te~����q�>�#}���5W��a~�o�l���L,� ��X��=���k -���.���J�w%���\���]��6 \3�bt��K�-uc�4�;($�:�@�O��3�B�i2�
гNf�P	����W��XH8F.����j!6L����%0����T��Kd�|�,&^�2�E�K� �K����ۼ�^ֲզH���?Zd���a/k�̒�
�(׵�+v���n��JC��{����VӉ}�u��9ꘃ8H�i%�9�Fu��H�$d %=w���D��ۃ="��Zb����l@��]��e��E]��+y�s��>��-:�c��(�<��J��=��y`�7N!7x#�Vi���e�`Xh,N���B�8�l盰d��+���@�\s�� (��k��VWF�%��)-�=�&��hD*�Ԃ��+��ߠ��z�J�C\ �^O����è�Mr�%��S��uV>4M	����b ����%��ZxE�N��4��p=3zxO@#�����p�\s7k��7Br	��I~)���k.��!UL�N"S;P�v)KV᫩|1=�D�	ް�v	a�c�-3nE@C�������LW@����1�\2t��P8ħ�E�w�eX#�t�tF�w5�13��URc�Q���Z���M�
�����6�/�A6���%���a
iy�F}�^а�M&3���xr ���J��`�~%�J�����#�p�)4l���f	J8D�^���/`I¨�&U�l��^�C^9�_D��]G�)��RʘĞ�)�� eq�'�7���4re�6���.���k��E�۸��7=��	�Bꖬ�c��?~�|�ưo�a���K����V��U^g%��3�'q�M�̙���꤫�c\�|��Ol����q�hJ�)����)�X��t�>Ѕ��ɃE�16��Q������H����gwh����q�.�?��� ��UE��WFs���]<� �t�uSɀ�l��l�-\����G�_1d�Kgg��#���%��_w�A(�y�p���e��E6.��_����<��[�Ί7L���פ�����*ǉL0�M�>����-m�7���)Y������R��5bs=S������:�#}.�<�i_
N�2�=�˺A-F�l(Q�ꔤ�@b���w�Q]��Tex�PIK����M�4ԋ����t>�>�T����|I�co�j��&| �[Zbfc��T�$ǊL�~j�#��
6��a�Dߢ�}�h����8i�r�Rk����5ʖ@L=��}�vЄΚ�U#)B�j�3���:_b� ^�υ����Fb�tE�F`�P�\���S��/[zf�!/f��Yw6��	��x��W'm�SJ=�{�";*}dg����PT�L�fY^.c�1Lǰ�������_����m�\yR+5���n:x�Jֶ���ȡ
���n-�%S�GLMu�j58�с+f`�#V��n]����@7O�,�A.1\����pCd�2}�'^�a�1�0��/��o�d���D���������x-�D\(}پ�@��+��@$=�*g�a�!9�L6�r���;���_�3$�SV��~`ú�L����_{����(�o�����x�K�uJ 2{x�����M|&�wY��Qrg?_���V�C�ڏ�`#���#�����Ut�Y�e��*�u�O\"���J�'p���X�Wmհn�ۗ:�����Hٖ��.8������"Ѳ�)�U�3aJS\מW�~!Q�f� �)���o,��ow�X��`�w�@03�,�Sl]�cx��sUǒ������6c�?��r�5�ƥ�N(�-��{�-��m�Tʡԕ(%A�S�@���Ǡ�ވ��x	!�haϝ�*ao�iN!��{�]��>z���9Kt9VJ Ѷ\���(�C�1=�
�<|�O[$���t=Zܲ��9�x�j��j�Kqq��WÉ�dj��I%{�C�l�%Lm-d��@qV_�G��z�&w|���M�<=����7K��c����{����Y����6 ����5����3���i"��7�|�#���%uju�R��8�IO����gٞ=�zD�џx�˓��G��Ok�{a穸9��E��kD���|D�߭9y5*q�y��Vn�)h�3��|���C���b᭄�>�ưKC�:@���Il�&AtJ@�=Q�/����
@�x�@ݽ3��|��Ō�9Bwa�s0��/��W؜��:�T�oJ���GԨ�I��mvcy�I��CC0��j�۵��(��(��	y�a��g�Td6��JrN�E�A~�Y���t��������
ZXd���N��K�;LG��#im~���(re�`��."�����/j	=��UdF��LSc���[�mr�����A��*9¹�FKA��UCќy"BZ�n�9�Dh�N�J��ܪ��q�����:�)������:�1����̵Ju�5��L�dul�P�F�2+����� Cȗ�
k�,�N�\kN�ZW�wŻ(�N�bgV)d�1���,�n��=�y�QO�3 �"���.�4�����..��8w��k��ږ޵�G��e��M�t���/�#s�Q
�C8�a�}��{�^� �^K�W�I{�_
_�bj	&(�����V�Ĳ��H����g�)`�m��F�ȏ��v���k���x��x����3q��@���@ϝ�#P�4*��1cʟR���؉2.�^���jȤfr*Ǘ��0с�j�'Vh��*�Z�,<ټ����c��;��`��m��_��R����L�k�h�x�}nb�tR���5�҆Mnj׶�~�A[L17���˜�4j� �	�y&U��=���؅\ˋ5h�?�r�'�{�^�^���۵����s=�}�'_{+���"��CI�5���&w�LLǰPz�"�
r�
�T�I[Cuf�E��%z�Ge�+%�@���Z�O[,�иh�� �I�E-���7��+�z�)�x@�D񝾬�/c0D�ʏ��P�\/����ZE�d�e˞{�@�L��P�ʾ����!���9zffxw��V@��N#�����$�׳���w����91?ٍ�2~XR�  u�@ ^ZI.��J�"W\�+�|y���������v�ս8�F9}����C�����E�ٯ�@�݄S���U�����
�*�&I��l���*X(�@Fr׵?h)6�i�XI���(%�}�3�?x.`�Zю�*Y��;/������@6h���gC;,zy�푓Ċ�#Y3����Nۛ�^!)獟��yp��9!/+�{�\׏C
�T�k��o�9p�Q�1���E���څ����qB~N7���Dg��§:���[�>�Jݢ�W�+?x�i���MMN`d��P���v1y2�hAR����&�`�[F#��V���ʆ�5>���ħ\��h�\�<�2ԏ���'C[BZ�i����8�α��&�P�=�X��h�tuL�/������6C��U���*�Q���`��K�=r���֎_���Ԝ�̳��֓p4�I�w�M�i�_����Z+��ƒ�_J��$?��b��
���f���rݟ�V��3�)���-]7Q�I���	>�1�i�����z����ֺ��S4q#e�y����H��X�n��F5.��dM���+ߵ�0��T��\8�4
1`����C;�NVt&��ɛ9�����0�&K�}Z-Y�>Y��	���)�������Bɀ2�OP��H*s!?F�N�c����&�񯦮JO���UZQ+ߡ�b��?OżEѽFA O~P+Bй����T(fz�R��$���п��!�U6]C5[�b�O�89�2�r�v A������O¯�e�ݕ�9�su㭃^	J�/�`
�Q�u����\F�l��X�z�F����^��cy�D`��5��4���'GT3�5B��N�ވ�O���9��	�.�N�L3�]�M9���NvbɓcGn�k�2)=*�}�X�l=�Z�KX(f9;&nd;�	.�h�����iX֪�EY�Cp_N,n06���\�(����i�� ����6?&eV{���}8ݗʪ���?���-X��g>?q̾[�������'"a��P���

0�s)�!H�*[����%�X\)� =gɴ�+�����&�� ����*���"���@��CQtN����T{Qפ�z8��W%;K0��a��Ȭ�Tv����~.D��y��@�����nZ��
]^���2���Tp��J�'iu]�f+-���Y���bWy��U�P$�W�Ԕ@"�C��^�����9j�UA'^���ʫ��x����2o�� �D |*��	��)(^'�5��S����m�i��RP�8	"��p���(��6/3% ��A�'|ņ��2���s��B������t�s4d9ao�ݑQo�����c�&���_I��������,�fR�y�Q����3L����a:���>r�7-Z��*�/�_4�hC�R�S�xQ�Q+Y$�۰i}�Z�n?�~�0G<k׮���u�vG��(�z�ØՄ�[���f�*�X����^�} 
�cA���A&���x��AM($��z��!zuGa������xtVzV�\�A+�	5��/�(�?'?�H�}%g�Uq�Mx�\��m�5�	�^�p'�5$�kʩA�� �@QD���̇~8�r���摮�D��%�������q3����YoVΡ���)��w@��E�,݈^Qo��b�B?�s�"�|�CE� B�_�U�4b�+0�ĕ�ځ����ڂ����A�ላ�K�{��-�+�qJ��	iiק�"��-�y��*�]|~�tD�P�JB>�룿���6F��\���b�c|kHc� C'�#��;�sz%�l1���gW�bD8�~���p���(�����z5�������9�.�e��;�*L�1,�u�����,}���$d�#�P��p�$5sꢴ����*��������+�p�b�B7�z[)��0���'�;R^�40NC���>�̧	̨Ո��-������`8J&�0]֎r�a)A�԰>EY�&ꢄ]Ѫa��P*�K�{�1Z5�,{����}y�a�)�Ԛ\�G�$������ki;{�n�'k�^mM� ������ �mi�׀��L���
��X��9jܓ#/ξ�����\�^�G(.�B��s�����Ŗ���pt�y����!.�pzl�w��T�R�mYS�
��߀T���!��:FQ����n=��Z�
y��� O��Ŷ�E�+�Wd�z�ֺ]r�-��H��2 f�I��Α�Pqw!	����>DL̞�t=�F�{o��;��i.Vh���#��d�����ɔ����p�9��I��:�6+���.���E�s瘗�"�*@��������+��*3���a]��fJ���H�{U�-�Û+���3��3;8o6��鬒�`�0>b��/j�'��tQ@8�����F�I=�
�[���x�&Ô4�'�e[{n�&@�3��㉋�U�7�����Q0�{%���vv��ȉ�%�踿[���Ƕ4��T��9�홚���6�q���0v���$wW����|���1e�cP}NCV�y4iN	�CS��� (�s��%C��$5�a�7)|\;�BѬR��{�����E���F+ܝ>�-ɯ�޲�S?��c?��\��$��|�2#X�,�j�t;���4*Y?K�Z��}�Z��~%*w���`�O(ah{��Uq��s���1�E��S��
�Ԋ с�jU8O�a�p��l\?����FO����0n�_�E5��%�GNf�M7�l���� ��␾8VHu[���%+g5�N���HA<�� �AA| �2Ñ 4b�n"Ͽ�3,�%��D���L�Қ��r^�!��@2 zw�1U�V!zVB�<\�]~�f����� ��}Ǵ>�ݯ.R��t��U�|��f�k��A���i:��!���,8*�}O�Eg�ԙf���gi���0Q�_=h5drw	Y�V��$�̍��1xJ6��3p2-(e�ESj)��ǹXΔ����v�#Y�<���z@�Y��A�z��H�"Q��1�'[��HݺX��ō<�+N�F�ȔUl���7��]P�����1�!g%Qa���*I���1�~ |^���F��lНA�k�E�8BJH?�Q=��Q5���@�Z�R��L��p�xX�+G���q̛�;q�Y O�]����	"e-��p�YW��y�BI�I��S��o³���X� =�5\���>$�.�*�����$��s*��/6����|�(X���}�ٟ�ѫť�,�%�&+�M�;I��p�P��HsD�RW�cRX�
@�c�~���0�߅���.��)��?�ʐ����i��:L��9�o�u��k�'���Ҧ�U�w.}�]R���!����	�����Vb�@���x�I�;�:}�.*59ؾھ����y���!U��,�{3��o�o���*�n_=)��5�~w�-O;���k���4i��J#(Ȑ��~+��U�֮�o��^��z��b�*��+�w�Do&�b=R�y��E������$3��Dx�� �%[�5���e�(\��
�J�,[�&���STUPl��'Qn�7V�8	M`��JO������f�������n��e`��>�.��QTֺP��jr���h-�F��c�8U.K�R�#/G���}�<�9#S�w�4( �y�����UN���X��rr�5�Ɏu�^-��3c�"?\��[�r�]�i�����������m�#9��e�����O�Ϻ�,�
e|����>�O�B�2Mn7k��3K�;�7�8�z2yR�
C�4StɴF��3J��/c�mb`9�˷�����6a]�Qn*H�����z��G��� 2�ʯO��zč�-5/b�:�s��9	�q�Xo��?���Uȶ��;���:t���ac�	�	mO���\<b6m*�d���R_t��8�+y'?I�V��L�Ÿc#MN^wY�����vaz?��H��8{ Nd;���O�r$��MK��V�@Z�q�"�(m���Ʒ��U`���[��{�Q�4��ԛ4�p�w'G1غ���S��$��Y="��ڡ
̓�uD�ES��	1��H�����Z��ɵV��|�+��X�l-$�J�ɴ*E�V�F.����O�%��Z��&��.*���1f�T5wTCH��d^Dm:O�����9�Y��CV*���� �\�1֟,�"#�}K���\��˄껦�oׁj�O<S#�����M|@�$��'0f"zU�Z����ϗ:������4Y�H��6���X��g��te���$���5�k�s�zA�I���s�#�.	@2g7��qn*S����ٰ�fP�~t�IN4� �&/×܄.e�9.v�)���C$��]X\RE"�!A1�/��.�D[\�}di0�D+ �(��h�-�IXy�U:�w�D-|�(cv.�XNy�nM�0�b��͎RА�$�@���՟@\Q�ir(T��'f��y�| J�}����+;lL�ӳ0|k���d����-v�f5[���[�ĝdJcE[kh��)W�e5��5��'�j�uK����&�����Ȝ�Gx��3�[.���]ys��E״��f���:o��A(t��	�o�rWUR Ir�a �'ͦj]���A�i�h�25��{���r~)V�S��K�>]��������p"��WxõZ���Sʿ:�
u��}��2�siФ���	����e�s0�e3~����;������3�/�̱��Tx�Y�5�����z�G�h�����hk[��:}TÌ ԣ�]0 qఌ�܎ʭtc��J�r_K`=�G_O�Yk�f�)}�E�=^x��=J���{��Ђ}����>�o�֏�A'�m_>T� �����A�M�f$��_���^t���k` -�k0�����Q�=N�A<�T���(,��<qI���D�}`U=�э��k�K����g��HǗr+d6 ���}V���ZC�*�p�@����DQx
6r�n.�V���v�vI��4�G"�$�X��u@�%�g�fΪ��+�(a�Q�Jض�dv�5A��:j�dT ;s3���ʇ n�p���,�)b�Q
̄��O���MvA7Q$�F^h��ҏ~Ζ*YF26����(�g�@�h�nȽ�B#��w�Wm֯� �M���s�-�����s��z�O�8�5o�p^�Kxg�����iؕ�?�������~7��2[�X��s����}������J�Nd$w�����lX�9�H�np�ߖ_�.��a�]>y3!~�ʼ�̙p��_ �Fu�p/5���S�&24^M����,��t(WW�Z�<u��x<�Kb�4�g�-���t���蔬=i��,V
��~��)��ec�,�d47�Z�*AΚ7/]��7�;�!�O<T����M`0j���_�C�prgA�I�� �c��p����|��I���:�/B,
i��j�OӨЅ��g�8pȐ}���!v���J��Y�M+8C����ԧ
��J�1�_�׫Be���.�����n�ᵯ���R�C`�gS\J(3�<	�T
;Z��|n�!P��v(F�>�v�[�և�F%y8��k�}��#n��n��(�:AP}���?a���+Y�;N�Eh{��%��6}31�$�@���ѵ�Y;��i���]c�z�`�`�l�)���Qz�t���ۗ��3�0B���$dw�E��ӄMQ������Q���L.-I�x�j�Ɵ���hh���3�ǽ�CK,��a��Yc�G �+
����e���z�LV����r��Ϩ�[-���d~�FQ���Z�{$#�ѽ��F͎�� ^����0h�8�v�@(
Y�m|%To��_s^^�4^�V{$g9z��.�>��x�fB�
���,��ٹ:J]I��,K��w�BjD�5*���qf<H�L�˦��O`�.��Q_2�e�б:��5"DV��#�=�.�ֹڃR���>�:zy��x1޼�,����
�G]Ky�;������d"�7pDv���~2��X�8n��� >�R|1�e�ˀ��j�J��d�*�he�2�v�M�ٓ�%�j�+iw����P �^{�f���=��Ĺ���R�On��������<��㳨
���=��6h����W�f?ཅ��O�f��<���{q�w��V�E��=�9:σ��b̊�f=��@:s��A�˘�iz�quN��<��%2J��K8�;�4D��B�tK����@ϸ�ևs����u|��]V��E�B7?2\j���$W��B���C\U C.���*����Q"\ԡ
��zE`�rWVqg��1#f�t`��B�Vbl�:�4��/�!�:k���ͱ�Y��n��'����9[-��l�L�����VR�|�H.�eJ��[B������<bsx�u3��[lo5�Oe`~(�d������4F�D� ���E��&��3��JR/���$�D
�<�/�����ѹ����'!h+���?Xs'�x��ٷ��4���뛒�e y��QCd�D��s��f��y�M���?�5�P���;j�l�ٞ9���L�������`��43	<4J�	�lR��0�	PW@��fz�cX��n�h�	��C��l��#/0����Қ�4͒���-�9pxN��mť�(��Z���C�i��6�p�d�b�j#Ru���V@y���N�75�F�!�a�$��i�qgy��7����L�h������Zx8,��t�<Ȳ�J�o�k2�U-�����\��G
t^����������@.��8xڝ��v$�6*AI�����^!�:�u�C3�����W�\w:�|���X�qro8(�I>BX�d�8R>Le��(��*��LG�CQ�'k�H�nSX�tW
�"F�`�~�ؒ�;�'S֍���pt�����O�b�~a�V����9�+��� �!; w#�����+1�&۠��_"(/�t�R�?S�;#�Z:����'��	h��m#�45a&�#��K�΄�FZdD�tݵ�����;�W�y8
�ȑ^��X�6��i��V�n�����O4�ݕ���(]L��Ⱥm('�!t�Z��R'��;|�:ȋ����i��T���#w��m�^�������8�&Rb�MIe��1:_�՝���݀�/m!M^��B���nD����>f��ȝ!VǊTAd���ٶĊ���Qn+��u�� .��U���})���ʏ��	��<�t���<V �>��D9��$�fT��9|k5��!�W�`�um8$\d@�%h,�@��t�� �;����"��r&E 0�7�j�ԅZ{��͎}��k$d.K>�ۆUd�a? ��6&8������,���IL�h����_�\�d�哛���Ќ��'��T��2
���C�&�mh⌱D�Z�_��4��6h��W�Q�zHRj˗��-���[N��%Ǽ�	�-��-�n��na��JV�����p�Oΐd����W���I����SEAcՇ˷2����E���ާUu�4��)�ӄbDmJ"Fu�CL�L���8��!%����9U�2�^k��L�,�w5����b�J�Y��p�Y��� uw��[�;k�q��<�z@ꍂK �^���m���$��5�L���c6F�#
����׿���xW}-)�E��J�8gťI몽:����/�
/"R���Sm?���.8����#�hWV�	
>��(�;���F���k�H���0��|���1o�@�-��+)t�8~��/')�QRk���/�h�nT�`M�;a��$�h�-9C�Scg�^!�3�
qn5��}s���Ѻd���js3�D�x�&��fzh��D֕U���Y�5<|���ɴ�g���c���Vꋦ켒���-���N�y@����Ƕ�	�u�Q~Ɵg�j���B� �ܙj4f�G�:�}H��
���z��
D��\a�����Y�d��'�`�h�"C�$��6�f���Sy��j<��v��1.��Qy�J8'O*�s�6F�T
>�=T:Z�J88�I��������&��h�ͤ����VlRv3ۤ�"���b����_��U����c~	3�j㽘9c,�p�pu�/r��"�w�-X��o�Y�������� V8�r�tL�lw�j�Y�O��)}Va�#�@�{�֐��pf���<�Qؚ_�SyP���ZAa�Y$��r��T�V�ZK"5��'��lL�F{d�QQK����b�ƀ%�v�� R�m��Y�MY�
 _2��beU�f�� $A���$�u���*��}Fm`�&^���HB��PR{�#�����B���T
ⓛt��{]G���Lԋ$xZ �,q�:lS��k�B��`W03�LR>,�k9+��m=��x�w4��;=N�D:��j�'Q��d�[[W/�CR�L�-P�'+,��Q�	v�q!L��,�{��Q�"Wd�ʚ�X��_2��]��d�C���-��P�aY�&
$��T��"O�jX&����z{�W`��5��X��a�U��#��Z�Eɏ�u�Ѹn,߰��-"���]�)"�e����
?�	�s:B����HX"l?i���
��C��e���_�U)���6"�إ!��������=��g��U�-z3Y7�2+���F~�3{A��Uj�n �NkA��ܚ͟�lݓo^g�FȎ�܄Ue�n�#&%���`혴��zf�ɕE�|2�y�������4v�v�S/t��Ú%pj?�;/�5�*`r�+!C��G�Y^v�ϻ�,��9a�_˹��[�/�:^J�|2�$	�w�kA�A8n���c��0��KU�����p�<8mΩ��b&K��$:��<��Vht%��
��z,�FL@t��]��Vu�R#�E�\92Ku�P:~��z�`�M��>_Y@�m>L\���.���CI
HD�d�5y��� yk�%\։&��6!���S�]0Cr죱8 �����'�z=r�rW�E�������p�Gy������vi
��f}W'@Ό���9���7�z�3�ʸ�W�%?�a�I��vq(�u�<i� ����oig�R�R:�z���=����쨳��M��ݪŠ, 1UJj7z�	�� ��G�&@.h��B��vP#;Ku�+a�X�<~��b� ���dN�ۆ�l��u�qVw��X�Q\�+�lI+�*G����<���mT5��(��ER�!M޴ID�m.iEg.R�T\�fiJb>��<����v�d^�Q����./
�5 M�%	��3��&W��X�1�'x�v-h�[�4�G)ֈ^�U�)��:;�F�w+�0��=��Ʃ��_�wk��D���IlĻ��b���ID�� +m��e*{m�Hu���?0����0�.�鰀_Ҵ��GCnք���/�v(�!i=Q{��[tI�� Qh�������LeM����
K�K��Ba���(��Y����~# h������W� �?f�ڥE�w"�������6K����jQ.\s-�}>��?V&�%����"��	��?���I2�P k�<a��h���@#f�!���f[O�PJ�"���;����{�.��g�v�N�ICޚ�
b��u�+vX�d��G��Cb;m垡k�8��L�
��N��Mc��Sɳ6A��~��=�����8�I�!*�Wpkh7�`SX"�Q�F��e_Sݖ�V��lN]�G�p�9X�oE�B�����ŇhOZj�Q�k棓[`"��vڪ���&?6ɗr5�ߪ�#{�hZl.�~�(W���(O��߬������j�F�-6���nR�0�<���H�1�������xnk�;BE����a��iah>~�t�xBr7�b$ +	�Z%������r咖�U��X3=;%�#��N��}�p��%���Z�rjnB߫�!��=OK��OkA�*��`$�l�,n�}�כ�r/Y[�w���z)�Y������+�n��r�� [���̧��Vk�.Ɇ!�����7�E����	�M���~�iB�F�����QJ�6yY�#P]�l��5Iq�O|�L����kE�Lh�g ���А���q	�kЇ�x�Ac����Q��M���3�]�ᗘ�&Y#��1�	�a�tL�?*i�?�?���zɽl�/��5��/�6�
s��bޏ,�ax8��2,�%�v��f�l�+IX�A��M� ����[��,!&qMq2{����rW�a	�i�=��C�5�j�*#}^>�g��v�w`_Ve����w���{���#�:��9�Sʢ��C���V�������s�\gI���?�#)�_u�j3N�#]��7?>�YD�������t� �V���C�y���§nW��H������K�.$�S�J�v�Wu�3?^����G�S3d�/}+�;�s��#?8�E�w�'$�W fZ���8��.o�y{WO�`\�E�k5�&���X��
��Ea�#����l��۴M��;��~��������5f[z�M��~@�������e��+F���trE�Шhj�Z�/E��I4 ���8$&�$K�?5�6;��S4@7`�ټ\����L�X&�邪�]S��z��ᱽQ�'v���)����,/q�j:
��P�PUt��ݻ-�C� o�T��˼)�C0U��e	�lff�S��F�~�2���Ν4�����RH/�[{?�|xĶ���(-D��M��V��08;�>�1ƈ��?Ւ��w����k�zX'b M�,�$��_,�e�=m~���3��s�m�Ny�
�eA(���3�v�h��D��ܜ��dZ�%�Þ�9v��wC,?F���cb��u�@t\�����92����3Q����QP��G�6/-����E߲I�L��&C��1>Yn�O�*ޖ��;���y�����W{7*CF���=qa�?����l۰���5�b��S���u�Rʞ۸�㣈�q�j
ts�QaT>0�lq0��,�.t�Dm��F�D�}�g��E�P>���l�Rl�����#��d���K�PW����@��c��NfY���ˊ������m�4�Y�Z,Ki2'�fr��8��l!�"�V��sq�֝Tf؉.���y�۰���l*��s���#��ϓ��FB�6���u�����{�"M�j�`���`��n�2��a]�0 2�:���n���Ϙ�����&��*�H�QD������=ٺ�eKp����Q�e3(�
C�u}ΐ�V��"��=Π���,���s��|.����V�}��[��r�d�aZ_���0��$L
~kr7l��\l9ڳ_1'��j�U����?�;/��#鎦�P��}!����$���~�̂��@}1 |Q���_]��qD��
��P�L�� Vz�C��Ցn�׉��;�E2��A���;��i|>pZ�n��<t����T��-��WIv���"y�R(�%�u�%�9�L$��d�Q>p2��#STl�E6B]�&��1��n����}���0H+�#��\yW�}�/����;j��~�C��m�ʩ���Ь'S!��J*:	�COh__=+:�Z�"�};�Ӧʓв{Ւm���/ڿhD���W�����m�/;�:�#G7i��X��K��\@�r}�O7�Q�J.ac�a��#V��Ĕ]
d>>�"^i(�T�:=��?�����U ��,@��w{�y�n��C��=���R.p�89���T�-Z��4~�'4l�~q{��������^+7�'����m>�	!�J��9d��������?��_����r0Mʫv��0�X��(骒!Qms��I#����K��&�4K��%tH�06��M��=��{^�հf�wuf9��{P	A�dTz����X���#�r�\��r�	ǝ1� >�m9x4�ki��)����]�7>9��Ui�1Y?��+D�/!�g�ފ���C��b�7e<�z����!�7�BQ�Hf�b�ďܞC���;A���`[7��BK��X��K�7�e���..�X�}�47���Ң-��>D�5ƪ�Q@E�[RA�:�Q���	�j��V2%�_��Q��(����!��k��*f�h �v�C4�'�/�<���yo�4�?e������	�)�'���v8�1�K	.��!K,�י�0�/���89�PMV���a�U�#	\@���Jy-�y2cMS.x�J^���9vk����O�P�
��:y%���Iu�}<4����8�q�zA(��A�?|L$��q�,�|I|��:�LT��GU�m��<K7��_���U�	�%��{n�VuclݘB�a���{�^��� �X�<�;����aV�B��"�P\&&}Z3&p�˴~O8>p��Xb�ѡ��f Y���:�_���m�uh��)|0��DX�v,��f�*��B�le�M�S�@[v��]�F��/;8i�vm���獥YZ��u�OTvM�e4}qǝrE�Ǒ��m��g�mP2V��(���Ǝ�	���b����I��0=:=VG�(s����/��&7]�L ���ܜ�'KA| dm]����c�|�m����������$�1�lU�l�
����&�S�}�����ޟC�|p����e�
9s+���rhe�Lx��{�>)Y?���c��7,�i�lgW'��0�G�G����2a�>�$e�x4�xZ��W����8�kْ�Q�-��:�l-O<t[M���l��`�p�_a��:���&���E�Ҫ�46en�c�i�Y��mg&~�W�ɡ�s��⇬K^�QRi���U-+(+�q7S=���%Q:q���j��ͼ�����{g�b����qp��%��~}����g"�b��tj4��O˽m�Oj��cdt��܂�"��.h��n[��͖�������i����8���'7%�w��K�d�E��>+r�*�\���m���q3��~����m�_N��mK��䅅������JQ��;�+�7�\BP4��e������Wy�uy���fo�[E��n�#�x!��p�?�� iY4ZF�1lG1����q�j�.[Ҷ��}��K��O�]���^ �"���4��R��9,�5�D�"t�`���)�6�L��U���ԋ�xC
� O�|�c'q�Ica��W�>�ㄵ����R&?O���Ql̲_Ç��=\"�q�����k)�*�iy�q���e�0Kx�.K�W{��]u��|���y�猥��A-��ı�w��;�l�``�k�uv�vztGi-��g{��Nz�g��%4JDE93�\�u�W����n� �V%�J)H>V��y�3��/�@�Ҍ�r]<�Ԓ8��ɹZǕjיMs�}���#�E��Mv�6<��f b��v'��IJFj��q���&��Bu�%�wQ�^j�]/������6��Ȝm��	�ӌ���?6U���+�&���{�봌���]�q�̭�zyO�_��~��;��qDMRY4�P����� �-�f H+��hw����*��!%.��5���������֎7�u%���� ��v]�b�2�8Z=B�F���	���"(iQ}Ϳ�~}�w� H�����x-&l	�/�$`�b��)2i^ҊAA���6�ﱱ1Rl�q�j�N���$<ۭP�ev��H&CΫ ���l��+��{[�,��R�9�H�4��J�*W<�L�D�W�3~\�y�����R
M�`P������"fD��H���K^��)+��E3�.zK�3�o˾���(�����y.b�]���f[�Un�M��&f!��G�
��jfbW �zM�eK�[�z/�!�5�+I���?�|F�W0T�eG�A�������ԣh>�#M[%��z>�9���[Gg��Q:�CU�|R]����mԧ�&� �S�0b(���I�讒�|�L�5y�4��
@j�c{=d|Щ�-��M���ӑ~
WX���ь&V�M�|����8�I���^@R� �9�5��W�C��ԛ�k�<�[���v��]��}��!ŭ]5��!A�)4Qπ_��}��*~B�ݢ�f�
9�=��z�75��ܐl�zc�u��ң��/lĊ�1�3�ۓ�˱�)�Y�* ���.���ʃVB���!5����gr=/i��X�]э#�C�]!N:�aZ�F�l �]�k��'�D6�����!�<��T�U2ͅ��	�ag*�U�9�[���?�5&	��Ճ�~Sebd~J;̇ӂ'S/"Nդ59a�z�,l��y���N��&�G�su��`:tnz"�<�1,�#؞y�'�rmj<2���^��$�z���Z�	�|��xM&�.�aѠ�g�XEW
T��Ƌ*Fk.ׅ���D���v����T���9ݛ���4���ra��)7>@[�Q�����e��wJ���^r:��7���k\��b�;��z�Ú)�D���Ŝ�&3W�q����FA��b�,q�p���i�uR� ���! �Q�u�7�.�`Nkn"�r]���;L�R���ۺ��X[Q��Hf#��xa�P����`�����+K�޴Ψ��j�c�D�Q�8R{��u2��޸]�2rb��>c�ĶX:��C�R�<��bt��f�;.|m����p��Pvb7J_�F�5��S�Bl�c��g�q��R>�V�W����9s��(�.�)��n��ņ��A2��;��<�] ,i�=r��<@�T��MV<��U�H\�#F�D�����hv�����"F�LS�׷�j4o������c��Tk��	�໰5{y�=���	���(z������
gYN�@;�pUW?gr������q���kd���c8(���*� ��8�x����Ed�QSn�.��D�	L�%�r�i���~���Ǆ�fKzQ�8����-;��*��UH'_W��V��)�4F�>j��p�J;���̨ru��.!pʠ��6��yO�H3C�"�z5��W�U�!I�����al|�aC���pw=��)N�5^7b���V:�j't_s� !�\��<�~���e~�ɋ����_�@�V�c�& d�̊2�fR%3}��(���Y8��/lf^]D��Ôy"L :XK���+�nP���d��͆Qo��^�Wu�����Z���J-�gۖqv�Z�b� !vΛ��a���e}m��$��M�2����(
��[�9�Z;�f����n�z��k�؇�s��U��;n+��f!�S��RT�A	5b��,�q�*��s+7�����PA�HWlH��6�� "��$�N�}���^���$����7���Q�|�����
@������31����_��ne8�\��p�P��1��}��}�ië��Y�AO�BJX}���eNڵj�H|�^�^(�ʷ��>�gZA׷���c��6����̺fu�v��uv����T�_�n������B��A��$SRw<y�p�$�Sg�p{�5�N)�	���v���`U�fO^={!jE� E�g���9~;��&�:P"?��!��>l�c+Z�iG����ۄV�O��DD%�|�Ȃ���G=co�2���}�+����s��:�ȍ�C��j!����*?=�5a^H)�n2̔'���^(���b�+/�>����e�1Z�} i9s���'��u(�Y����Vw��_�`0)4a�Y�ď�c�Q��d�u%�����D&m[���x=_��CJF�M~�Qэx{���[JP�M}
t����t�t�4QQ��L��ص+f�h1�4�w��?U���*Kc'f�}�?2Vm��� ,V��V��t������9F#��q��н���br�J]��:�d�Td�]���v�JF��.7�[v��h���$��>i�=����)u���HgA�g_&D��iC*)h�C��|�/���"�������HL�:�<�z����W5�>e��>N�:�E �Ȯ-�_��`?=�$ Vjް�cG����a�}�8.7�F,���e�7�:}Yj*`���p]�p��d1E�.�K}�H4�����\ܵ㒳�goQ�6��<���s���a�MD�7�3�#�S5Xh�:��� '�k{�[�d\��c7ݟg#�W
���)9ˉsQ��wՀ�k2�����ؘ\ݻL�`�S	ґ1PN��OV��ÒLPe�XțuFp��-p�3��前�*�t@J*Y�ʓq��^6-��*}��o��k�א�"��t̢F�A�V~�Ȇ�
��� ��o�.YBIZD�z�	`#U@*�kI:�+���m�>���*����$�s9֔wς�ցOx5��uŠj�Y��|;���IS����T�����a٥�4��u�Q;[��U���]F�CfZ��Lw�z9y%�0^\��(g��_sE��Q�2h���S��	�����!�������
��6�Moy�e=��D3,�si�āK��Ƶ�u���q�
Х�h\h�Ie^g]V���1��Xƭ/3�*G���!�9eyg��3R��BT^48+P�Ͻ,�zܢ�=_q�7�� �i���� ��er��-K�S��{An9a��>���Eg� .P�\ ơ��9$���Z�/�9iۨ��6�oG���+);�JG��ݿF/FDwi�b���ή^�!�̄oY��q~��P���e/���.�P5y���k�C��� ڨ@P�j���&j+E�"q��sZX ,���� �J�	���dk������̈�2b)D9TfiF�ls|��[t"g,F\�_�Stm�Uc�ڝ�Z<p�8�:��n].ԙ����0�������B�nf�{f�ٱ�WXOO�[e�zImX� ����dXE̋�:6��7]��7�Ɠx�q��ϭ���L�W�sB����EڱA"��4e��8�
�BA�����Ȳ�C���	k� ��ᔤ
�H��$qG�<dl.{�A���zi�H^��D���p��>U�D���~��g�v
Y_P�5Vζ�\9B��b��/��
&}�w,XB�(��лl�2&�y�?�p��VߦGR��3l�Jy8ۛ���9#pQ�����3���῔Ik`i�~�M��m���� ��o!��GO`��p��!�j��39w��ݼK�I��q��6`���|^�n��Q4CB}���XC����\>���.�]�vFw-�j�9@J��v�Չ�;������1�K.�cE1�䍍}Q��!4xX=?OZ�2����y�>��*���+��fk���G�R���0�_nX�lpF<0C����V����4�k�������+�y|��]z��"��p[��A8�ft�̈́�g��Ȫ�"�z�I"�嬴K����x��,�
��� �^�����<���%�T����Wg�O���6y�)�~����x�U����@8&\7l�J�����P��6|���5�\��Χt��W�E8N�¬��2�A��]�ˣ�u����5����:9WK\�bu؂-a�<�l�{֪;�!Ut�Le�:#{��8D���c؀��l�N���%�o�+�iK�g����*�o%d*��ؙ�J��'�tڿ� ��V��5��ʯ��ơr���W��e����~�ȨW�]T"����ΰ���g/;4Y�c�3?�G-vphs1���#�2��kg������!uۍ�!�C�,w����}ܴJd�DH�@��l��2c
�^l�)�E��Ҵ�vm���SY�v��2�w�"�M��prh�xT?�*�c/����"֧+���R�<7�*��g�ADwj�/t�Ubh5�lh}�%$��0��?´i�ϓ���C��.�O-��R�ZQirL���`cZ��4���RN� ����b�%�I%�֧˚���za=H=�P�Ɩ��c����祋���l�c �-��V{^-�A�y�}����x�?���+!�Zd�BR��hQ���A���9p^�V.ĵ!6d�J�+��YnH84�en�]����N�Ҡ�:Լ�x	��c�C�F�z��w�ļΞ^�&�%[;�[BPK�S�V���)�q��/����)Pc�W၂�u0�R�#��UA������5;� &Z|���Z��b-��4/_��k��|͙�J��]hP���bn���׭�=-���|-bI�O�N�wMu��u3y���c��{.�����dbPD�ٸJ�� *
�I�x[ҫ���!<�w[	�0E��O9���͒�k/� ɘ�5_����F"=����ڜ�QG���奢�"��k��M�v����6[�lˉw�GP̄��JR�~CXz�b��\Ai2L��c��B}�7����MO�`/�@��� =��ؿGY����"\2�֥#(��L/jK]�gG���"���ۢkWe��{P�+��W>�:i�qdY'[0�����z"�pN���:�*U��Ҙ��F�{�=�#;�mdz�V�kZ$z!������P���bw�������ބ�;����������-Y���Xqݕ#��^�odK0�F���HOR��9�  Jk]B�d�v�������?�| }�Y�ʒ�|i^���M���H	GZ�Ci����P�?��Cow�,��M�#���.j���k�n[�;�r�5Dؖg9�,�Sj�ۜ����]Ȳ5I�B�Jsv��׾��{R�c��ݹ\]��>Nn{��O|�Bs�ZQnBW��G���U�V͒ro| ^��d\"Z5�1,�3��������`��b=����`�� ���;8���W.ۇ	��됻g�@��T�?�\; �zx�m0��.���j�`�H�aB�c6W58�_��p��G�W`(@ }:6)$C
�I��4xw)E'���F86�����-�ԁ7m)>�Su� V����~�{�0<��#ya�	3�<R��}Q��NFJc�p��>�;����I�����k$�=������w�e`eb��&P��\f�A��>�7�~��eޓ���^��G�X @�T0{!�!��J�6�����IU<}ǃ�V�+�7�m���]�����x$��:��k_�}���B��i� ����*�²�!�k�W ��P�::��
������K�g��N᯽Y��f1�f.��]!��0��5�F�/�����T��4�귄�`���f�_+M�Y\��*:����)q+i�]�_R�Ԝ�Ș��u9
�HmL�z�m74o��D0]�}w���Wd�NZ���
.�T��>�fD<JE�Un��'Vj�Gۭ<rE���P/䠅�!��#Q����a�-B��� g$>��]{�R�B�ϔ�C��ЅǒT �E}�������F]^�bWM�d�լ��1��\Q�!Q����`v�u�zBT�F�և(��z����I�i�r'�T]'�2��VP�s^�"�4_,��w��W�f�����6�+T��tIVP 
m7�(nM5u��4�X$5�d*k��@<�f����ĊK�vp�tG�vok���!��U�$*sy�k-�~�����hhK�����C����R��ι@��&p�w썹����6r5 &�]�i���tz�"��%�^�� �t��t��]�U�9,nY�>l��z�B��ӑ�L�����18��ߝN5�i7�1��y�|X\��Z�6i���l�7�G���J��By�]�1M��|]#[�u�����Qځi|"�֑(J)����nG�u��)� ��Ǐ��`1����K��]�VI�a�`�g�q2�-~�Faת��P��@��ੴEm�du�)�:Ӏ��j���8��m^�z�!O[���)���DE�����9劲*d�(�@|�;L*9�ӏ��t��1^o�^"詴����4Dp5J�H�ٖ�:a��_�p$����l��X*�`�ķc[������	Ɠ��ON%�L/ᨛ�r�gt��)u6?� I��])�̐����d�~�NK��f��6��v��'��������z��	� ��Jۑ�gu�5�_�.J~�Äx��t\uMt��2��;Ȯ�ѹ�Ouj�@7
`�AN("g0-8����cz�"�'��'b\ZX�A-��]hÎrj�����#Ɏ��Í�����m&(�jES)�ȟ�؈4�@�J��
lB���̞թ��uy�@')n�Q�a�H�iq�Db�O��Ÿp@;f�^�1�n;d�����}��8�� g�\xg<����>��,��8bY��r 2��V���J77Q�r
VХa�:a� �ZFb�&
�E�}����yn�=r?����`c�ZQa�ʅ\�i����S���N�Y�@y�Q�A!��<��q��A�A�!�Q�&/�ph0����&(���8�۰&�L��S	F����I��U��Y���W N:j����";��ĳ�LmpKꓞ���*��8}V��MM��Sc^BǦ�-E�;�j�@��$�-��0��c��v�*�^S��r�>�kq�OhtH��2P���l���dS��\45L�a٦S<�I'����Ȫr!*��RPr��{.��y�lÑ�1(���cU��|�S�#߂7o`<oU3֐NDI����FTiZB����ThX\s^���$7�HU9ʘT�P=7��裮=� ~���rO㚃B�kz��b����%��XBvǵKy�Pi�H�
�%��(���mI��t����ml��'w*Bij�W	�+[�|'6���X�	u��2z]���5z��!2�Q�?ne�ґëk�F��2��X����� �&�\q�0�e1k������(���&�iU0�L
�P�jʱ�tx��>=F �#�	�X)��yB6���/��x�}	Ċc[�6�~m�Q����K1�*��
-�}���>�T#����ؚ�.�|�	]�&�m鰳4�H�cы�l��6F�$}o6�P"'��+��wto2zV�%g'�	qz�a�K*���ZMe�ͪ���f}���!��O����t�]j�<�aW�&3h�\]���%B���<���FW3z�'y\�F���.��I�i�CK���9>�棞�����e+�)�c��e�M��<���A��5�8s�S�s�jpC�y!%y����g������"zx�T�g�vegv'�Z.�B�b���3VL��%�H��k��Ӎ�κI��=��!$���:Cޙ5��2[D�޺�z�H�'w�t�HC�'d�S�4�&��Hy4{/3�I����� LlK��9c��2�ʎM���B95��J���}��.I)���
���9p!��-%�{:E7�zb�S��ms#�>�8�ț߶#���U�?U��VƄ��(\�k��o*Yd`0v�9rf"���T>6�2�k	�t=�/�)�"��7%�'W��"�N�����	��F��Q����f��Pp%̢s�7�Q�u� �eq��Rfܐ=`bO���A q�z(K���$ǒ�T5}*���9��5zwEc�4
�}���dQ�F���`�C���{qg6���)�j���<\/���m��?����<���X��i���H.�K�E���?����+��d������,�y���1�@;�Xt��]5���G�8�wk��;�q��3��.~!�����c[��:!��G��A���5D�D�_h���Z��3���Ҭv����@i8�0�%���U�h�$��\��5j�O������~"m��]��:��B��UP�%|/����W�7�X��Ɔ#���JG�i����d���آ���&�#��g^..�Ì�XC����*!jH��䬂���Oݶ�r���5�jT?)����n,%*�r5/����(Bz*���d�����L:��h�J���<T���¨���3�T��y��@y}��O	 5*� v�
�-�i�q^�f���[Ox��ϒ�`�����%*�[y���/	��`���r�h/��R�gG1�Z��a䎏��D�R�!֙����C��H�MJ�>�±��`^�E��&Ɉz�(5�[)�*�\�B��|�]��L�lD$EH}iM��<tŀ�YQ×~�d�i��*��y�e��9��T>5�&=�_!���ջ����5�E��tWB�~�e���A�(���ū�Ɠ��T�=E<�U�2 0N�_-ଁ%W/���ٙ��2M�A`𥉙�{��wkkJ�y1s%kc�Ɯ�Q@�1��:j�Ǉ�Z��;��w����j����LZ��$���Z��tc��KN�F��w�xZ��)�Jp���M�:��t�c+szq7�
���U�G�// b�)��1��� >�[%?�H2z$i�F?�>2�kz ɵCm[�3H�˄>���7)Zuov���93L���,tk.˧�n�w��:U�ӣ�Ͻ(�ޤF�����l	��Ÿ�k�Y��bH��x,;�C,ڹ�����4���FKCH�T���Q�A�Z��n�ļ}Ũ�-��ZQ��B��|�r:h�R�Q�/]Nn��Γt�C������-������>���K�yZSis���R��9�
a��Kf�Bkq�B�U��;#;������'�D�}�	b�ၭ��Uw��̓�	�oB[��=[�_<�6����_�����ξ/N"4�S��Jfᠫ��Ê�<�͎sL�}ӳ[+�I��Xy��΢��mh��Ch|>�3Pgbn޲/�u}��Vb·f&���8n�рx4��s����k�]e L�G�l��Hږ��;uT؏0Äb��cQ��{�;�5�l�%���_ǆs��~׃!w��s��)�N���[��MsjQ�|m�c @��g|�?.�
�vs���E̓L�y���Ⱥ�_�4�i�M*���V�L�Zz�0mڧ��H]-�)W�`_�"@K�_�����=��M=����V|���l�G��VzU��!��,K�6�'X�C��v����"�`�[��X��6����xA
�:�~�+#_Z^ݟ�J���/���L����_�;������HgV��j'��8�B��3�Bt�U��&J,;&��4J[��T�P�
-��2�}�������=�e}쾲��t��2'6�)al� �΄�`�d��h�c��B����e+�>e|,q"�>���FfR��.d��Ys��\�\^�*��Ji�����[2���(���{w�����i��ϔ�j�Vݱ���|�b�v
d9��w�Z�&�I�R�_A(`G����0hT�]��MM	H�Et'�]�A�4Ǵ���=J��%V<ʼB,i���=�à�[e�_C�B&.�� u��6.]��,��l#j6U�\1����(�@�ŒU�����������k6u��Ռc�JL@�Աa^[����]D/*nI!�������.����v"Ủ� ��:���YZ#A<5����ŕ���j���48c�x5���{p�n�k��存+��m�nA�����Mt���S$���/^�<$�X�B������pSή�:uT�����46)�'�������1p[�x�I8�Rj�c�e���U_�c[��x����D�wj�:�m��T�
�4[��<��b���� ~$F�O�;���h�p�껃��6�h��ש@	Yԏ�v⑔f���1d��;��}��B�7��D�����M��(Þ������b���IJ��`1X�D��ϴ��D�5�O5@!#y�]���y�c%��Y�Uba�"�����B��q��O��C���N�_���v
��޵�k�i�S�ѳ�x�0w�m!}�R��MAM���uI�FQA�ݎ���;�sֳhnaR����A����6�])F�\�~�׍��N��j��|�A����◎_B��m@Ӻ� ��b��}_Mo�!6��j�θ�<3��SGN8�2�%�X���U+!yaug�i�M�N �p@9YK��6�u��t+�!�e`�-<d�v�o�O� �F"8�_ϥn��r54�YC��GP@5�aDe�I+;�w�--�T�@[�z����0�t��x�_�R;r�?V��ˤ5J��|I�u�Gh�r�u��.}"tj2xo���"�eWC	�L��~ɚE� �ɲ����Ś��S��r�y5���r�@����}_ύ�L�mZ�g)�XR?A���R-gOI���rikGf��U�6x3PH��;?���qL�0y��gDba9��2|����\�<I�$�&�R�`?
�Ȫ���xz�>8N9��V 5rѺZ�H=:C�2� �1N�|�ݎh88��O���� 6F��rR�FF#m3�R���S��`KN7.|�j;y
yc��so)� 51���U3�����z�\ٴ>��>��љC耘1��&I�
��A��T<��$��f�b��°�m/*�V��"m�9��X���_h)��L�Q͙����ʗ�Ta�,r�,W�i��X��^b�����2���
'&���-s�qE|��|��#EpR�m��'��P��Z�����Ά\H@�Mq�꠭��x%��7�?mfD�~Y�c	7�+2{��\*����w����-���=/|j棅2@M*o�.��]	�.;gV�l����7��V;������e�L����z�Ŋy�A:�=P���J'����=�2���% ��H'ٱq`ܽ|��o8���Ȼ�*N����AwaoLD�1]��x��[�9�����`l��������GI���R��!��ރC��J��Vd������0�<�!*AL-���E�_�_(*�d �*a�-ѻ�OK/���щ)w�)S �����A P4�ѿ�%G@@WR�^&�p+B4|������Đ^u��Yoe�Hg	�^��Y`z�j@��b�F�K���2o+	�_]D/od1>�?�b �|������5�o�zcT��h��0�����`������#��<ql屈zܮ7��wՅ(�3�#D�2m����?����i'B��wҶA"�������+� ��yg�8��u���ӫd��q��)/w2ǫ��+��h@�E�p]�?
����DE�3 !����IgK1>�LaH_P�e	���<7?j-i�|Ef�7����3p|}�̟��q+Dd�;,Rr�S�⩟pk�}C�z[�Q�:?Főt�c���S}�#���0k����J�i��jh5)���w��>\�
'�=TT��,�]�r�k�|@�NV��q�<�u�N�ɻ0��䵆9��2����: o"#�� ��d[ �i+g�����Q�}N[㹁т���;C������ @�?sJ�#�401���Ѭ�o}�s�M
��G�h�۝�^�Z!Ӳ����ݫ�j�;%B���=A�*U��C�A�[׍�@��$�g�Or9�K�9ůSE����f^R�8(�$�
I�e~�>����0y&���K�Q���&^j
�8턿�x�����p�.;��Q��~�/�+�����`6�k;��48�M0ٮ�/�O���˥I��x�"�Z����,Pj�W懬JID�d�����c���ڞ�1��E@E<�W�Gɺ�&��5f��`�
��Xy����	��ցǃ���|f�m��dp[����8uA�Z�rݕ�O{�f�0?s*�T����a�@���uX��y�F�=��й��vՆjb|�:�:��ui<�Κ�Ւ�R����&�uA.��$L�K�=��I�&˼m$ͯ�}ߊ�2x�Bh���Y��#-�|	��<�`�L�����J�2����MFd. !�y�l��H���7v^�BRg��,�I MY�<���G��k�6�R����g�v��� �5F�]FL�1!!��g�E�(�1����W��	�'_�J�ef�b�u8��8�d_�h����n�{�����7ӹ�c�g�eC�5��
��pK���/(�ԥt�xq������;0��l�觌Z�E}Gp���ЈЍ�z.����i��ث��d�8<#n��O޺@���f9/}*�C�zRI>�ld�p	�[�=���4�X|�Y��H_���cw���q˛�ݪS�U�9x�ܿ�Tt�>��2�#J��e�R"QкM т����˹�&�Y'�l�XQ�)��W(�L���i���P݂�	?lYx���(�mI^�b��p�c�L���t���R�����~���{3���9�@��p��\y1Z�U�A��̙��������뱞�j���Y���GH@�>��/m�5���׌�爘5�$WJi�����X�.1�ֈ��(���Tr�wBBԋϾ�Bg�F������V����z��� ���8��Ȫ� 	��U��D|���<�فZ��/"����:����8�t�X��AT��&q���Z���!�Q��q/LpR@\L�~󓦨bD)$��S�8���-�C$�E���.�phA��H�*���tE�U�/�����=q�@�P]���Kߚ[z-�hm�;�O��~O�!�%��[;�T�t�!%�,p��j��wH�]1ߞ178�vv#��T 7�/�����ڝ,)����p��㚊[Ű��9\6y{��8�Jr5�[/М���g�������egJMxe���.�������=yB��<T��u?�Џ���	oAR	ْ|�<�g����>P�˭������m�'�'%��cqqyv?Ѧ�S����9b2�n��q���X� �4;��!X�}�K��]%o�EW���GɄf�֢[ѽ��O���MyO�Vv�5-E��<�;��6
����j��2�?c�<�AO��{{U>+텎�*x��3i%�⭋���@%'����<b�\�����R��;������~Ef�vx����;�D�R��+��)T5_mo����	k�d�p�����<���-�k�������,�Љ�/I���<.��������浂�.9;;uzN�7spȆ�~�日����8�]��K�\�>�5М��2�7'��,��匞�sHZ�SdO�e���y�GqM܆x*��ꛛ��2��g9�������iS��D>�+Βf�Э���������A(��O ���rŔ�A)%�D>������*�oMg�c���6�h��1Rߘ-NAyO�[kC.�)��ּPyp�P(Ȱ�M�I���p%]��&Y�Q���H�O�L��%�Ts6ca븕1�1���Ӑ���?�x0�~��>E*֔�"1�;1�8!�N���-hz�v�-Q^d�X��]��d�oDS �2�$��+1m��ph�*DK-c[��╿����o��t�8��s�3�Zt'�Z3iy�U({�b<�N��|!ךU�����3;9g�#O�M)��U|�����pRV��5:��+��3M��vz��H:�&m%���,����k�~ؚ���(O(	�;1�	~��Q�s�W���|���),1�'S�.=`��6�t$X��y�t�*}Wj,3���U�ȸ�W !�N��ە>��O��b�:������=�v�S���>�XbZ��3C���:96�
�+���2Q�v�B�vc�.&إ������-��Q��w~ {���0�<5��J��͵d���S<)���:�M�܁[��̫�{+F�����p!��R��E	��U��{���������W���Ar�7�*��I9����ۤ�)	����Q��8��r��TYZ�+�˩7 υ�֥1;o��p`D��g(�Uz�Wcq�G+�X� sqzɼ}�mH*��3�@�JY����4/����=��Pv8{�sq��3$�6妴�c��n�Q���@�gܾB㡮��������z5���A{{M+^�Z*'� Mm�΋i�)��h�0\hn72�+��(�?�k���p�xW�Fm�*{翤1�'��lA3��"V��׌���F�9��~�����[�������k�, T 3�7�Bn���b!���~C��*E���sS	��:���2�"�$ƾQ�Z��2eK��b1B13��1*Ǡ�����Y]�!��P�?��^����d�a0^�&#�6�<�D���D����
�)"YBj[�&��(]��>A9%�-t�,|� v�;��vo�$>Jց��Q�Wb+��|�⓵Sz�2�ۭf!�֔��h|M�E�P�x�����<k�X�`��v�͚�\���;"#���9�ES񕬦/G��F<3�,��x�>\�wvW}�N��+�1��~�꤫�zy�����@M�T��'I&n�b�tm��y�|.��UГa �� c�-��Jʉ�T{�\��F���?v'�G�MMb>bo	T�FZ��_�|��+M�o�����<[���f{;l&�e��`y�[�w������E�s�!��V��.��h�v,i���f��'���߆�@M�."���Q�؛��4p�����	&H�6��.2/ Y�0��S�ñ4���Ϋ*{�]�}�?�(�ϐ�*����E7�#Y���2ۗ>�I��\��r
m�o�x`��cfD�ts �05e6��+A#�w����ҙ�WC3d�(��;����S%od�]7�ڐ�mv�㤁=_��37
t�)�3���=S+�T�qo�y̼g������	��~��MZ!��j�t�4Z-v����hKLC׭�gxk�E��(��=����a�Y+���bZ0�U;�C�Pf3�R��b�A� /b|)���c�Y�u��M�x1X��\�+k7�R/��Rm�⤶�s�l"��P�	�cHXb�_}����b��U��9���jnĕHv�e�Տ��SS��Z-	3�
�qT�J�◫K����)�#�v�-��LѬ
iUz��oQB���W�Y���4�_��i��7���"JQ.@ʮN�5J�aA���6�-�`�!���+��:m���|�C��g�r��I����6rY5�����M��v'�O�yǲO#��)�UF�?wdyO+au=�9�����Dw���Q�Y/'�eר(G�6�I}a�N��5�|u8KU=�H�?[&K����S�8*^��X��Z�ٚS+�Oq(���Yq�[-�
�&�s���FV��̈�ҿp7#1��OP���p��\������X:(�t윘b���ɬ�U�f�Nt��+=�"!*y%d��+�/���
�"t���N ����F�ސՒȈ��@�k2\bn~�V�?�n� �5RH�aQA}�:�0sE�� u�P���ͅ��~���R'��l��WS��v��lrf!�>9g�Z��cw������e�$��Q4�U���7���9	?�Fc��ݞ�x���[��FQ����%-z���̝�ɜj�������Ws6�8��"?�\9�����[��U�p�+B:�.��Cr�鉈����)JY�Έy�Z�jMg)�m����6��\i���S�+6����}�%J��1��^��6�.����C��Z�,�d�Y�X�U�׊���K�f歷'�!]?As..t;c���z�����᳾�H\�ِ��eSP7ۍ�������z�"��_e�08gD�l��QbU~�j�{W�~7�Բ��V`K�E�\I��|O�i0SM�r�rw�����<@��\?�����h�r{F)���(��QmK5��̛�6���3��r<��#�څ��U�tQ�j5�v�) ]�N�	�G���
�$��qlk���E��nX�ѽ�۟U�w�~�Dє����R4E���[B�@�=KdYcg��qO͛߻�q����=���g��!�#X�t? �x J��������G{B_����?~Ӆ "�+�m��xmy�gb�1�k�sk��Z(��
{@�����C$w��C�w|�}����nDC��A��\��H԰�vJ�B�T�"w�(���0�<�ͪ.NBL%��%��ڸ����k�� ܁�r|��-=�g��.(�!��'�m��B��'�F)�q7�G�#����6ŧs)dP������E���UU�<����'X�V<���lh>Ӈi}��ކΧ� �22*y����P]�nu	(:M��M�8w$���P�}u��\������=�u�S��i����ʧ|̚`M�2_�A=����،|P5�Ƃ�ln!�F�gfS�'I�Z�-h[�><H*�&���I�D�E��
�0��X�����C��V�ب���T2�=f���#����Aq~��ʟ�5� ���ֽFᑾS���V�i�S��ܙS����>ۧ@�����Y��0>|���PT+b@wB�ǀ樯![^W{~~k�R; 46�!��#y`�q1���y^]}�+�]��%�+�S��t���n�go%��t����YmW��W���?�Z�\\/����[8�	�Wb�@��L����߿=x�r�P�۟�n���&�(�4_������}@�#��FO	q�Xp���Q8]F�+�?�,X;�y���j.$�[kV %����a�#W� ��w���u�r~�)5��^{I�e�=�XPf8IT �^W�Y�BQ=[r����vj���h���������$.�Z��if���Þ1i��
IMU+zu�g�Q~n�x��b�b�|#��ܣ�ƛݖ�R�w�4�|4<�sȭL)�� PU�z4�4�uҽ��x��n�����ߖ�_��9>�ؾ8�"^�J'J�0�nK����ë-]�U5JA�#\���r�e�4��x�95B���=�qB�f_	�z�@M�'ut������e������tT�	<k@����V�Gn��WF��»1!v��SohD��NP��Zb-�&C��m~�B?�����u�ջ��-�9��8��S�� V�E1��J	��}w<��H����M���eަ2b���~�]�m��(#KB�o$$���B�C�L�5���դ4�6��.yU
�CCM�j�N~���c2��b��i8tA'{�SB���B$~�/Ey�K�m�dY�2���X�B��Y���U��3�F�p_F��\���g��"�ԁ*48�k����+t^�#���ն߫dW�8g��ל�kZ����g6�?�8���Z���>�B��[��TÕ�U��[t�d.�rf�]�Tw2؟� ��>:@����z���R�IQ��
T��,ncaY� � ԥ�Z�|��<���	Z�j
=>�)�	2�n�ܪ~�u^@��W�K�Gj�=t��7�Z,��օd��ۈ��N�wu���^��l»��@� К
4�nb4����U���B>�>�@�`�ǖ�A�4�&��p��)��ѹ^	e.���G_Ѹ�� V`���䙆k:���;:6��u��`��}�S
Hۤ�	i0������ԣ􍠰���sw��h-m�k3�d-;��[�L��)��y0����IL�~8!c��Ձ�`:@F���[�ܷȹ�������D���\	�ЧFﳭ�\�H����a��	g����T��,v\-�GW^H�ۨ$��셕G�@9O��x�2�.^���vD�(4}�˥����i%f��ON4�B-��5�Ez�����'6���-�\	q���		ʡ�L��Hq:�|�z�3�aW��H���
�>w��;���+��߮�}q�Ԛ�:��ޛ�^ث��Bļn�l-a��P ʪК6��Pץ9Ӣ� R��hC7_O��׸����Q���S��R��nc	<���Xi�p� �:lA�	{%�\��ufG���Ώo5����J�\����c8��xo��Z��&^
RuU|E��g��%�r����,Ӱ[�����S�V*J�6�����q u�.���)�co���_d��8�:��0��FB�I��G��N���ȏN`�W����u\O"}�,w��q�Z[R]�I;?�GA�
]�Wo�h/�/w���8�_���0m�${V~IO5����b�M����-;E$���h��o������g�崈,3���vۑ�,V�t��7>z�c]��j�u?U],���%�gEE�?�8�s��ȹ��b��H�;�+�IEd�?7)�U���\c��p�ë�lS.չ8<rs8�) �:T�y",e��4	b�S�"��2Pbώ�)P�`6A��4V��z��ps�24:(�T�TF/���Pa�镕�@�/q�����l��'���g���9�� y���j�-�H1��&u�mb�~�4O��QՁ*sxr�,Q�t�&��+����v	����u]aK4c�:�]���܊����ģ�/��x��*�-���&�:0f�}&v�j
��3�t�nAN�w�;.h@@G˻8D�r���j4Eb��e���u�m�L�ݻl���Q��c]��z�c�����É��3	C�����Bw��1=��?a��[U��1�O�,;<,n��=�޿C(׫J�k��X'\�7M��m� �
:6]��ln�v{;g& wlr�ڪ#�}�����er�N���Y�ي]�y��PU�����+�!R��=5���*�s���,)j����LhT6v5ݞ$��.ס �33��\�=T&Hm�"��`���zKX�c�j'��
7�=-B�c]j�IO_ã�3T4�2F3oU8qA�_3�A[�0BJH5��C�%�Hr��ȈA��-4[��b��'~�Ǜ�δ�AOM�2�|?��Lw�\Ŕa7�%������}j4H�E޸��&��*fU�]�Gǲ�R0,�p���[JT��dGƔ"�2Ӎ���0�����m�r6�6_Qf~ke /.͌����֡�ͥ��Ă���6x��
|���?�w����n���Y���ͿZ��?ܑ'�>�/�����+�J~/��>�P6Bz�LjZֶ���ۛq_^������sv
�3��\񡵄��=��K�I��6/ƙX}���I�t�qLd,ua�L[��!*��6[VO������V)=��F2r<�Ë�;����>��VA5)l��8z�I��R���2\l͂�/��L#��������@�N}��4U�ٍ@���m_J�&�DC\�����Qڨ�G��~aq�*���]����I�Xg��tp4�Ow������~�'�e���K���ȳ 	��Q�Ӷx"~�-[W����c'�l�=��-s�ifq1��4&Y��	E_��q��� �p��(���9�v�N��M5�=�Ё�9�:QN��hcw+�/�D<҃�\���a�N��q��1���Su� J�1rt�QX�����B"r���$Q����T����)H_�(��0�8�᫡�����a����!4O)��&O�����<Tk�+�NX�K��`"oudO�T�m/�v��a ܆'aU��������1��\��x������h^z!U��B���+E��k/���77�C�*l�)���:��$�ף	����bȓ��K�G�oػ��L� ���k\<���^���?���|��,W>�7A��s=�����c@o���~}��+s�#��As�}�3�]�E�	f�*L�>���r�:
�!ă���e
��
�����_ς#��a��u�!fx��*�
���9�33S+ �L:cv���ʠ��v3u�ᶹ4x��Xqo/�����ޗD�7M��p�8���6�؝J>�6t�7z� B.:��!�!6��
8�>��X�B�r�S�O?�tG�����wq��흤�שPë��A���(5K�C��&Ra�ULI���elt�W՘�@���L��2]���#�6s�Ve�_��ޫ��3�1�=���#=��!5�)�s��C��(�װ&�4�kNn�+
 I�+�w�ǟ�b ӯ�x�r���r����=Tg
l!h��;�\��1n[�Si<]�P���}��Pq),��fo�����M]�?ו��"�~��^���8��NՈ���#D�\D`���5�E�C�n3ԟzVG���Q���%9~C��c����˨�b�� '{4y����%Aou3����4�p	�[�
2،��7��E}�pغ�w�M­	��8�e�� ���yv�Fo���j#��K��I%��q�$�-p-]�d��S�T-N�9
�D���Π%��!���.s(s�p�*����X�B&�S���2l����#���-���	s�ڑ��4��xV,�c�FAՉ9WI$!Ř�7.�{��Q�"��ݰ��\	' ��{��rlJ,��Mgc��c
�Z�P�-��T����W2��5�rL�R� aD|�~��L��WO*�o=O���p�S���ݏޟU���F�\��,i2�d�t�d����C�ɝ�ﴻ���R-�SI��r�e�mB_0��b�2�"���C����#�Sb\�o�t�[�F�T���q������L+UU[פ�r����ѵJ�6��P�F�3�/=��a��3R?q��V-� ������D�J��:&sL'2ͧU.�P]��2�����l�1�T6��W��z���ޅ����P�-�*�VnB��2U��/jq�^ ���������n���~�I�H��\���X�}Yc4��u��/o����Y�"�:��R�(@�ޱB�.��~���n��qF����p>�_#��"F�O��9�4��J}H�,wc�%���(X�mhf�w���u,��@�;T��Q��LW�Hh߻t|Se�����\�A*�w�<���'d���ě�����-�߻V�!���<&�kW�Ǥ�Dc�˙�:������ 8�aP�;^1�s��=��6	�-ڙN�ў���.��4�@�󖩪şt� U�f�5����+���N���U�n�����\#�Y������a�����dP�n"��X̳��'\��E8�N���q� $u�fOj������)�>��)T8���9�w�H^Ua�D��jð�}���.��(���Ѻ5ֶ����b-����a���-慙����5����µ��Ǜn	�j\_EYy�G�/Ean����:�']q��A�`gg�;�R	V�zxj��y�e�����p�`�0�g��WJǳpo�j���2�hy2\���^�{kCe2��|�Of�n��P�p��0�������������e`���ݢ��?��r�4��K!M�Ɲ�?QV���@����^WV�t��0���@Qc���Y�]wg�� ���w;��tcy`1B�r2_F����K�G����Y��YP���a�CN.;]��C,�b�mq0�X��0�y�X�5���ܶɁ8�R�l�@����&^/�hi�{��/�H����+팲T�G�>6�\�C��LCH��FNf|m	��A�̇j�Yo��/���Õb��,��p��r��#����c
F'�۽A?L���nLS�/�Hm ff-����D�S#^1����'E/P7��+�1�ِ���3���.�)0�[D�X[�Uc�*
v{�J��G�uY�<��\	�g�2��[����I~3T ���D��E`�o��6��	�M}Œꬎ�)��\�4� �n�J�E��턣�Ҏo�t�oMi�]b���XHx2�p���xpz�]�M+3�^ؾm�d
������y�@X����<��n��4���F��?J|(D��|7�du"\4dq
L%�|��w��l`�כڅW)���x̂	?>F�q" �,�!��ʥg��&���Ô��[�� �Go�����Wl����!D�9)�Ϲ+���qn~�O�K�SyU�
AM���f�a�,e��Рa^j>N��2���ږfY
�,�;Tͅ�ENW����3�`V�F,��t_[���O�tt�x��uIOړJ���|�����瞥���M�j�H�n��;�l#{�Qе����6��am��9|���E�8䩥��Q'#J٬�)�˩dJb`ݫ�.����m��˔�Tv5�$�w9����ߋA�WY0�M1���	��O��(��7�WwvM���Ӿ�*�w��1D�H�?|�����n��.ۆ% �%6z���ˇSYĐ�������gd:������@��Ռ��+��k���5��
���9m�x2g���k����h��m�T�D�r�UY̋���R�2��K�\E�ӳ)�M�����^h�����꺜o�'��4#ߘ�����o�K<��_4�c�K-���7Թ�p-]��~�Ă��A�����	9��c������ɷS]�Z����cI��A�r)���k�*L'D�tb�1�|��w�Z���e#2�p�i��S�'�t� ���xp�d��$���>�wC�R^�O}�m`�A�w�CآP�@��}<o糏e�I�Ӣ|��6�͚9�c�Qc�T�f ������q�$$b:����d�=F6�60��MhJ������ǟ��/���H��a9���e���ODaa4{9颙p�|�%��(�1Jb]{X��e30\�_Q�`��4��^��ȾJ��i���,����UR�Wa`��^�3��5��j@�)�}���J)��o�N�H2w��6���4jJ�+�5��p�*R�KT �)��o��F���R�y�$wu��`n��6�P]�HK�Ʒ����6I�ӥ[��'y#$Ի�)2J��\_�����ɰ������ZMs�@��e�p�J9����ځV��=b��<v�>����s� L���\�	�.Au�S�Y���Z���԰MA;�2��h/�{|H�3KY˵+� �����/��W���z*EX�����$�O��z���g�m�
�J�<6�b�}�J'��R����pa�g�`�"�*���
���Z�E��,()a�0f|���"�>H׵p�g��c|��2W�ŘF�O�� �|s�*���.-����e�U:Y�ߧ��c	���`��^6�C�0Yf�y���*�b���sE.+�)v�ji5��OH��R�l�3�o�d�&:bL�9#(��aG�����1��,��*~;WH�l��� ��:� #������(�8�v��J,:�(-��`&�����qq(b��J,�Q�A�
L�ج�L�>33}/S�?"��o -n1�fTG�x�gUG�l��z�ԭQ�k�)�����Se��5�l*��÷����߲C��wFi\��X4T�<�\��Ͷ=�O}	 ����ld��t��5�4�Ci�X��#�J��Q����9_�t�P��0�@�#`;��.Q?^����Xs%�YUCk�5��X�O%�o;EG e��+�ɺ��HE��C���˅�ST����>US����f�����1�	k��頨&Eϼ:dqg���"�_ݨG�s����+��Sde�������,��7�&��\�V�a��{Kأ1�{���i�(��_z|���L=��4$���H�AVAB��ݩ��[� ���< �K��Q�G\~� ��d��i�|�V���`�_`>�\2(lڏ+:ǩR0��I�.Ö,#���.�|��n�՛�ɲ�A5��;OU�����9�h+���t6�sg�f�M��W@�L��Np#�������K�sW�&�*���E�5F*������(��.�P#�l������nh�/D^�
�?� ə�y�D�/�;
���[�N@�E2�c9m2�`�YS6y]���\��
���C/BW���m��e��g�����������!������uW�dd�6'�_�/��ſ���U������k����,�wy(�O�՗��:��g�gY��^Q�OVo 5yL;k�����]ʆ���m��g� �ɛ��
Z;�����@w�$������?����4bLF�1��� $�E"�
?'�Mr/��Jݯ.$c/�ߎ�?�1}u0��d�'�	'�d����}���'pՠ�X���g��W�ϓzE+����A��4��=EʋQ6@W�����-I�%R�2����	+��[�N>wG;nJ����H���%�;+��`I��5�-�c<������i��l�����shOB�ܚb��!	cFW�]�>�"h)�'i2i6��E���1 �Rpy.<r�yD`B�Ƃ!�2�]	-�T��cO�ذj�
X�2�|�)߸��S�#�P�:�����L��d8H �b�9����i[a�|g���^��G���YQqO�B�ԥ����LCfLx�H�s�g�ʁ@/��6�Ł�s����x�8<Ғx��?���0��|�o�@|}]o]a���yC��5"6���v�}C4�"��,��󥗠�����G7f�XV�����+�o���MN;�َ���8p��I�@�s$PB.\$����q�.:�Sg����D�����t'V���݊�2�jU��P�2�d�y��Kh�]�[a��:�a[v9�\�k����9�O0L��*Q*ނ��-Q83�#i8%��Ci��ܥڻ������/�Ô3ŵ�����U���\�5��78��O���*
����A)Q\e
�щ}7-��҇*ODC����f�J�0,�U�^�G6п��"0�CZ"Ed�˫�p��e��}�X���M�ඉeo��b/b�)~���^�*�����n"�ܵ��&S_��Rn'G���Zg�j�,��?�.��5�����}A�AF��j�4�$=�Ǎ3�f��=Բh�����!(Jޠ�[���d�����3�b�IC�J�ljL�@ ?�
��W�=q\Lv銀?�#�t�,m�$���Yјgg�i���O4M���G.��4����8��;�p�
�/�.�g����Q�<�-����0W�ײP\d��%n;AdNG�&�M�ޫ�\�Soi��3/��)U&�b��h��c��/�t�|�Cv�R�~��>/�Z�!w�|a�G>w%KX�b��%K�~A//d�.I��K��T[f�P���u��=���/9�biӔ���)r�r���&��5S��<�4+�s���b��3d�V�_��}W��E]Fm�$�^��`���'VX2c�����e}�*�4Z=3�노
��}����MCip5R���	��Yc�B9�n1��!��뭣�M���������Rq�c��W�;�|�?�1|�yD�n-4c��'�{^��#��C=ܽ�o��R @����e3nG�U{�U��+m�v��1�͵F��4�=�j��o����k|��P��Bzu�7��j�ח��B�~���������~h�����6�v����Ӕ��Z������ ��_Q�"��ʩZ��Xj��4:X�Ѡ�����3�$�h��3�D���VF��u�F��bNMz�2xv �����.2.]Au����<�P���.=Z�9$����H���4�O��@2=p�ً6#�9�<cD�*�չ1���U�@;ʨ+�C�y�:(>h/�'�`�~�I����K����{9K�����R�`�|���#&$�b��1�}���i�����HkU%n*^T3�$�d�hx?�M�2~ eiډa0^����ٔ�9W�#�s#n����$���G�����N�oM���9�[���!\���Y����N*�܏y��!~{�E���W֭�X��J0T��=ﷰ�ʕ�`����2�O�zF�Lͪ�0�������o]�*-RȤ�&ع-�F�W�5+���e������0�2�;Re?�eR&G�4����xV���#(>���Þ}�8�0�������P7i�rO��%e �J��z��)�G~���Xl�_��ȡY_�rK����5��0w�v��γߦ"�����ݑ)�Ш��_�z���Ҙ����� �%�t��KP?�А�}=�h��i����-͡���c�ׯjiHV�HUa��kǋF�+)�o�}ӝ'c�'6��8����Б$�6!�m/<���j�f4ל����H{�����I���-O�
k��WT<j�~�r��~�q�J���b�7f��ǵ쟄͔z�v}��C䀳i�d~�C����XH6����ݎGnD?��:1�ʹl������f.v9B�gD�p�
pMՖ�����"С���ۖ咁����"ۂJ=.��H�|�􌲄1V�~]B̾��謫���|e
������M^
:�� ���Y��܊���Z	�OH�7%�K���Y"ί�E�r�0�{':�O�Wղ�+�eͩ`�����9t8;!ƣ�Z�a0}A�2���EB�"���,�BJ�']��!�@X_!�����n"���ɬ��ۜ9A���zu���A"� �#&{���}�5ʡuUҶ�~G�'>��ţ>61qR�VCt'�-:�U�GiEl4�7��B�֊ٖ�V��9�3��������ԛ�Qq���d�V ��){���V]�Fh6�@�B���Ý�}�0&g�O 1�8ӥ'�nƷ�.9��C��n#03��0��}�6�����"�ϕ�ݯ��_����p?� (;�c�B+:�)�MؿyT-!�� ��}k�&��vi��ŷ����`�x�J���qP,3Ս�
�%c��7�?0����7�t�U�9���#1�[�_H��#Q�LO\7Ɠ��9�=C�Q�����c�/}��CF*�#���>8\m�W�ʀ���)�F���Q�T��g���{49��2���wN�{�q;'�yg�g��l#N���i�Tt��<�𪋶�	���Y�)�s�'����<Ӆ� F��OR;@��n���fO�ڛv��þLB�!�]Ѵh,2��`�pjm���;}T �]��ϒó�O5<$:	��MfRd��8]�}:_6��iO�������@��\3&��'��N��M'z���n�j�r�՞7�yM��T%,� �C��|��c���af ���7a�N�I�Cn�#{�J7,���(��5�:4�6�-�δ�0d%���7#��v���s?���(���mvv��7�oY��C�%l� ��АӢ��3_�q(�<��
@���i#ߝn���R�L���޼�2�L9b�������o�U��ݣ��n]���|p��lM-�J��4�p��3Ѭ��JG�hK��z��U=�<5���G�>�xrq�V��:����|�X�l��zK{?�G޼��Ȍl�>J�C��3O�5F{�m�d�Oq8� y�l{bZew^�t���ʼ4ƈ|�lxV8:��L��;�Z�oUi	H����L�?t��$y!�.q����.�>�^so3�j��&u NM��k���$�?g(�\��j��d�[3`���$��O�4I]vE[�y�+&�R;)5� 7�<���j.�%�о�"o��(�07AK.����@*�����z��=6��uL ���@'/�����'2'�����U>���y�oOx��{}k���נL�M��D�*E4���o�!�Iࡉ�d1���d��b�h=^ٖ�#�|�p_�۩�b%|�a���<ȘEv~�G��?����C�
�z�i�QM�\����n�����c����줅9����2�)�R�)�x���A����_�k�Z#�+GY�c����o��t�G�C�5��m��T� �4��C͐��J(@e/ @v�Ix���䰱J����ۦ�	+�H�T]b�3��Z�rF���`Ϩ<�S��a>i`�Bm\O�Gu �47��������a���'�>��[$��X?�נ�5�o�E�Vs%�c���y]7XQ���3�h�M��4��G�فz8=�eݔh�𤗍��6-�7��X��ɂ����X]��B�;)m�i��m�3E{+�(K�
I�a�s��y��_���j8v���za�8c�9��n����%��w�m,"�A��@� <�H;�` LR��� ��Ƨmr�PDo����ڡJ� �ϕ ?�ֵ�+�z@�=��jo��ֶ.�x�`�5��4���?C8�P,[ Q(��E�gh�Ѐ8$�A�يS/�5"�#�S�H�+��2%}�ݑ�xl��[oj��T9�
�u�ʦ.�;��>�O?HA,{�F�
��N��ڝ�!nU^,����`���逇��(�w��]CI&�_���~b\�mv���ݠj �,A�X	��Y�a�ҏ�0��ASx�ؚ��tã��3N�`��ϤV��ͰU�#�0^0��"<�)����-���+0a�Ni*�=��=+���w�T86e��g�� «P~�����a����Y�-rr��|��,�!14iSٶ��Ȁ*㧤4�@qnA艴	��D��"�Z�Qku�"@P�XJ_��9TN���{�ˊ��a�
tL�5���XF�r����#�)K�K{u�d`���q�5#C�R:��4)�ix���I̲��k��|�G-���p��R P>����*���jK�Ȉ~�5�I'�H/���Y�Bl��