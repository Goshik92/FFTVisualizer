��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��XMXl�M�x��ֈ�$��/Fק�t'��ĩn���}��_�]S��W'����Ēʅ�1ëN�S�]A.���^�&����N�!Ci�6�E�.�(�����)"�?7R�.�l؊�|)��ѵ>�/V����r5m��Tt�&r�0M��T�����L�ތ����vg�P|�[������6�1��zjqj�I�CO��ĝ�U|%8�FZ߾c�s�� '�����]��r��#9"���;\!���)����У[X�������MUB���!��׻��ZJ���xЛ��$��������
:��Љ�):��%����$��T^{��KD���7P�g���U�UsOX΋z�
��7�����1�v}sj!`w�ʊv*�k�	�]~�d���ר�f�7�d}D�V�]��L�-�s�R�
��v]��e�L�N>�6	���	sj�%�/~�KX�xay;O�ڤ0�7l{�d0bKh1<��A3��z*��olvi���\�Xۓ��zrJlL?�1B�Ns#�$�nC����1'�����w����Q�ąf�á�J��*���5������ H���ĔJ������՛z����\������/vy�  ��Qy�P�$D"a�B������#3�@s<CxM��v��{��|ȳ�>`D���#Ј��9�[r(u_$]���=��C�Я~��|
z\(�	Z([���g�$�ɦ�1�h�2 y��+�Q�s=��*�����F|��x_p9☇+t<H�٢f3�4���,zD�Ѷ�R���+���|�g�u�Il�ئ��-���ԝ#�ϾQz~�L�;z##�m(�Y�j�R�[Dc��/���\踃N�ɿ�l����3!�e���ߡZ\��$�lB����\6�+���î��x�݋��i?&���y&�Kr��SA���T7I�_��� .ѩ?Qo�"G�d�����{�7�ێ _�+WJA�g.�*���C����^7���6�g|͍+F���e�M��Ô���C���ؠq96�]����@�3�c�7t?'��撟�L����\���1i��.M��MKbPc�@+tS���'�?�l�tܱ5DA>�1MP�*d})�ef�)�ZhF��$�����h�������8�.���3��AjK]����Al�vy�*~]���u[��?�X$���<\��6�} ���Q���F�wO�sY<�n��t=����/��V	���dД��u�$
�v+���a��^YS�f��������b�a!pOBг�^�,�Ɗ�/3�(>����	I��LJ5M7�����i�[�6�-X](v�T�;`�<E:6���d~cn����D���h��X9�O'�8G�秨D[M�<���W�i�%F0҄���hL@�������V���k����9"�s�R����OV�:��y>v�yY9P!�}b�� �F	��6�~�;	p�R��:}��`�6�n�W��ŉ뇱�p�D�q��<x��U�"�i�>�����!r�;�#䕵j��g�П�<,�"��jz�AN��Б���qFV"��-(h�-������K�-�9��d_[��j/��ʉ�+� ��Xc7v�SX�x�����?�;M���ߊI�ҳ�U�
g �3�%6}�ч-�̀���J؎'���~��|�_�Y�
gɧ��W��vh`�UÚz&9#�p�9��m1l��[��ڧ���c��Hq��������Ȩ'#d�Г��3�O`@S-$��vGȋ�q?3�^��g �0wrv��+�>J*��K�a���"��˒m>�Ծ�����N��k�E ��s��k��H���O:Fv���'�٩�-򡣣:���]���O��$�����o�A5�?"OhE/�o���!���u7q�ɟ���l��#0<'AV�o���VM)��)"��u�ŏ������T *wc�MU�	;�R��	!k��	�V3'�T��/�ﰅǵ<���1�>@�J���3i?�V�Ƒ�d.��"����\���i���ϑ�7�{e��Gn����Q]h�r`�yE;،ְ��8���l��h^+�<gT�8\��_��Ԃ���'�gC�� ���;C���G�Aۣ���5va�J�1,�2�˄�w���N&e�î��\�˜VU!��rn8�KUi~|+��6n�e����9�eA�0������f?�=����7s�d��#,�����4X��v���A)1EKC ����'�N�$���MҾ�����j�;��7qc9�J���}����@�R52M����۪N�}b?��,�>Xz��Ljj���G��ݸ'�tΌ�1Z��՘:~���n�yU�S�!�CS7?�Z��Z��r%#�}l�������=��e�?� ��G���s��t�RO�*aB4�\H����Ѥﶎ!ێ�p.�=(�M`&�{2��/�,�(���������O���P��-D��R1qSj�/C ?����4� ɮ�\�?��D�P~vN;�zb�)�Q�����@н����TM �O�n��I�S��r4�Ũ����[�2ۃ�9a.��f�� ���{.�Ge|����Fvh��Fs�c���l<�;�<�����k֐�>��=�U���s:#\�2�����1�����r�r�ؤ�_���^�[w�>�� �2�j����%�Ɖ�:���^q4>gH-|�35�Փ_�R�@�V�RI� IYCV�=��_�y���|/P6���8t^黾%��-��luoz�92�.����m(�3�?�n˯X`	�D������<������	O}xA�!�3_1���%{��QFhv6'f�t�������X���A��h���! �$���t��VoL�
G�h�r� ��N08��Ӣ�t��^���B��F�R�Ͽ��$��]ب'�c��6_防�APB%��sZ�Y��	���Fk���QP�ȃ��h�ȋ��esQ.�����%� ��������*ټ\���go]�5\�!51������*��~cᘪ	��)Ց�W�
�ٺ��&T2��֍INs�eN{P�l�COY��y�/̻	1�f8)���Z>x�@������
�Y�P��|����R�]�U����5?�N��>��`�1+~�F�*��-I�4��*M)`lߠD�0�C̉y��Q�mGiЅ2�dWH�N���6��k	G_#*4o�y�!ǴI����mQ&�(/{6k�-b�&T���J�Sڌ��]����Q�G*)�ǩ�K�h�0�#����"I�V:`Q7"�(�Nr�p�%kEF�{o}�-��/����-q��l�H�|
+g�#sb�s5�hzA?'�p����ݷ��4^LЁj�d���M��f;;�����(����81R{����m�P��"w]ݷv���Т�ǥX[�]I�1`�Q�Oa��5Z.`�R.y�-��u?�ӣb�����A�������i��H1e�88P=��+�r�'Խ�XD�l	
W�^:*�a��P���� ̧Ȁ׍���T�3���>��ҠQ���z�&v2\E�Ej4��A�찝��e�w펂�J��T>��,qZ��A鑐*��5(�m�c�^[HTO�ٖ�G~�-g��PgޝH��M(�*.��Ű�	��"-X]#��1/�Ԡ����g$��(,���*�x0f��4W�ܒ���x��Iuѷ�JR�{�SvZ��_���pݐK��u�;M�lhN����i{l���H������������`(\�?�#\Zy,:`"R���	�v�r��=�����ߧaw��+K��}�;�g�Z���K�.+9�y�2�'m��Uu��c�v -���� f�>�n���cbڡiM�vkQg��t$M����$FvmL.��Ql�2�hzQ��X�mT�;����Q;1��բhESXҟ9��l�(FN>���%)���r>���,�c��@\X���A�]�����/�[�	�4�4�
��X٧HƃW�j�ac9Ѐ
E:��Lg�V�s�"H"��du���lh>��I�|�1�g�E��/������oQ�b��t%���ϰ��6JW��#���|"�������V#�rTD�������V�3V`��Y�K2�}���p�ĺ�D_D���k��R����?�ϊ���,bD�圢��-�8����-�0�ꑔQ ��{��.��-m��=���b\�BM��H:B�&���f�^s��/\VWT���Zzj@���;�{�.��B��M�q��R�.���@��eٸE'�Q&9�_��A\�G^��
TH�q���wq�8{��]!9-�:�K:��d?��+	wctJ�G�,���q4�B���B�]s.�����ԙ�<�/J/]xP�WNlb���$(eV?��u
�'5�&`�7H>J{8&��f80�����Æ��:V�V��B��ʄ�ك�܉m;=�����+�ɡ�d�+O*9��k�1�0o��+6 �BO�;��I�nKQ]6����I���$�ucҙ��F���u�8�Z�=Mn�i����A�w8_@	^���p#:� 9��H�oh��<Y -?	i��H�ď=�s�{�껅�t���@���_K҇m��Dt�9�c�!
�����$'��M��"UFV���Տ�����(�W��5�-N:�5qS�����3.9��o��B����R	P�Z�q>X�t�7-�&��T�T�Q���<