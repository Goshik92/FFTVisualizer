��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|����z=+���v������� ���6�\?���������b��q]�rf��<Q fUk�â����2Z��)����UU�1��� :�^8�U�	�|�E�$��s�&5�?��w�2r��K��\�m:7��6b�r2��y�g�T��C�(����g\�"��z ���j��Q���Fѭ \S�r�(�3>C�-��bu#y���Kc����m�<��c�Uk�2�0�՞7~鳎�g���!��؍��@Ҝ�K����2בڹ�$�dI
먘���|�<��T6ʿ���|w���W�ߧ����c�������/+
b��Q���]0��$-w�S��!�R��4ɣ����"�\I`�F���nq4)Q���G��rZ%֠d�:�����sfeY�a�i���[�>%�61�-|�d���e�h�CM�S5A�lY�.��.�)�t��ڶ|�q��#��J�j�)�|�o�i?��eT������a��4@�:�r��gM�}b��ݾ��-�=�R���.򳉨������P���oU�3�h�A�.����3-�x��M~�Y���x�r��5P"ק�*���$b���!�'���n�5ܪ8N����Y�cd�ۣ��2%v���ޠ-�c�'מǞ�����a��N ����r��Q�{��b�=�,�独�?�p䄲�<�N�����<�G]Ιw
ܘ�|�"xQ�ZD�ɛ=A�BC �#�����ZB3�'��_���h��|�2u�6g�P5�VM1]����}~u���3��$�i�?.�7�:Q�]I�K��Yb}��vd<+��$�w`}�ԁt]~�R �K��e����:?W^����J#�/L�?��5a<"^�(~;�s8���]:�:|�~7�h���CW�󸄑����sh\輅am����d!��!���E(�"�~�R
��3Mņi��"L�y����'��5vbi��}vD���/*��|~ �8/��49r>�MQW���`)����6\�4��baЏ{)C�y�φ2q�1�f2bH�������E����'w����x�q�kbE���%�
��WS��~�3`4���gG�@(������a���e4 `⃻I޽;܆��ϒr/�\�o\b��u��@i��7>����
�[�ؽ�c����7�L/no�)�+���3%n������q�艛���U�T� ���]�A�� �ę�sfz�!߿��o�9�w&6���U�;��r*��d]Z��5bk��Q)��.Sb�L��{��r���,I���w�t.PZWi1Û�f�owY���J�6 ��3P�d^�Ӄ���N?O���Ne��:�*�pdѺ+Y�L/��G�4���Ͱ������t���P�t���Ή.Ɖ#�Z������jk��s�V)ƾPE7�cR�4��~qD�3�e'W���*�L^ۖ����O����ۤ�������3fjΙR���[3�|�e�{!;~�fF������'���6 hCWډ@Ҝ��FY7I�3F5��.����g�^Ը�>l�aF�}����@���m���ҦN��f�=l��8L��a*74b*�O���b[�.x��@#1ͤ��V�i`9�[�ݱ�}�HJ���e!�u�T~w5�5�zL����Q�S�	y�FH#d-K��{p���qv���o_��<��@9�1�02�GN��r�w�o�e�f���h�� �@?���4�
�D{Jm�Wc"���]�M?�$(\$���vi$��F�Wd��m�O������I��F�B4����������:���.&��E~�Rڠ�n���6�`\e�6��z{!���[K>ـ=/d��y�)�a����S�wՔ
���ok;1�+�AC�(M�_$j����PS��CJ2b
��{���H))ڌI1J�a ���;���:�v"��_;��k�v�-Z�,�>B�|g��b��_���;)h#��I��uX��!�>}�'ەN�N/��.~��)�j�F���M|��t��G�c�
�����l�;7���Ƀ�e݉�mD�s�w�MF��o�o��s��1�K|F�b�ӧ���a{�'}���p�pb.�d7��g��X_5GVgM�-PC����󒈮�v��0��7'�� 9�*x�w�#���C��U�Ze�-�	�L8�3B�,�E��,��q�Ҏ�P�ͤ��<�^m����2Z~^$�0K���C���R�#���*%�Jpp�T~f�?��O�%��߿�?�U,�n֨u=*R���;PT�)��IL�+0�A�Fj�뗇 v�mY�� 0b��f-�L�
Pzw"��l����q�~���bUyJ�]�$p��C�RЂ��$C��F�Mf`���t9�z��p�A��u0܂dH�t���m�x�A�rhΜ�-s�@�1�a?G�@m��*N����d"��@qތ�U�����qwӆ<���`�k��U|�	tg��[*G*K�)���������_RP-�:���ؼ^�d��e���0���	ƆR��Q�B�;�5�-�:];�CQ��x�/�u�NS�B�ʅ�1��j�Z+L��{�<��˕��:�?}8�z��L�F�тk��J��O]���$@��� ��G{c�	�/
;M� Ez��m>$�8�<m^3�=T&G�����{^.��h�!��Z}Q�H�<��eH�$��������V����۲!ߊ������
I�[�-|��8���8zm$|��7���Ze;�����e���h�ΝO����z��`���"���J��[N$MI�Os�GL	�����uť�?���z���R頨��x���~~`�(����K^*+��F�zɽM��5+HԘ(����nI~*!��M�>�u�UM �`�j^M�׵��"Z5����:�
��?~��g�w$9�m�x/�`؃�D^�4BS�%$���L��r �B�`j�$J�O�Xnvj����W�@��bP�/�y��k7K�9j���B+^�r���Q�	�A�����u���0�O��Jz�����[he�{���RLӔ�1�7�1 :��Xy1��d�fc�$�~B>Fӊ��h�TC1U����+a��1h����X�c�:Ҵ��;�u ئ��iuO������� c�e���^�1�zGBui4 �gܤד�����S��d:ޣ�� q����P��.���H�B֜�PiƦ�Y�e"oД%d�d�\&~�hMYTD�je<�� ���@��3��1�W�fp��<)�C��{�`��G��0xe���9Z�_�_p���%�?�a^�7G��Oݣm�_0�e��TKӮ-5�Qh�+8ݳ�4��l�9�ϣK�v`�L@�6�	U'2}wM9I�X�Ł�1��� �~�T�^�ۖo��9��je�d?p��HJw�e���s{���y��%B��;=�^�ZW����iE3�����v0�)kl4�u1�q���bI�?T=}t��C�C5M���`���(�n�=�@L���6�%R��ꥻ����-��иF�<�9,cN�q�I��:�R��#��Y�-�(�������X� �%"Yn�"<9�q4�ˋ�0���O���0i�{=3e�m;�דh��2���Q i���꜋�s�X���