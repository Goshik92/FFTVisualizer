��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y��yO(e,��.��̡�+P�FuX��d-��N��$%�I߽7>wN����u�]��j��ܹ�Ucל�|�=í[~��k�5�P�ؐ��T�5�����#�p"&�l�z�Fr&b6��,���Fԟ�Z�_�X�;���93	�����Ǘ�M�~���٘�2�c�D��������f� 3łߥ:ա�;kv��ތ(�}��r�{|�Z�LP�����!�Y{������I��܊7Է^f�L5�:�	�͎������W&��b��wD���Jݎ�IK��et��1���Lt�:��6�Ui�;F�o��!b��\#�Z��k!�Y�#Ao��U.H����Ƈ'U������0JN�]�[�萙��5��!M��	��1چV�)�MM�.$�uR���4��m ��Db��8��"�H8j:j��K��C!�Pv���l'��S@���Ӽ�!�X����W�2`F�.��֜�S>�p^�`���U��(��ٺ�+��KIZ����s4`d�F��(�dźM������-�O���+�ra>^��~��y�#)T��Ɔ�K\U��_nmx�)08��V�����$���F� �����M'K�6	�cU�JѮw���n'P�ɩ�������4ԩ`G�@�Ɏl}F��>�X�8�F�Rb|��L�����1# ��"I�ʶg���z1*�
_:>�;V��=Lӏ��-��΁+�Z�Xo�MZ(��be��W���s����d�-�O����5��ӥ�%�W���bh�zcb�	�N�t�����-�:�.��w�b���K��_q�f:�f����2����\���a�jU����	�t����e�1������B��%hޝm�XK���MH_�/v��<fx!�K ��B�)��-�G�V���T�XU����B��� W3F"��a7�w.��N�"8"3�K{$��pvB��gT7/87���	ns�&�!Ǡ�x�H�|]��U�*F(�
v"�]�]V��S[��?IϿ��v���kK�Lۀ��g9[�j�D�W�舠-V�/�:����dF�`9`��/�V=��~����A��Z�7@��	�3I=�@��j�����bL��'��+H�^���O�G��T�z��d�m���֎��i'���:Q
J�"ɻG�(�������ɍ���4��v�;�˘�D�I�^C-�hO��'����_��N���3��m.N���x@X���l1�< V���iJ�ނ�(հp��e�Z�K�z㵄j�E��P �oVUa���B�XQD�QT�i��Aa����U�w����cρS��܏%��G�9>�pi���l�1�N��![��V�%��� �xD�l)e:�����.Gګ'��9��l%~��
.ŃP�^nl7��M��ƅH�KN���c���j��P+�\�P���N֭/��3�f�vb~�����I~�\3�1~q��}
���q����Tc�ö�TyRJr|�F��/�	���-���M��살��N��h���z�6ncĥ���2�\�w�N�-�
��j�u!]�v�cx+G��+x9j����?b�W�2E��p"e6�:<ݨ��O�#=��pRU�ѣH �z-ru�����D��]�>Y���L�|����R%K����X	�W�v �K�/�O1��T���Z�����s��<�h���>@�������|ޔ[�1�\��[����d�bS��5�����D_ԉ�=.��Ň�'�X{s,����mc?��t�8�"�`�G��6���[ M@���U?��Ir���]\����-�O�X¶R��b�A[�k���{L�����/� C�M�	�8�Q�����;�X��<�ꕄ���{l�_�p-L[4㞢��w3P���lt����2��/�
JB�?9��$�<���?
���6�䎃��a���f��:�!��������]�;�� 2߄V0��_�Wݦj�d��fI�-5�6l��S�:�-�o�dvY�M��.@(��j&�^���f�AG#���3�6΂�0x�e��r	�vW�M�� |ٱ�OnQ ��6�7B�zǗ��W�P�	������~�Q���l��Xh��1Zvd��K�8fr�J�a�p��Xb��TrQ�&�˃3s&XT�C��9d��S�^�qx���A@������ ^c}N֥T̲wsX*�Y��<�ǳ�.��2���JP���A�Qh�>Ϧ�u�� Z��Ο}[�P��K�{�i�*x�,���M��j�����w���y_�Q��9�-��՗}�Nu���u�X�<.\��9����>��ai�J4Dq_g��N��
x�6W���\���]S�!���G���1X�P'��%N�92<�&TB�6�u�x+���+sc1~50c[ ��l�v� p���K����|]g��F��5���
�ļ�·���J��b��9����|l-�Ӈ��[Z|�K��.�[����\3�~c�o�r�EX�t�