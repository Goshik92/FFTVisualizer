��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|/K�^!�� �Ϊ�I.F3�h�]D���� �1x�ϓ�k�K]b�ec���9�̑�2�۰�}EW��E�aǧ�b��S��+�/Aė �d��׫�~^^��y�4�4pjTK��~<OS[�EI|�ݾ�wi���tW3|��.�O�AC�Dl�w��;�|�y:�	��gL�0���\X��D�0c�8�p��!Z
�O�.s�H��/�hȍ�`���@UR- �BϤ�YgP�C���/7|��
���EM����\�Ұʝ@g����JDyܳ�b���bH�7a�ȳB*��S�!0�PDk�|�U�S��D:�Gl�p��q��لe㷗"�Cfe��b�ߺᏻ\5�2wϺĒ��S�;~��ж�Uwr�ޫ	,S�'>�q�Q�T˞+�A'^Baf�AC�1��~*��W23�B!�->n��$�-;�])x�Qḡ#ۂv�֌��䱥��o��n�^�_YzG�1' h6���Z{L~&��<���E���h��Ә�7���&��qKܖAK�����] �� &͢$m`�&[(7d��2ȁ.�i��h�Μ�r��n�2Q�*��W7{��{��-�	VT�׹m�א@�e��H�;1uW8�|�X�"�l�[�����$�c�@���-Q�}񆖕�k78���^@���F��B4�q�(�o��� �!���,@-r������Fa#L��dO����`.v�ћ�2��s��*�Ћ����9�-]+}8=��
4"�8P��<�1"t/Hxץ�}a��`�ª�&�y܇f~��z���Hԡ6���Њ�1��K���/�Ң����Y��@$�����T�*�x��^��jܐ�$������=�U� #�(�oS��?�������ڑ[i(q �.Ai�o���.�ܜ��n�@�]�+�i���+D���TU�ܰa��;=O��+U�h����&5K���������K+FQ� N�T~ϭ�Rj�_J�zfjm��X�����}�����i��!E{1-ߟ�t4�0����JJ�Y�۫�2"��]��q�b�lZ�w�q�lF .�[���H��ZFr�=�p{���k�	�7�� ��%B��'�ȝSGff�Ta
�Z��8+3+ʃ����>3���>S�� ���0�������
���u\��P�%��=�1��J�A�C��}�Z����(�{�'|�� ���:�ꂝ]s�c�:�6���A,4m�	tD�y�GOO�h��w����t�����#�	�?�a>����q�~'�*H3'��4"Y��'A�p��`���8���9h�z�������O�:u�$�(hڹ��8\���\f����&���:����A���<�^ybF@�!rRw�J<1(��n��`�
�k�y��V:�10������pE:܅��]mr^J,d��<�9�3�эtJ�+=j<'�.�������4��֤�?;��VZT�$\�i�n�̜ʵ`�)v8�Ih���^7��w��"�b;r<��#�d�Z:� :�=p�b��	�\��	AV@�2�.��BT֝)�Jm�9��k�y79����{�k�S�_���و(�	�Ry6��P򪢕bB�jJ�Hg]������ݯV�w���Ѫm`��Z�� �fa4�H�ؾ��ɬ�~�!��`����7Q������[2��{�p�X����@G�͸�]��g��GQU9�|�+�
Ǌc9���m]�V_�u2�Wi�r�6��ĬW��{vZ� eO����6��r!�fy��X��v��� B�i�_]�L`���ce1�ϭ��k�7��k�R��𺳷`�7{Ǹ6[=���՜�mu�Q��7��,�:Lvm�P�^.�LL�����[@��")��d�C�ph��������yY��-�+TPf�W�Qv�ߚ��$5z�)9Y@0�� ��0}4�� d��L����5>��jk�/�ʴ�Wx���6b��{�4sę�$����fS��3�/���vA'H��w�q��Ǭ��0���4�Z �(9p���#��;������o�a�t>���-�MJ��x%U���!pU�iݤ�rf'��,��÷Ae���k_�jk�g�8}>���q�1a��0>���ψQ�^\���s^�v^��7����gV]aR�Ѻ[$��Y=OG��/�`�E������$�c�D!׉����*T�)���n��-+�q�d�-�7���ȩ�I4 �-\�s�l�꒗��_;��	����:�����- ʐœ{�HX�4Ɓp��yh�E�FcĮ*uu�!]�Y:
���FTS��|T�_aM1 #��'�T��3^��4�|F����&{� 众�RM�NLu���"�:*� �Y��g�*ȿ5L���S��Lf��A�v�v3GB9�������sd4E�uMg���r��DU�|I��������LQ���sĘ�ke�;T!��
���캓�q-#p��cj�ϱ6��Oʡ���UW��\@i�ƿ��� �hŌ&ՠN�ļx +����E�����c)����HÊ<_��\���Pq��$��V�O$�$3:mۀ=�|G Μ�s�Ԩ�B��5���5�7��5� ���#��1�~5~�`�Y�?��@��
d����w�AXj��Nl�qٞ�������J�
@�Kg%���,h�����NZ$�6�_'�8�l�d+)|���WO$$�d�<���a���)olb��ed�@{��	g�f��:�B�ֻ���X�ޝFp�*��w�G�fC�}��!K��2N
��9�Ȣ���V����s7\I���sAqF
�跛$�V~C��T�6����mm������HM˰y�,���}8CS�����R�0��{��{k� ��-\_�K4�p�GQ�$f���I`��/d'�! *�*F�u	�Z󉐬�gC�Z+�2�?�|�g8��QM�l2�:̊q4�W
Н�,���F�5���PMK�^��xpI�e�5��=/%����'�,k��TQ
K�����ǓOAػ�FX��H�G:�r��tcI+fW�P�i�
0@j�m���I�i`��R;���S�{�isּ�Fa���;<�Ι3��"8�*����IEƵ�P����F�t�:ფ&�\�����xΕ��g0>RFx�-�Xj-�"|��ݯ�1@���D�X|-w�[�&~a�Eu|z����2��e��ɤ�0��D�3Uh��J9B�*E3�����)�7��C��h�Y,k!�ѱ���R>+�D�`���>�ݛ`�L��������O`{Iv�̠�O�2@xI�;De��9��g�������ޠ���ad�K�^L�0C�aS77��d���<���ws�&�Hӱt�R���h��Vj`\.�C��J�q$Mqɸ	��G0B(����ޜ�' ���ī����*��|���@?�`�'�cT�N���X_k��V/�%�`,TkJ�Ɗ���N*��ɋ�QM���� Q���\*c\Mu1j��G8�?�x\T�NK�}��Y%9H�b{]�F��$6Z Ӽ�	�|?c'��*��l%r�� �.TL~���Q��[7��3�V�T�$����
�ȟcu!�?�ԏ�7�W��B$z�^�p�4������u�:��dF�%{�;f�e�~��ƽ|t�Ϲ޸>��.1�J�|��L���IKQ@��r��ޒ���{[j��fl�m�f�;z��k�,��Ib�3�Pd��H0L�f|ƀF��dXQԖ/L��L;a�������g�-��k���
�̱C�.ocZ`}�Z�W_�F�G���f�����:܎���B�(��l��u�uL]h/���C�Dp� �=#�&�C��ԲM44G?���*�[��ѣ���K�E{���H��vBx7�T�D��'%�QIa$,K��LC��7
9꜇DΑY��T�>�^�N^!�%1#_����W�8�D#ޣ	�t�&ٸ��=g�fj��LE٣tu��*��$:�B%����y�0u��(����FdKcP�i�=�����}�ά�+%�1Q����������~�>$��y��]Ǹ�:��Nƅ�j1���1�I�|��/l9߯��dm��O���`ӆ� �'g�|�d���fC�]�
rS �sի]�0�%���F��J8x��)��IE]���yA�D�J/�։�5M=�����]Q��l+x�Z
�-1H����4O�@�̱��)�n��y��RH3}@A���M�m*lpmx(/���ml��KM�i �`�̀�}�B���Y)�Nڪ��,9�U���h�!.���ɇ�W�����F��v��Ғ���$P�NlE����b�V�d��Y�=�"� �ts��D�a�&��z��[��5�����p��?������TVTK��m�]�Yɐۧ6��h�5�$��z��bF0(�I*��w.
#Jhw�^sP�cD���봑���VЄ闸-}�'�Db��0�(秏II�φԘ;��%܂�	A��;ʏ�Ek�U�tC�KT�A��rN�(�J��ͻ����c�֐�ɦa����]�*���Afc�������x���N�Z�W�qh�L'x����#z�9���:�j%�SE>��d�$d�K�Yy��D��r\X��dYDuq4��g�&$ʮ¬.d���[����v{xq��Ǳ`4:�
y6�8��`%u����A�ފ7���ך�H�f5:1��kd..9W7r����D|�,��TE}H�9e"� !������M��F��*n���B�Y��`���5@&?��ꡑ�,;uG�"��4�I��%(B��8u�2iB��|˛9�;t~⍢[�Ե=��f1j���y��嫂״b0�b�����{��%��Z���ME
	���l�@:����XU#7�^�&���~K�)y"E�ӺOM���{H�T]QT %x�O��1�a��J����[r��0�'����/�q�y�3��⇐A�t4�o樬�W��Yhg�l�e�l��$wǮ,���U��Y=�es�f���d��s>\��{�?��o�;@��m3���/n��Ɇq�*���������fYVK�s\�ڱ�v G��Ǟ��&���s�^g9��Þ�vL1a��>v*Ȱ�SN\b>6�!�`������.���MO�P�z�Cݚ>ޛ�z��Y���Lde#��N��M�^�#t:( �)�	̩�_��l�bP�֟zV@�641e!�<mq�r��oS�I)��`���A�f7%��oI���\�R�I��!5gB������9?�	�"��V���8�wŒ�V0�s�`���ȽuL6̊���QC�\	�y�ق�#"���hk�~��՘@�lVz�Y�MG�; 0���'��'���G9�*J2��IVJ�ڀ��rv��- ��!S�fI���S}�3S��_g�]���*a��\�x9�E.@�?�����J}��N�owf�Y'�3v<��6wz仏�F7�D��[����Tԣ��S�����a�E�ϲ������;��b�@�x?�\���2	�]�x��������Ȭd�4����d0�G�)�i����3�b�BL��˺�ܼ�H��:��>f��+p8\ǥu��?_RɃbM��T��+C�/6[�+���V�cec��7�l�,'�c�6F����y�6
�X��ED������uiQ֓��m'[g��/3�;"���5�v�[3�+p8p~Lۢ��,<V��ݓF"]���%��റ��	a�ѿV�&��d$l+䪇I��9�@v�+)IQ��>��1cϑ�˗��'�T� ���bz�6�?�� j� ǜ�H�[�.xA6����Y�?'N����K-?#�����ʲ�߰�9!U�nܨb	 ׻�%'m&5�%�g�*L�2+�O)�C��4����̠]UMw��-�:���o ����ɳ8��؍a���s���C#o4z^�~�x���U��)!���N�)�{S�JP�U�y��\��m΢�+����2�|����=~�l��`o�1�l#R��Y�'І��b��d̣r���~�K[Ll�<+�����9��W���M�g�oؑP<��a�AY�J�"?��(�֢Ϲ7�4����Wv+bB�q����'z�OL��["�Μ8���7ed�78�F��Hr�B�*�O��޽%?K[�Q�]��Rȕ⮂�b�BH_]�R;��8��������i>���F��zI���"�#��,�(�Cj@a_%&b��!���'�VW�s�Ϣ�c��� ���]�6��G�C&��|�׏ﺉ���
����,!��)�/��,_.��k8n�ž�c'�!�5ǭV�A�x��~*}�Im)rO�(%oIA�TOݱ
�͐�<,�Ŀz��rǆ�T~�au��)3"�^Qw�1㏥�W'j͇1!7+v(7����/-AT�<yR����{YU�K4m��"Q�����f�>1O�ȳ��+���W��%s����z�bo�զ��>�����ԉ 
 Q�{��yk�#��Bb{��F�QP YTw�EO�?�0��(�g�t9v:"ץ��q]܊��,�����ۮ����b���Y����-M3[,�� �}���9G"zTsӳT%W�M�c�Q�i�+V�H�:dِy9d��}g����>L�V߬}b%?�X
-r��s����7����X�>3�ȣ(bs%_1� ��E鍑�?iߍ��yc��z�W�� dE_�%�^��9��(�9��'�s/v&����������. 06�����\�L�A=A���)�bj���^:��%�ǀ󶟚�L�~C���6�'4�9��RcI�%Κ��K�y�F����Խ!�Si������#n}����	��ơ��)Tp�d �/ɿ)s[��K+D��-���q���{dX!��);�@��v�m�FQ��ۉ�C�Ǖ��Y�����ꚃsY��6K��)G��vc��<v�)O10�.�b׷/}�c>L�n�xr���?W�9�S���rL�F�կ+� �/�L���u��N��֟I��u�X�b��P�\ԙᛒ�;"���?3��8?ĉ�5&��p>6J�i�B��j=6|��	�[ظ���-�.�^��_7P-{���d�_t�C�{8�;����ٸ7&����m),נw��o���ln$y��ʶ�6�BtZvq�ŗ�8�l�ٞՖY��f�=��� ��C ��&�5�?�vv���u�Um�RS�R��ȝ_��%�/���d�ꩁv��j,�;�L�yfEd2�#����ĥ�>�X*��N�x���q�9��埯��b��>�"ܒ�Q4��~Lk�͔��O�n$%����dJB�IH�P�]op�J�zR6���:�W|��r��&Wz�*��)�:�)�