��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|݅o�@
�nI�֛TU�PP.�����+���u�Jf]�ϫ(#��$�r�jO!�Q%y����m����T}�R4�?/䃭0����AU�(�ƾe��������f�7�m��v����of� 6�{�
N�m�H2
��j�Y�?	l�Aō4�8�����>|�f[؁���
Ζ{�����0>��������'l�d�b�%#T���QOo�Rh��&42`�-�R3Ml]�Gq�]O��ל��J���('���Q�5�.����p��� 6�	J�/FM��8���b�)f�ĐI];�^�EL���j�����D�1�5�1�K%M6P�]���*"&	а��u��~ٷn$5h����k��O��L���׎D�y6"�  UD㍺���"O��ܣ2^ �4"�.��d_y&����V���k���ƭo����`���%ȯ��e��εA;�3Yй3V��l%U}��N��������aUiJ��������X(7:�_0�Ah9�[��=�2�5�����,�_���i+���C�m���K-?�qi�b<�-�a�!?@�3��w"�[^�J�������+��A��W�P���
�sYy�ŏ7j�S�����h����nK�L����E��#��-�\�9Ú��U���-|{s֒Ѩ�y0z�]�C �_@Jn b�K� ��A��a/�F�B�!�Ma��Y'�����G������]�LQ���|��gE���,\6���Պ�E?��d��򄻙���R88���Z�c��5���G��{,]n�M��������ܵ�l�{h�W�2;��+p�εn���>"q��N�G�T�����o�-�m�%�xG
�o�]n���	l��'��a��qB�d\|���Yc�Z�t�x�塳Lr��X��/'>]��59֥�'�w�ƣ����2I~ٺ}���Mw�q�ckg�<�B��<�� �b��ű�G̹�[�(�R����Dz��#hu ;��9�`6.z\��".����X*Q�dP�So�4�K��z�~�n�^�a��W��3	# ����k%��t��S0��9����N� �o�����.�Nj�z쵱�G8b�1?�v~�W��e�POOs!iъPU1��� ݀���e7��o��^�]F=c�59�s�+7�ҫv�J7=���z
��_�σ��y�\���h�_��s|��Z.����*ô�XE�@�L��:���e�P��E�U��2���Ἒj��iu�*�9*���^�y�Y��ja�3����qL%Q~����P�l8���Y����3p�V_�X��U��2�p�R�
J��p�ӥ�-�؞7�;���
����ԃC�B`)��Ђ��#�L.��FbOx�4��w�6�c��Y���ia�W�le�\�L����
NBR��@9��+����dϜBF�5��q�>��&�.{a��n��k��/|�i?ڜ��J���|�pP36���ҕޥ+�ϻC=�;7_!�g}u_�]�(��1Y׵��B��r����Z���aqB�������_��2����<�g�$��mִ�Ga��)�f�"��{(�3w>�R�5��D���t��8���A�����VkQl�"3����}�� ������z�����T�Q��@f,�V	�
�ib3-m�''�)5�4D���{�c�+&'��'�}9�5P�g8�����-;iaJl�$��W� Cǳo��zH��%N=����Iq�>n�0��| �H0�,�X�RhKM�Xۇ��tQl����Ge��j*��x�G��K.�"�b��.�o�\�����Kg+T�Z�����m�Ĺɤ�
��ó��&��)5�&�+�m,5TPY�Vw�~%8A|��=�H`(���JآD�ދ�(�K{B��ҝC:�%X�?� #�4K�������lTH�C˴�t�ԕ�(�<tۋ�$�� �?�R�o������|����O܏0qt������4����/a�+&[.b&����	�Vo�-�0�,�ɽU��-A&4�#[��u�d������y�e*��]�E�����1rGz�D�b���������?��C`�� �̲�	�Į�j�>|e@�T9�K�q-�C���7���C�kcn��DqZ����!d��su&����p��µ-��f,>���{�Q���X���V�E$�%�����%Z��2��<L��f 8}� ���m�E�� ߑ�8�a,�D��FxEu/��/|^[��%�s����J�jJ���e_�i�A-P�YC0��r�wI���uHi����x�X&��t��[��L�W�v�h�RUb�r"��78,r���,��5;n�Sv�VA�! �b
6�|�JS�G5A�7Ӧ�Z*.-��\���#��ê��CM��8���U|L���(Ɔ���8V�����^7��d�Dk�T��L�Pm���v���P�]�I	bf��s?v�'��>�@��0�W([j���έ'�H���"كC}��9N����H'�	ϟe+/i� Z�@�k�V${K����*�����n�7v�:�7����ܒ}�|ʹ��ڙ���Z���t�u�4�h����9��8 �֎�ol_3)���|����܄����p2�ZK�)�u��	>���t����-O�Q]a/S�������\��_<b�гGn�ѻ{��y*-���_���c�vH�}t�Y�\]6��yZ���
q���7����<R%;�H��Noo��&�j`��z{-����_�6.����W�md����G�b��y�\��ˉΈAk[�x�UNa�� �F.��cрM�U*�,//~��J��8���.��jJ���%��y��]�7�+9Q[Yݕ��<ѱ��������\zw��só�@�ě�MĹ����d�}�sB@e+�U��JJ�Jlr��>�I��8Pp~Ƒh2%dֹܽ����7a��|��2% s+���j��{)$��h�;y58��[��6�ITJퟳ1��+�)�QϮ�;BR�a{|x��W��Q��@{BR%B�iU4�߫:��w��U)����M�%5�@���OE�-ǿ�8-��/�=8w&�h����Ѯ�ޖYG��ͨ��%�XBz���r��z��)r��ո9yྫ����R��rŜ��yU	�Tc(i#yۥg4]o�IZXĂ�,	� � �x �.#�Se?[(�P���p�J�yh�Ě��7A]<�H��;�6��;I�t�8��i�w�����C��Y��$�]laQB~~
v��u�=~�)��M=$[�ݦe�h}Hp��zX[I7%tk/�%a��t��@CLz�"Va���G�c�`��l"��u�Y~P(�:�.�J�5���0ې���d�;v�#Wk�/�(�P�e\�J�j����"�2��7��7#��ds�+�f[�/�r��Y�����q�Mv�][~k��]:)Q�r�� �У�H>@�4�3>j���Mp�԰�v�ꊷ�y��M��J�/}i��<�G'���v��#�x��M�nFv]ǜs�FG�;WCr��?�q��W���nm1�f��[�}.�M�w���D̡�4XhF-q��ֻ�,�$�Ŧ��L�%��`{�Bmޣ=;���Ej�2�����SZ��I|��aw>%m�R�hH�@;g�����;ݽ����t��)�{�n).�7��>b^˓�N��`Â��͟/R���?yk"�z�*���t}���� �)2�l���+�<%�$uG�u����&`��c���k�Rً��G���̧Cr��h����g�]�V�mRDI ��e���oJgy����}џ�u���>�閵�!��
0Lk@�&�1<����h���>�l�=��"x��[:��>�FQ��B7d�
���5�*�qMP,:)��Av����E�V�"E?\7e��
*fΤA�V�һ�b���	�$꾇,���a�CU���~��2�N�-��D�Ց���j���e(S��w�ý�~Z���>j�ѠsH;m�|6��ܜ�����2c� �F�ېTNԧ��XVX֥�/�y�KF[����01P��I�S��w����(f�O)0Z��j��-��%�W�����\�^�k�	�EChK<Wi��.M�c�˄t}y1�$�����=���A����O�	��S�r+�T� �|�P �-��t�Q@Ad��{}2��u�xr%�L��JW���ȭbe�:�9�G=6!�!4�l��r�#E$�Rk�m��;�e�wR_�-gu����ۏ�Ӟ(%W܆Z���b���Ԫ���(��)��
T=<D+�vN�;�Tti���:��ć�W��C�t�>*dJ�^S���g3{���*�İcZ*����o��|PD#�%V�b�ȉb��'�;Gv(�z�Gg��n�A������sD�� h�:����Re �D�p␢���5�_�6�ہ���L�)��#|��TOc�:��^Y�M��z��/]�4b�&~lx>|<suhx����(Z๛�y1��������w�c�k�ea�����4�jظ�4�������xS���Ɗ�!1�vC��D�v�ꦼ�����XBo!�'h`���v1N��������ïW[��)N����x�LŁ���Ap$�@T���%(��a�'���4K�lsB_h/���P����tsA�p��D��و)I�DuTodoT~��PJ�[5����J	�' %�v���wcfD�Ds�h�j7�d��S���V�l�\S��&;�5��_-���S�D��+eAsn��O���kV��d����`ֶ~�*!����1�,�˅�PuWL�� #�z�2�h�e�#�Dig��QL,Z�E(e�� �q6 C~��2.�=W6+{U)D@	�H�b	b8��(���B�LzP�w���'εg��9.̔;�~��r�nb ��2J\�,/E��۾5a���f7'���ؕ9-�?J{@�t�{�p	�K�r���̘�Q@k��s��䙫`v�{]Z�6����-����S�R2.~�@��s�x�1xo�*�E�(�ؽ�(/am]��wt
`���5�;���eJ+0)c2&��]&�'Y���iT�`��Ex6.T"+"@�ݕ�Z��I:�Ʋ�5�b��.�JX��.��{#N	��3P�����
jG�#���E\��4�h���)��6Bm�3��^��#��[L&A��Z��3����?�'4�c�)eY��]	�B�O�:a�*�q����Jd�VU��˹h��2[��0�3ZWv�/�"���3?�2�
��*�X���Os�]8��3�Z�k|���r �F^>ƾ뛓q��H ���S{k�n�ɇ�y
����Y;��o�N�9}w8o�Zk��X�*�����	}�!4��j}�Ǆ�e�|	�CA�Z���K��'gj#���`�p����H���N�^Q��!���PwCp+��1x\��>`����S�5T >vU/;8ܦxEX�]��؊'�l�G�h?��W�dV^i��$���F�$a��5l������uΖFȠD������H�_Q�חi���ҏZ�d%:�-%��hĂuK.���HV��[��Q��%Җ��Pi�k�/;��:Lx�,��]$c�N�
�/tW�7��|��7E�u^]�h����)���
M����T�Ħv��	�*m�2�>�&��q�g}jh��Hk�9B�f���OG
!e�&�#[�� ��VX���:���2&~-C����(u�V��zj�e�u�B�יv����HuV����N��i��h�gt�ʕ����P��ۘ�tPŭ�����Y���R\k⪭uX�y�Z|��&��_zLh��I��=�������Be�3l�Uk}UU� '�ͮ�`�[ZW�f��ݜ��ԡp���a��5wL�/���u�u����9�s�Y�ė�/�Р�l��03C@ԅ�YI�Tl� inNأ����	6��B1�y�]���q��V��Lb!���¨��KRb6�D��Jqz�kt�Bm�D%%�uI�[�ʓ������3[�u"��� �#�5U{䣝@����8�|6I3(��6�;J��xW D�r4,t��?M������|{��u���z\��&����0-�������b�q�jkzƨ�9�¹qFo!^8R����T,q�\���Y6�c�VG3�LEk�+r=!\��{�/����o��˨�b��2�	*<P�Z�҇PS䌐�#_�����w���xG��6`�o����|� RO?��׉��a�Bm?	w1�A�{��r:�f�n���ڄ�̒}$�v��n=��r4Spǿ�6��A��	�eh��6�j�������y���]��b )'ژ6i
�XBC��"[	�; {	4�z�cu�hD�n���ɥ���ȫ[�D�&�a���&�(d+��n�⢟m޴��	�o��nctk���!&fR~�L��(��EK\1��6����*�h�FiZ��x�b���Ğ�ҷ�͔���;�� KҿB3T�*(����u��,K"�]��k����Q��800"�-7�ɪ�-
��96��l<�!y��d�uP��Tj��X��j��{X��S.m�$-I7�B ����P~�@�N� ��-j���{���Ø�	�&5�i���p��@`��(!�~l��,�"�'h�e�L�q��3(�&]�����%���)��5X<��
��Ḳ��D��h8���^���~����t�X����'.T�67�>j�o]QA��7Y<�G
� �1	���\� �����,�פ}b�חt 2s�sْ��5]�e/����6�1�HX1�Uf��4�g,����� �j^��JH��=�{�K�1�����H2_ՙ $OH����t�u��}{)D��������;����~*5Tf��B)NqΊ.�4��E�V`k�G��������C��t�A�WJ�f�E�z�̑7�䕂O͒6ρ�Ӕ����y���q�F��]���?����h��)���˝�(Zu��HÁO)�M�q��roQ�*�fC�U��g���=���8��st���W�j���wS~����8X\GQ��wv����hP��D�'7Qe<���U��N녦V��FѸH�SӋ��\�����@+߀l�sb��}t�*�R�}=�͇f+����U�w��ҷ���}H� 6Ξtf�r��kS���B~�T@GZ�vC�0�E�\o����p���w߶dhQ[�>'=NN,?'f����5��U��t�DA�'qb�Y�v
:�瘫j��͈l�)p�j�F�$
d۠޿d�=�͒�[�mq�(G�iϚ+�G�%\�!���R)hS���K����P�q�hLұ+l�>|��m��Yeiҥ�l�$�E,wT+��FܢYC�L߅�G~h8���'�5�(Mx�ړ�TO�w��ʅ[jo��m�5�*�3�f���y�2|8��v>.��~<�H�v��91REiȣ=�G��1uhAG:y���v�z!&�`O�y�����qE"*gd����e��G�!<Bq(+#w�J�!�Rq��M��x7��ô�E'4n9�d�C��	u�yG���ݎ�Ͽ*��=2zϢ�F��2O[xu_�K {'R�&����Y�d�F����y�a��ZfI�+
��4���Q�Y����/Z��l�a*ז�:bf)�ʊ��a���oV;�uC���z�C�I���DBABo��1� ���������:�:���U���> ����qݐ�*/���Z�� G��z,�"�G�@�#�=���{M�L�hY ��'<j;Z*��r�>�����F?��?//��-�'�08�UPX=�PO��E�+|�"��ښ���2x�q�&{}�Z�@;=$�8TU�F�P���uv(]5�d� �?\�"�c�~�f2�GVa�^����ثգ���כ\��Z@��QX������lr��P�\� F�a�#��R�=&#�w_A��<���gd]����P��0][C�ZM��{���,G���'t�"����-�W�P'm�`��Δ<Ϻ����h�f8o�+��"��?B!R�_�;x���v���eC�
�x��Y�OQ�JBX�)���SqԸ��{�\[��������k(�U1T�����{|���,<2|	� :<5jh7���˴s�k�h4K��Le")1p��ӽ��x���ro_si}h`����Oc��W��̹�٢]��#�oV�Co�~{�]�:LdP}E{M�
��w�
K�vņ�� =�&6p��>�0	J��2)�����r[���UD׈��,����Dŵ?;b8U�-��Nũϒ�i/pi����_��a�>Ս� \�8J3U�����d�:�`�=���L�kvba�vzM�?1���d\*z�u���{��ݷ���r
Bt0�Q^r��7��u� fg��W���-�z�f��<_(��o�D'~�˷���g���)��Ol^NV���]�h���-os��YJZ>ɐ�&�{�^l~�"�l���k�I����$1yud]�!�*��B�ǵ2��ej���Vy��1�\��.�A�Y�"O˖|��u�ᑮ�&_=?�R#�,�qB��ٷ��X��6Ě��!l������B���|�!�p���g<G�*ب�!B�fm���q�.xx��5�ZQ���
Bi6�B��92�A��ev�#����oP����,ȡ:�L�#�`�:�}l��Y�L�1�;i%�ɉ>i�e@�S�b��^�U��1A��㪘������s�J��Y\:�l�r��Z�&0��Нz������N{���K��n���)Y�f�4!}�捎��tR�#t������7�'2@_��zuY��B~�����ϯCK��gJ��h��84�J�At�zg��ݽ�Ԛ����Tb�ji��o�V����[��+g�<�$i}��\�Y�N��D�80?S�Yh��$�>�b�G� @&�	�;\��xr�!�9�KG�#@,%��WO�#�i�nJ�����SK�ӭ^���}�W{lY&͉����s-m�a�[���\o������Z�+_oS��1���%��T�/ܚg�a�z�`ܿ�z)�'��)UA{fKt��1�b>���e$��\���Nq�L5}X�<�F�in��� %W�^���0`�>��0�j;U���W���ٮ���[n��$�l�,�<Z�\��n�ʗ*������c�T��
D"�l�~�9
����	�al���f5�>3������G1ߔ:�� ݹ�}t w���gF����FnSE�#4 J�z ����=+��3>i���aM_�N��g��r1ظj�O�/_e��m�X��S�����|I�R}_����X�P=EW�`��� ��U��H?�1z-�J�����b�=c�&Eh�a�q�烧 ������AvHu���:o|J'��(��p}='>������Z����VB<J�b~�}�[B/dx�p�2�ݤ]�dd	1���~�
��,Ņ���,7'���hG���__�~<x� ��@MU�t킨g]�U'�L��+9LiE�,9�	�5�o��︶���f���9{�s�)y�����[����L7�8ݕ�<����{���`����JÍ��E�e�&���E�KV> ��q2�a��|r�G@ �n�8Z�o(c�NCCH�+��P9"q��3��
Ey'cf�]{�b�j�Q'm>��;)�|Qg-�p�I�����XʎB��:��<��K�����d���l,�B�a.�%A=�h=�٥���61|�E䶫��� ,Q=���׋V����l�	.sw�j��k��"���#qwb H̎��j��i�T�n��6|n��0W�H+!{pswF+D�?Z�m���w"�-s_P٪�
:I�� ����al�G+��@2�"� _�jѤ��C�vW�%���;�����e���^�Ƅ�w�J�L��g��**�p�Ժ�Y��������Y�*kͿ�
���>PZ>�ު79ܰ��� �CY�8��GT_�F��:iFm�.w�a�3�$V�oY)ݠ�/����1U��Z`؋��C�G���ﺵ�@�����?�]����u�C<+`[L�`���]�Q�%���'#�,^ja���q��A@0Xg���LEHW*��G\M�zg���J��s�8�^M�z
�)��U���F���WkY�l�������`P������Ȝ-t
����U��ۻ�����Ob]�$�c�fV7�H�*	(���}ڈ�u就V��E�("Zn�+��[��ev��A���A�\��r�Gnk]��� ��^��sj�A3;�^��Qq���5�yx�wp�FS�~���w����Z`��h��� �7�c�^D�����ED�0}x2��D���i��hFRTچ����Պm�tY'00�ո�o��2��I���#-AT�+���9�A��!��k�����HٌN��I�:%S���
I!�
iT�L:��$=}�u�5�Ԝ��  ����2Y����3����w��_�֞a����U5ץ鹬�G���6l�x1�<j6��!�\��� F�\�����MN2-��_(�^�̽��q+�K�����"� �B.q�k~9T?��͖䰐�}�>0���ڈ=�n<^#�n)]ɵ�J�+��Vċ�#3�ӆ�c�|��#pe���7����*[�ʏ�L*�C�Ƚ������vhƠnt�[w;@lZgC�������/�qc/U��-�ak���<���)I��&�ѩL��?��_O���;���@)�6;Z;M�_��+���沄P�I��Z����ŀ+�ny,��yy	��-�f���E�ı�ͨ�}�:��փ�����yt0�j���t�Õ��*J�C��g'L6;��Jn��3��߄1��^��Ov��p���F��a
 �����!�
9ͬ���|��oG�C�&�G3e����r�����P�ͷ�wP ���&Q���I��x�+JO&t����@Z����Y9F�o�b�Q�pw:_�Gn�n�D`T��u�,3�h�L*��DX�!�/-&r�-�"�����|�k<���]"�C@UQb^�Lv`d[�������������r��\:G�W0O���f �����������2�Rc�<!kM��x�h���ۆ������SAP��~�����(�{�u���y��@E�ƃ�]a��� ��UL�n�B��tta��JM|�ׯ�8kڔ�#y�:��rv �I��a9�V�.i�Qߴ�o#4��Z�g��!�����(z��|x����*��q�@x0
?��x/y~������q����=�U8j�`��΢����C'����JZ� ��Y�]R{$�2�;�EbE��u���\h��Ѳ����L8L�}1G��we��Ȝ��|����ѣ��|��3ͤ�-��#*ѹ��,;��Ҕiк�-#M{@�5�d���������G����>���EtZ`�G8�B\�K$H��0i��7���XQ��FD�J3�DE�&�}H��ha%P�ﾾE�Q��^~�->�<�����GS� �3n��+:��>IwZKM(�4�6���.��C�B��+$�6�b����Z�y�L��}���ŝf��^�a�gسhTцO�7�y��;ݠx�x���?/����� �#���>9�g�v#����]w�Ÿv\>�v
G��$�4�&wܚJf�)�����7�5U~�LFt�ݬ�l
 �+��2x�4��sj�e���9��Z��Z����HeT�/�~����(�h���LR�7����:�����t�4,���yμL�����C��_�}ĭ�"Ⱦ�/��r�����]��ÞK�(Vr���N��O b���7E,�(ja$_U�4C�+�BV;���g�� ���m� ���u{�s������ {1-p��0��W ���y��	�Udp;~P
u���˾�Ü�,��Q(������&�k��TzT"f��C�E��K�&���4S�vN���¿�G��:�^�ci��y�n�Ƌ_�.Ξc���ҭ�oƛ�Y)��?�V�*���Tođ#��k��G�/ށ�.�ֺW'��$v��D$ 9��@ ��9�6�i>�˂��߿�.ۄlXP�2&��L�
'׏Yc>ݭ��]�0x��K}U>�^�G��\_b���
a QG|�P��c4���f#+Z�|�@qwVdd����%�հ�誌W9o���S�,� <E�'cM
���.����$������b��3G�1P|]�dÜ��N�E�ua`�U������e��?biӥ]�Yu�5Z~4~fw!��-�0Jp�r���¿W�s���
$��y�>.ƿ2oև.Ȳ0�quE���0v�9��`�P�n�-"Ov���#��q�֑x�1�x�Ŵ:1��6h	���ðK����<	��)�s���m��_����"��&��i㸧G6z��Zw��}q܄0�2G꞉�(���d�U����Y�t���$;��͑�a�o[\�K���W�b�v�7q��Z�@��|v5��Z�"ޕ*�H0�I0�����".�Bi	>�6���	�v��קUӨ	gj~��E����qj�&!Yٍ�Ggz�tڡ���x�i��4�1�{71��.��*�{���t����g�����m�4�O�U�����㄁T|�Z�>R���_3]�N{E�U�6��U	O|�o<0'��Ma�%m��H���툓�Z+V��FL�!`�=yǧt����񸬶*vE���H����Ѧo�>0�4�ϐ{�H��ݢ��e��(�<#'#V�j�y�����H��p�|�v��бib��~J�ʴ;ۼO�X�*0�Q)AZ�;����l����5m~� ��%L"�����س��I�эϠon�jd��S��ՋY}	������
�ߑ]j�l���`ܶ�f0�������[8��9�5e[���q^E��xq	U,^��b)�U�b��푯��[��o�[�BrDO���J��`�����X��hF2wv~��>6`d;���,(����|�����d	��������<�m���� i��V!�;����-bl�%�X��f/S���͢�W���m�����;�o1dNd?���q[:���Њfy�`���ta�Wt��y���:7�O{oRH�j�t��p@�_d(s�E$��޼lW�����:L�]�r|xNo��У����(�����t���IOˮ�r\�;)�X�{Ů:R��������k2�57�}�8���F��Ȧ���B���_ �m��}�_*m`UB��01�r��2�;U,d��+�M��G��g^��4�T�/�W�/��p,���{2LH5���Ωx�3���v��yqDS�A��\���{��������Fe�nb$@`L5�$�U?�R�(W\sk���<�+e�d/�:���Ǻ]En3p:��{Qf8 C�N8�%S(�k|%n�J�*w��&(�¤�,'ָ��j�UPN��S9�-̘��EG��k�'i�^<5�C�"~���s��s�A�hRm�T���
zaK����f�D�
r��^�Ji��(b,,*߉�=�g`� ]���c�0��	�=$ ��xX�K�(�-��JD\cb��WL�f�k�$T��`�� �a��
J�$�?�{�Q�o�b�C~>}�������'X0=p�'CRD���L��~�p�3@����Xzf�D`ixxN���
cW�K�T)�Ԡ�UG�)B=.��՚;���7�J �qd�~��o*��n�/�d�3o|�]t]��͸��p\����+J8�M�����I�L��,n�	Vy��g�L��>�$u��n?�#�U����Ǚ��i�0m�Wo��{�}t,���Y���W�0��4p�v�; ��귽�Q�B�Q����nH�M�O�@� `nRP��/g�QnT:���dI[H��F�
��d��,���;���)��_��~X�؊>�~B�A�g�D�`~2��\��i��à��9���"�_
�Ƈ�EH��[fc��
���B����'�� /G+���	@�@��z�/������W���nm|���Jj=��lÓ��{j�x��=[�Z8ۯ��u��]\�ٕA�鼳�V���4d����},��/�1GPL[���툠Cֈ3�W��˩I"ed��ߗ�tL: ��������+r�اF�! �̐��4�%=��*�2���,����R+/[��7�Nd�1�g"���#�g���y���s���4��
4&�"�ҙ"��4bɋ`��?�h]9w3ݎ߈���
�*�@ȳ�����&^&W��d�2�Bv%��y;��C�6�I���J`�|[�5y�) ��L��X	���;��(n����c�R�sX��m/	+���n���Z���o���_<ݠ�k�F�A��Veژ��?��OA��C�+�S����~�)��ѧ:+@ٟ\y�P���%��B��
P�����.�	���t�|�y��, �����ȅ4�9�q� �oAv�eW��J�v�������Hjk�Ɓ���S�&̽���L��#Xld�5�r�wY	������!�	���y�v�<�S�� ��Hw�ު���񑡓I�e�T^F�Z�E����	/RD���+�e���˶U����h+R~^�2�4�4����N�|���/�O�H�)kF��b�H>�k���:�g'p)����A��ʃ���.PJd��~8�+�S�AP���R�P*D׵[(6���;�Ŵ=�\օ�&��t�w��xD���n����55�nY�s�O�I�!;Hm��O�r�2��	��� |Т��
ͥ
BIu�|���7 �E�K7=�⁛Q�Du� p4�)�ܾa�*K*�L�?o��	��c�ℼz{��Ҳ<<(�.ZV��~�n3��P������k5��!�_��\B���O�.��շԢ��Ro�l�*>�^����i��t�����k G�v\���Rkc�)��
1�3��
щ�^�(��+/g�M�R�Mx��ѫ���
�)X!������HmG���K�����6F��/�=^1*tk6`}��'L��^p�bE��h;��e�?��K�7+5��I�g'����1�o��YS�n�^�?��=Y B�8�t�K�4N2���_� h(#_~���[��:%���%շ�^���>KN��#�$��=������%e�$[��
�仟K�'|%YR�E�j͞|z�B�>	�ͺ߁�-W�'l�M9m�dE&)�:�1 �P�����=f[�O��N�h+��{�p X�DI�z,����L�b`|���N¯����֘��Y축�B��^2c��� ��s4m}�D������.m�"�(" o��
����Bbȱj!�To	�5ʻ��h*�Dx�|��T/>�����4�bLH��_Zt]��:!�D��3��LwW���5�2����y�2��Ym&����	�L0 ������A���מ�'r��*�"��&����J9����Q�o7`p[��Z�.6·H)C�:�Q�1�	1����+~}�����B�%�RT�u�sP-PL���ؾ�/��^_mJ[_`���c�d�G����\1��K����~�"a(8@�9G��t��t������<Ki�l�Ǎ:�o!���_�e�
0��4c�{���\N�2�kg�.�+����Z��|��Ub�'���{GS!�)�f"w"E}ݼsO�+�E���GG�,�#��tM	R���Z��˃oPJu�LU�8�W�R	����/�	��"��ҝ��-�+�Ma|�OH�������O�,Kb��`�]��@@G� �s�d���6�׀Tb�!|n�jW�0_ruN��>���Xe
�v�d5�.�Z*e�9�����n�G~���Lq���,�\$m��n�`�;M�
9ދli���'��a`ʽ\��ɏ�Q���X]u� iU|)�Vċ.�nt6�WAƂ�J���V,7�G@YC�(���!�x�+��eH5��_���v�A���`�m b�?ˡǃ�
�#�5lZ�	H`�z���`��L��;��(e��)P!�e~6�s.��s5��a}l�o��6z��j�p{P��P_`���2�������5� Y^���P�MyRIZ����5M;��,hF�fwK���x�©���J��2Re-S�~V ����w3چ<�`�f�����""9����Z�7:�_q�?��.�}v�c��C���87G�ފ�{��>���v]�����t����v~����L#	J~���F����x�����
P��C�z�j�u����G@>b_�h;�nr(��+?Ĝ�`���� ^�z������4�W+��3U]r�7Qz-E�9<�o���H�Y�͟�IQg�hc�oM� ��o���]9~!P��Dޠ���d(���UQ���9H�q�&[/.i��mM���o
�����
�1��̬�q#k%@K�#iZIS��l���5�^�-�PPr�y��瓊&����h�=�Ll���g�y�=�8_$n I���ۥ�opt��}ϧ�I@��f&%,
��98��R+����&4����o��5��;<z4��:���1�Xa�.�ӭDqE�N'��VT�d?�)x1�~��8�+n��ji�iπ�w����
��B\;m�RF^��,��!Aq;��8��q�sQ�R��R��9�)Kf.,'�����X�g�|]�7���F�������<_��C��s8pK�4��XN#��g��x���@@�����*��/nvp����2&�����O�<G-V��D�¡��z51Z�	�0�S��n�؛`oY��*������h��'�Pt��0x�B��i�n��rb�ҋ���<���e�pɴ%2�m�Z`BUN[�ض'l`�"W�|GV@�<�\��Ya_�e�ƈ���y:�Yu ߓ�')x9vA��$�P���O���<�s�-�eѨ���K��Ol6�ˀE�l�W���^�.�w �p�n�A���t����yx�2��}��l>ќ�8Ѳ�U	D��3�F��<��A�nfGN�g� D����ܞTm SѼ0�~A1���.�Yꤗ8(\uӟ;���mm����@ՙ;;Ԙ��Qem8�I _ǐ�hu̽p��s��՗f{�����y�Y5� E����֪Ԏ!���T�W���(�V�J��-c��N-���A@�W�}e�x�IsH�B��zL��5�#{f.�qBՔ�0�.idm�\ۿđ��u�>�� }�>�fU��UT�td<001�iA��u�5��/Z_{�4a\��U^�XB��߉3����X07��lч����\��1�Z�����u��n�Á%ΧC�h�Y_��;�/�ļү�mî\��0$���/��]5�㩅=����w����%�&T��v"UT��#�c�w\��?o�	�_ޣ@��co�q�ɱJ�o%��A�<�n��Rg�A������c�(�I�ly�E�խ�lK�㼪k�?A�$�p\L��O��G�>�S��;g�
O�3�R8C�+{��T�$��E�Y����ph-*��S%�Sl\�����o�:���c\xGQ�����zdɕ�}W��b{�<���g��dO�� Y�Y�	�.̼�J���C3T���ւ�`��@���+X����տ
4��&����dt���7m�n �v��e��jlmѱ���8ɭ�V��{Hʧ'������G!t���\p*o!6���h!}�L�ȡ�h�{��`���S�q��]��@P���'��oxD���a ��OeZ��i��b�O��^���9IB�,�+�()>��r���L=�H4��	�X�)�$�ip������/r��}ځv�䫣��P�x�@:Py�+"�-��A��S1�  ���M�u��x�����&I��q��P�WO'����k=}�����4=g��|g��@�J1������q��re�@8+�k7���.�Li^�':�v�]4C� ����v�)�y�C�Y�O_�5�f�UE�1a8���8[��^��:]@t�C��AǍʑ{A��M�P����V�T���n�Io ��N����߲TωmM�}%�s��f��Xڿ8���6A"x}�"�˝������W!I�'K�����k��v����F�ܣ����#ޓ�t}޷,��`��t�����tn�x;���>uu�~���CZ+��t�=��1��۳�����-�r�q�7f!�4*o�s��*+���L;��|�M�Ĕ�ѐ��=����[��T��Ψ�ݦ���46����m�2~�֪f�/�+�p��;��KL;��ԫ
X���!y#X�w������,����Y��f��,z�	 �����[��O��6��Qĥ��9�CIǟ�������-���'����T�B_`&��gT��n,�~{�R1�����Q�I�g��N
r�����6�dG� �a����9��t�S�F���x@@\�2��书��tD�Rb�h<�-e���lƔI�DH.�1�zq#�O�|):�����`Tӻ`eNA�w੻�����o��p�^��������ab`r��Z��>�Ш4z��K`����N>z��բ�.bm�=ת�Q��c���"��$��x}
h�	"��I�.���:���ʐ!L$�� 紗2.�%�!R�_L���ULVi>ۀ��d�����ո��KײT~k�B���1�cw�!�y[��q���t'�tmb@O�eI7'�3r���#��'&��׊���}tk�L(}�� 9�~���2��
�E��?���r1d��~����4ZN�٦�uR��G�a�cE���J�lCY���TGo�P6�鏏%I��N�H~aꛤ8k��t�K��%h�KX�*U�T�	�a���n���(�~<44H4{s&\&�g�Z�N*�8��1�
E7���%��ve��w�&fgB/��WB�\3#hS�{�X�bqs䎀fiǍ�!ױ���y-���9gƻt] x�@������&�JFY���P����=�^.vܜ�B:m�"X��.Q�[�ܞT��f�-sЙJO�g}���,y�7Ģs�9WJl��y)s��}�]@�T�V^P��	ޟvv{,&'ϐ�q��l:S�O���ZF����q\�A�u�\#�n��<�k��м�l�f�gx\͞ϗm
�.wT����3���� ^��9�	
*��?t�kjX!�C��HG���-�\0�r���+�rĭ_3
��"��#;���H��x���g�#X��Ň0�-��~5P�I?�＿����Z��ô�!�P0m=�\�����BY��l��:�)CM���`5�+�LR��H>�� �	�F��+��f)���3��۠�^Yg���.����h�5u��C4�z�vv\D�ܵU�����\M޹Ov�nƇ�~햣�y�w+�lp����n�͸!ֺ�5���|�p`��YP�.���ga=O#Q���wt�{�H��:���Z��K�K�	I�ǒ�ɾ��T�}L�W2���f��{�X��)#8i[��z���by4�@�Q�k8>��,|���sy�V�Y�C�ػD���Xaa>�^��r#y|��Tj�$�]�ն<��J��t�!�n��fH��s��D|E0���?�w�_T�ߧ�F����װgg1z?�|���[��z�?�b;�P��<�/��M��gІfZ�58�K�x��
Io���T�ٱF��ѷV���{�������ZE:��h���ה��*�ouE�]_�
�8�2�L�Yi%`�Ǻ�*u��ySo5Z_�N��9�K�,�c��^�Wc��a�,��y'���*��!v��]�����m�%Ҵ�7`M]�p����7m�A��٤�Cy�aΖ:�sМ��%W�-U�XQ*�����T�r�A*� �V�o�&�1��p�#����/`݇���8,m�!"�pG��9�/����7l�̝��2#-=\;�FѰ~����YC���:���Z��W��zܯmK�~�x�[�&�5ojs�i����;�Gv��F�^�ݾ,��Z�9ں- �Ǎ�ܗ����}@|�ROs�#c>��s�J��*=h����+l��`�~���`	�iJ3���P6��X��ԟ�j-�3���^���w��,�z�"�^�[&I�;���Vk�]Cɍ���������ް�3S���鉂������;��Zs0&I�w�G��y�y���}�� 魊�YqS��{	��,.���(����g����4Mѥ3W��I�Z�5+Z�㷃�n�|Q�'n�^8�"�0e�Z|Z�dE�����!�}ł:c=��$�al���^r���)�TXгِ��zѰ������ ���P����s�}7/���'V�ܺ�,w���R�уwr�:�h ��)�I����� �{?�z�im6�#V}b�+9�a4����%ْ��LU�?�,O��V
���R�mz��[�%F��㤨n�4���f�0����d3��tq�N���H<��J�3��-�p�wA}z���P�q��),����5x�nX�,*ٻ�8��|҇	�FA�NC'G�� 5������X�"dt<fM��.K���4yF��Ϛ�	rn���^t[1�����d<\ۃ�!g$��/~��F�G���K/���ŭ�0�ᒎ��(�x/Z�~�o�<�i'70y+SZ}�0o��p��L��¦����O����������$E�	B�)��ɠY��9�~�`z��~�$��k�6 ki.C��wT����hv�4RϷ��S�7��[��c�xWzd�C��+��]��e���;�Z�I�kB{Kv���9)TnDM�wγr�����!�v[�Ѣ�S�c1�i���
Q��&��g �	ޛ�m�dAA�RWҋ~�`[��l���,��sW����t{��#4W<,�k �Qp��749}�1~���j�`[������ҿKe0�d��.�5	��J��htx[�Y�i��[�	�.�nN�·֚ɾ��>B�pl�(�x-J���9PH�`��~������)�gXEf�ߛ�&~���E~�Ii'G��ǟx���f}��~�� ����sf�ͼ�T^,s����Lq��@Bǅ񟶧�[�HĿ8�@�X/)Q��S��8����&,�8�Q�s�3Z��I>��"
!.lr8�Ngg���/�d��A;�H�Y��✮Uu�yJ,_�w���/1L0Kr�L����=뻞ه�K[��1�2��]GSSR��|����޼xv��R�=�<&}�!�`� /�~���[z�
��f����֑8E��Z�a�+˫���(�C	���ȉ�pL��x(��5���(������i�V�o*
�7�=��%����L��a�Dy������s�Gr�����k\}r���sƲj:--n�l�2L7�|t���2`<B|��c��*
x��x�U ����s���C}x[�t���]��,H�Z�i�wِk-�.�cՉ{�4gt����Z(2eV7`'�5�LrR*l2����G�5��J�����o���	~JUL�.���-��;�RcZ�Q~�N�7�n�]��4#�ܮ]�#'�Xs�P:�b��f�}C�&����/})��o	{��V_��+�Tt]�-�L�x@�6��@t!
P��c;�d~���"�-�$/��8;qY�����[�4�%��6�q;�3�ɭ����9U�/}�����x8��F����e��<F���	j������P��/���P������h�^~>0��lQML�t9���4ٻ�l��g���K�|� }��X1sݎ�֘�JiFOH���C>
C(�,4�J�u�g_2a���)��rp��<fu-���^eC�z%�	IV]EE��Cj@�;�q�3����A�	�{�ԥ���p�-~B�SNc�}���<���ɦ��/v��	�'ʯ%��C�F�"�,��?�*�+:3f���,O[Z���3Ա�]���$*,��}a7FD�=��FbOk#�N��=�s]� �^�Q�Q��JE�8B).�M�>5�=8�Tϟ�2������Iq�:��o�"v��&:<��P�X��[mH�3}��[@���Z���u>E��u���E-�v�Dû�$'ʙ�OM�]�%�s/���B��&F�aH�c�yzNP�V1h��M�!_k����r��<��
qZ�̀��1	�&����%�!�&��4�׭���ɟJ^��:���K*Dx\� �Q9:e�w��5���Q΁��in�̶<Ȱ/G��;Ir��� X�*gUa7���w/��Ͼ���F8c��w�o����5�ln��"���G�%}�����**Oz���eG�w�rY���j�0�#���k��g�A ^R���ĺgG.6�|�ص'3�Y���<�ړ�0Ġ2t�~��e[f��O+%K��@ �׋��_(b��g��Ί�Fʛ��ź,|���sw�y�=�~�!�L9���ڱ�x�Gk��R����� +vܐ�s��Q��	m����(>��f{�ss�L8L�S��b�I��"{�~)c�QD<v\�I!]�y�k�ë�@�9@u�G�̀q�g�