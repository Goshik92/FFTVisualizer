��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��r��U8'��q�L��)���� ��I=���5���J�)ȋ�Q�b`�ۊ�=��|�JA��u��aʆp=] D��V@��!\��j|U*�sՓ<��0���1\j+�`ڭ�L���oJW���3��ZV9ls̰��gm�|�]32���WIZ�T��l&+�d$z�;^�Y���0x�.��0��ziAYU��:!���O��뻤���Њ��HF�	�u1��$�í:��-M׆�	k������� �*K���̮φ]�{���E�j��i�_X�߭"�I����T9���zs�ؠ2n�1{��^cKMkt��wZ���H�=�9?ҕ�o�䝔����k_�d�8
�_5�*���q��G�X�􇿜���GJ��!��'��x����'O>m�$�J5-De1�Yf��m�>~��+d��}��m�f��Y5}���^��8v}��P�KD����@���0��ߧ"ߴ��)����c����5�nD��^L0U5Fa���e�4#���> W�5<��c�C��ܟ#,����a8~}
��U�����,�p1��f�r�d[��TF�)�SMͤ%a�EG��<LW`�\�f�ޱE�ly�R��_����f��`��<�e�f��i����2�]���
��f�D��0<4��<!)F���q��hc5���|kr b�d�~ԣ�-��/����]�<(�rWM����p���{��"pCև">%�~>��d)Q�fDuV���sI<��E��l��W��e|A�%�j�Ȓ���!=p4�D��|	�7��T`#�[���\z(�l #�-&����#�Q���f��i/)h�y�c�,y�c���	x����o����76�_�C�ئ�d��j'VĔ����j�����H?��'ԁ�On�� 8�#�À$�q1�,�y,�N	�F���)�[��Դ6C����~UEo����)�u��7L4��Lg��d�j���h��YI���g]�[����*-`�Ayх��d�󊲫S��,����|I�h�y��|ѱU��	6g�S�5�"��^�a����D�\���AI�%P�P'��)�~x��X�Up��%����ppp��sJ�A���]Z�-��Z3�xD� �y�`x2\���*�A�����D�b�iD�JI6s����Z�k����M&��Q�5�2c���o�C	��D�Sc��F�Gm�Q�K�]?~`�kݛ��1���;�� 61�����O��f��fF�E����s�\�8���RW�d�>);V���3��wHwk.^���o�n���2v9�찁D�@�,�\�z�ܨ,<
��hY!��&,��>Dr�%N&F\�Cx�aiV�b��E�sm�ᯊ��ץ%}�'���)����p���]�j>�� vqRƤvX��X0U�σ�1�>�P�?�:�x<jEq����+��P)1����Q��j�~sH�pw�DI.����m�:G ~+���"�ƒ��)e���es��@_:ೞ�^ԏ�;��T�����ˍR�����#�0��a���"ڇ&+~�uR] �to�' ����2퐍��EC�o�u|˿u��ձۇ?��i�8̮u�[����L���Y⥡����_��&�h�������w|j._1H\��1���G��1���^ǻpdEP�=y_E��,���b�t��D�����5��ph-���q�;�(�7y��~��$����xC�Ѵ���}ǄEm(��	�	K$%ר��I1�Իx;?(HɈ��H�|3��P$4����(�O��ڞ���~9�
l�
�]�5D���ۗm2��tT:��_:�1�m}����Uʀ��@@&��r2}x�M�s"h��^,M͌!)�'� �P>��g�='�m���s��|r�!FyE$t�QY��	9�1��%@�<c� �X�;$�- �"���T�:,h9�l�C?�%�o�b���ILA��>��+VX�g[�W�U�ְNV��\r��;����O�\���6D糌#�/k:N��Ȟ�6}�I\6{`���]˝�{PYR�p��\j6�$o�İ7L	�";~=d���#[*�_4��,Ž�gQ�}�#���c�rl�'.R�	K������HQ���	���{d��_�ra�6/��D9��G�d�j����h�dR�]��s��=.~�r�^��u��-��Sa�]U��S+gN�4'��B��$�95�;��6b���58N҉��������Ȃ*����<�P�N�ZCK�z`��@lզ�lSv�c���iE]��m�g�a^#rZ�)��>'^�~�-�9y�'rP���铒jR�l�5�z�����φ�N��%�Q�50��FJ=%�K�\'7��R�F+���'w��v|v����9��/3_x��!Lj��f�nu6]qf^!��T��讴��R5�b8�"�u+{��쟫%��#���-��'&�M��>m�p��Y?c3���n�:��T�+:�-k�%'�Dj���5�����Ot0<�4oXؘ�� }'��8��`��<NAz���/��f�n�>�uT�Uޓ6������7�!�0�h�rZ��̽���j5�!�߿4~���2�T]r��>�� �|6m{eY\�h�#��bȹ��~��G�˻~ϕ(y�+�FȆm��#�9��Wqgͤ�3K��<�K:A����bz-�KQ�
�7H��ˬ�K�C�%M��� !'6t��	r�ܴ
K"L����f��^**���mA���^ 㡣VWˏ�r�������N�휗B̛鯔EE��3����D����|��jȢ�\@����A�-�f|��u��iI
fK)QT2�u�}*�|�9��!x�{
Q{�!�uQu����U#��2^	z��ܣ�C�p�wxh#c�?�*$�iV��0x���:�\�G�d���Cw���h��	Ԍ7qW��yg�ƕ��G�q3l��>�hwJ�D����_���B�~�b�yD8��?�8��nRl_�/�#����ҷͪ%!�	�2ſ�go���D"�S��T�{
�����µ��٥1	�P-�
Z�4 �:������,E-O�\�ԃ;w��oA���}�D2:�����
U�M�XjB�I�-f���M��)��u��J�������P�|�*G*}��O�� ]��=�%�-��LRV�������$��v >�'�DB�x�ffs;%#F�S�k�M6�Z�S<#}��UT�d��(})�77?2g�N���8B�'�)���Q-�Mx۹r������?��LAI� U��ٔ�*#zpמp�o�T���.��hp~�H�Y˨�J3�G6;�QM����������fq^j@$���))�LKF�t���0����a`rE��ua�y-	��}�>��n�2ECQ�T�W��</���`2��"��!k�C�.�wkvMx���*�W&AE�'������Jֈ�f��񆆉��%W~� �R[�*���^)�a�BR���]z$F,tH/�FU�&M������g��?��[��YVn�U[*�J�D�C*�.\v�r��.�$h�� ψ����lp
��e*j���q#�`�2��h�������)��.V���ϣ�t���g������ߔGӑ�N���2�g��5E���.��qu�]��נ�9hB+����LL��9ٱwd�@��M9|�p�Z�����S�.�i��H����9͇D-�k��d�4�	�c�5���r�t`��$GZJ5aU3�P�y�H6�izS�T��"ν�d���Wnz�Ϫv9���l�M�1�3��vH ��<��w�$�|�R3(���b'fp����q�s�bdڐUhW����������\�ө�迎�dp��&[��}��s"cgמk�2��D�r����:x1y1Vo
I�N�,��h����2I�4�J:�c ��ҝ��������	��<�}r%�bu̑J�k��Q$FU׌;�����4H�99_�ι�Æ�ē�qLАfM�����ё�N|�2%����vi��#�K��Pݢ�( 2����4��Т�N��o@p^2I��l�Xu�Sֈ]UT�=���x�D� 3%��~�$�Qfl��&Y�������w��:<+���	�;�������a�x�v~�����?.�`��8�yN��5{����A�*iܞ�L��,c��b���{z�Z�C.�{�h�y�����<Z�~�d��suk<wYѣ� /wF��*�����<Z��h����5��/�:D�{ >��2Iݵ�c�D��b���mN�e�0P��Q.b�]�P1�?RǞ�dd�����:7�ɣ}�e�2bF��b�ʕ��F)n�s�U:��0��-=�����Y�\�g"�ȩ��f�p��$�s&��(��K�4�W	�ɾ���)]gBJ���f{$�Q9����Qr��#�y(?�0��C�6�k������~"���N���%�a2�����BB��ȇ�/v;N��G8����*�g��Tg�(-�xnz����������RYm
�[��!���@�KD��p�آ�3����?��g���F���\�mQi���5���:	I���F#��9>k�V�i5�u��
)^���qv��4/&��ۊ�U~�6:$
�;��M�Z7���[5��bD��f���|~