��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��XMXl�M�x��ֈ�$�(r�\���a�C@o�V�宅䴨���ڎ�Ͼ4 U�ՄHY\�YH2�U���i2��V�l��rN��\��z����\�Kw.��p�o$�MM�q�A���M��B�l��B�}Z�$g��B�M�[���:2���i�QxD�"\���(0�{קR��������;�s/r@*�2�N���kX�x�Q����`��,l���Q�YvDX���w�����:;a�� �_;�M>�`�2��`?�]��4A�b���֥�Ҵ� ���5�������˚]IG���۷��MF����eP����C>�Cqi�w�V 	�*�|u	��g��tǈ6���'B�V
y�Q"�g��,�ww�G#��]�K��\����&��J	��鳬�b'tOk��Qb�J?5�W�J�E�ѷP���V��ψq����Z��BF��.��Z�,�����1:.���y�����2��N5ޢ�ժ��&.��ɒÅ��T�����߫��s�}9�O�0�?^�e4:)�wK<^�;�P~�t�������Mf���k��������.mV���]�w�P�?Ώ�(`v����4\2��g�r�]8L�Vmk%��&eE)��_�Z�AjQ���� oc�z�*���kdG��T!��z#�^b���T��~JV���d�艹�lCЙɎĒ�ܧ���Cg��wp�i�<j؜̷z�Gq9L��f
ۥ����5],�Ok�.�$s�X�PU\�3���K_�/'���E�'�ZC�����Hԓ�	$M���n^YG��� �M�eF9�Ȥ`[�׫�²} t���̎Z/5_�QX�O(C|F4s�W���6���,�e�E6�:�k�Qy�.7ro]����d�a���K��Ы���+�{*Nr�kR�1F�^�P�Z�j�j��	�ȹ���r�f��r��b)`�=�~)��a���3�� W 9�`JN�R�y+	�����H���o����dhLg�l;��u�p��7�C�%L{�ڱM�(&���u##k���Ec�Y] ��V��lN3�ܯ8(8Y	�O��<]��h�X�4�_�K�1Q������J7\��(����Z>��u����(*Z&Aҟ�H�^�������X�D�Fڒ� �^���&xE���^U$q��#���R�v�b�ߕ@����5�����I[���f�W�
Y�bz�°d0��/ܕ�7����.��~Ie%��rz��:�o::ƪ�����8f�-�_��]A<�W�Z��%�b��j� v�b��t��/�"؇���k��l�G�����b:}Z��ʹp�Dn�]��〱~4^�./x�d@�;1����W���b3�� {�0J���O�SEr����+隆�ٝ�ۺ4���ZŦ��i�e�je�1�~\K�6�aޮ�C�f���4���I�=���7���Ѧ�w#��w袎r���=\��I�+���S������ cOS�4���`��#�q-1�_��V�e�4̠a70+0�.�������ZZ�*�'tCpZ��4d}#�1a��d��4г��D1�k�:��U��j2���/f,!s�Ϟ�*	H�,Vc�.�7=U��4eЂ���-D����߷���TF�Ā^ڬ��te���N"��ɢ•��^
�޹x]	��u~��	Ӂ�4F�@Lͱ�����ړ�;���\ol��n� ]D��S��a�)���^<�m� �S��؅��seB�K�Y��T���v���,��E����I��L��n�,K�h��g�V�ǧ-��E���m�ȧ�AU�QBX6���+C�3�m�Ha�_���J���u��A7�BE?W���E "X���V��.�(R�?�,������Q2M����1����L.�L��k%ᄞ��.��u�'評����j�Dxa����)F��Z��.m�f
���G���E���lb��u�O~���r��YG��6�%X������s�Ƈ<A
iM�ēyq�p�YF����y���=���S���T��!��ʠ�ݚ��V������8E��kX1�e�qa�*;?0���ةw!gP�7Q�Y�$��}V�Z��r`�� 
�cs��߻��`<�m�z2�!��⠊��I�8-�~6S �@�Q��`x~䰃-����;c��}�*�����>m���ζc�W�'SN"M�Z�]8�����;3���H�t����{<u_��]��5�U�������T�+Ql�v�L¶U�@iP�ע#��b�dͯ8_|���z.
 L&W�j��t4W�]'R����e�Le��͘N���)����Pi5����}�ܐ�� �$�?7�b�"�rc�?�Ŕxg�Zj9�C�ӌ����w���ab���z8�2L��h��[�$F������:4���!�$8梼����v��xWV�V��tk*Ӛ�J�a&8�DL1�֊����U�AY�xg����kp��a:=���D\��ߤ�G�vk$K
sd�-�g᭘]J�C����ϯ8.��Q=��Bz7#��Ry~V0�&�0b[�A��A7@Q+�*�e��>�Zж
�������rSe'�7�gǸ���T\ʃo8s��C�)q�@�2R{�jp�c�����V��o���5�w�Z S��A�2*�8�Dޔ�ٲŵ㇐�����k��C~?R�u���UZ�f��cg�N����0�6�8�����{ ��r)G�uO��4I��w�`I�@l���u�_�"1k���\FVĕ����N�?@�ȼ��p���� <"|���ľ�(��`�Q�eU�<��=��W�=���k�5��j
��iMGm������b=�Tr�-�T�\��F�f��
����%� �.�x[Qt�L��"�}-�x�#�V YӦZ!��|`�`�~����h�~�� f�DZ+����Q�+n�@���H0ݗvL=�x�<��5�����#k�S"�)2x�i}����"��=�]b���z�6EF9, ek����,��w�/<%�s���^ 
M(z�-�p9P\ ]x]�v��U}��{$�����]���C���'�����)�
�Y��� �[�mju��=�ݶ%�[�.S��W;׭�n�`'�s�zz��B��@'��j�1J/,*0=ª�x���_X��e�3k���+s�3Y�ӊ�}h3�T�o"ow��o��9Nw�I�aMaG�DT5�N�R![������.͞��"'x��fs��u���J���B]��'x��VfÛ�s���V&6�V������>B�h0��Z� nԃ�,mM�i�&_2*ύ���!�1�F(Oytg�ªp�q�Zc�?�0`�ћ���
z�����`�����Ƶ�'=bI20V`)�W���y5���r	Dŕ�3N�6��G@Ai���A�v��b	��Jj���6p�B�	i@��\���W�-���~c��J���KŘ5��f�.����2����oS����-X�H�HaO��K�Y�|?Tɣ��'T֐��1B:�x����S���2�fTM���TB䦯.�:�!�t<��E�گӛ�ݖ`<��pHYV�d�3���ym�}W��G�UO!B�02���HԦF�%R�=��m���N/ꁯ>v~RI*�ķܞ�Xa��z#e�����0�Ѹ�C^^6��Y�S�Z!��������L bZ�۾[pȧQ1�#�K��%��=p\��н+Vo��i��_� ����x��e!��i��7��d������Epl�m��(`��9G0�M_�gJG}L�_t5r�=�>F�蓻������@�B�֙)�g�"QN_�@fJX�����,�������
F�<S�a�>q����1����l�^��(����5|a��ژ��N�t��?]|�ENtU��]ˉXC��:����>2'�Zy�ʣ1�y��k� ^+���w~��+H���*$h�g]~x�~��G�<�[ha+�? �:K�[�h����y���y�Etº�����EZ�yb�K���#,��jzaX�Ss-��B��_��*L��eQ�7]�ݿK.|3(lb���%�]���͸̼������h��07�ӓVI����$7O�2�%�sR<�캲n��ȿR��'"���������BO@�9l�>�wt��gۉ�H �!˶�%3�ݒU�	�FC���9S��h�F�����տ- �����6Stte�ȸ=��-a҇
�^��V���iN��<�4�m(����ƈ�����A�H'�R_�\"N�"+�����2~aM!�E���x>�C�Z��<�ԴSr�J��Aj��&'������~���ٜF��Q�@��2�ㅚ��(m�Ί&�� �=�?����B��d9;�L�4(�i��Yw�Q���T��&ױš���t}fz��ZQ�w��.���L��z�v|;m�α���mᯕC7���Zy���
zy 7N0���^���b�zW��h�����˚�}�)�$���̱jb�����ƀ�o������g(:aB	�䃩�x���Y��*��S�;��s�9�PTb&m�q�b�YB�0?��e�<�PKE��s8Ksw�sJ���J���G#�^���x��5��-���� ��ƿ�~qh�����%d>�l�cXh�"���5<ǈ�<����Y�a���y*�s��}�\'+e�Yk"�H�KUVml�+ܓ��cH�.r-�r#H	�WN�|�_B�B�D�F\,Nx��F����=s�o.���qd|�!����gG.��h��}�����t� ��|�����L?>m�һ�*�ڵ!��Ւ�(y��H~�K�2��F!�2�UM!�">��(_z�f
&��
�	N)�QCrr�4ȻKs��	o8Յ�}�� �I"6p[�+�9��^$aO2��%��Oq��,�{���^�^��-@��:�a��]pL+_څ��k�p�cg�=���u.�(c�ކ���dAR!H>��v�:�p�X Y�5dM�:�:�m(Z��]q�5��������`�F<���&�����Evޫ����s�p$O��#֤�=��MG���k!+~qME�]�ҹ4��T����*}�H� �an:�iډ��)�`Þ��I?!Ƥ�����%xO>|����]���� 9���'��!�p����
4=�Y)�jjvkf5T.}��F;�^������8�̰�b�����YcWm0�� ����Np��>Y.���zϟީ/$yf�7Yr�0�3m���h%H:�'���u����{�6y���&��E�@�Մ&Z��z��u����aO(N,�
��3UC<5]Q�7E�p$nY߱"�N�"���QNr�-v����G) ��~�����G�_�a"�a�,��S��٨������Tǀ�r��CQ4���%m �b�w
ii�th㚇�T���Å�#��K�I<�U��K��w(�������O���̊��k���/�rop�'g�	=�d�^���o{`�)���A6�*�6�f�����@M3uh�P��K�L����O�'%��=Z��X����o����7vW���X�����k.^�*�>�hz��Ϫ=E�����^PpٞY����MN]�V�,+�^+�7��V�"��J2�|����^�Z����R�j�ޢe�
�����$�?����?L��u��'�T1~%�9�&4,����� D��<�mċo=�[���׵�s.�;��&��#`�u�� @J�g���rp��:��]�M[�_�e����כ<��x���]dl�J����/Ws����7�C�?��u�ڪ֫�h��莵�	�Ñ�"�r�L/��x�K���Opr���<8f�5O�߶j���s���8��_�[����9+��
5t�!�r��ߌYT�I��qfT�M��8hD�x,t�ֿ��|4%�y�����U��@B��`O���G�ٲ��B���	}�17G��w��E^�`��a�.�BE�.z"����H@����z�4F �o!���z����
ZS��=�B�`*�����u���v�/OZ��R�������7�����_t6w2�0f�FT�lŒ�bx��u��c�ݥ>y^骄�1@�R:��b#�tYՖ���������Z]����bo>b�|��t����+M�������M7d��AS�:Jx���fg	軚#��Y����C��N�/���]p�K���;2j��SV���ߋ��WZ�#�0�?9'��3���O�DJϑ;����2���>{Q��h�~t���U+�*�*2���Β�!��� r��iJlG�N��K�E�����.�ժ�����k\�q%ڕ�]H����K�*��E,��%�B�U��,������^z9��)H<���(����д�w�+��)4�\�5�3��PZM����Ǵ�@�����§�e������K��kX���f~�#� 	���cyc.�j�޵�`kxCs�ʲ�]�!��V��%��r�l�#�De� S�#я}�� `_Q�-�����dt84⢏��DZad-�o���S0���:ԓsU� y��$�L�9-��K*jHC�;+GH6�0h�5��f�j�T�`G���f�8j��V����񆑠�vv#�B�T�_�.ө���jf�&�w{��68�������ni���4�e7���诨����cѭZ�8�ײ�`�JUY��p?|"��1:�Q��WN���\8$Ȗ���]�9d