��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ����"WYj����i� �N�7A!�@<e�]N��?�jj�����W���a�q���#����MP�F�pdoF.8��+:���h1�ԭL��L��[j�1���߀/AP�0,r�F��x�N��>�RziB�M�\�P�ua��B�MɥBe�U�����v��+�R��|BC�:6u��8�B�����趟���*���I�lklry�.T����b��`A>�7��UzVT�*��"�}m��0�W��wS4ZuxxW/�'n���]�:kڗ;�޸�	��Ү���G�V�m!�������"������ ����J'"a_!��@v"F��z��K������W�Y�����Hw���5��Ip�X���
����1	�,z�蠥	��clYHް�x�N�5��9#��8f�r���~썁��x�ɯ��}��]�˂4�D6�1>@��m�����������@�Vo�n �S��˂���U�+�_H�̄ �����[�6�m?j;�jB'��DT�,ɅzYFw�F�q:7�ľ��5&_2,��j�l��XDr��Wf����0y�Рx �0J�#5!jb�	���B�*��1}c�i5����w�D��M��a	� ��\��V;~��@Az]Ԯ��3vK�%/޶ئ��싾í@x(i��Z��K*;�C�H�	� �Z_,��G.���V"�h왑��1�}��*ɡ�z�F�|9YBJl��������;��������G��(�ɿ@�ٚo�Tt��kBk�e�a�D/ݼU�����,�]���d�[3�H���v���ad�3�츈���/M��ϲ�&��t���AF���9F���R��"I��U|�)�6��]��6�.�~�����a��n���,�S�98U�<߲�y\�9�m�(��ŻW[s��C��-,��A�u��ˡ,��͋����`ĎГ�!4��n�≯8SJA�����}��7��h�o������+��|�0����T� ��.u�m%������BQ��ϓ�G��^�"��n���A����ͧ��1��,���XJ�BO�	)X�/����cz���H(�a��5�}L��;�d~�������{���ǽP�8
��rg���ON��T�����1���=Ĉ���X�1�yZaZ�B�6<Ck74s
�4�ぉ0	z�R�Ɍ��b�4��O5�I����bke8j������7���;!u���x��*���?��ka��mQ�D8ק�%��(�^2H�lS��RM?Ct�<M����9��Ծ�1��N���VUV��T����4)�_�,P��S���Ӂ�0q����U�����[�WU��ٚ*)i_�Qb.S����-�8�&����JE�U�,(���݆ZT���9ҳ,���7L��zt��b��s��"xJs�h�?�0)��!�ߺ��ϰ��㔐PR�f�	_7��2�qB��.����u�wYR#ݨu�>����v���	s[����4�\S_3��<2l�H&-�1Q��_{|�=�`-U	�I?�a`��!��㊩
&���C���F��������4�:@�'��7l��.��㙻�*�'oGS��x���d9�-�2�JR	5�r��0NI�(d�`2��%h�,��
]q�Z	�@�a�d���N�&�j���V�HH����E�c;���[��C�/P܄���;�V����)?�}+f��	���v,�R;�Hػ
b��0����9ԓؗ��������a:e̜�E�INqD��_��x�ѝ�(���U�4��s�#�v�!.�j�Ȁq%��Y�{M�L�\I�oQ^xY��F��)�,q�.�_`�v�+R)�V�Bи����ju�7}��!k8�>X��?]�r�y��P�6��y��
�2h��pm�w6�8i�ӽ��̪-t��Lv,�.$B�w���0�r1+�
+U���K�=߈�_�Vk�G-�`@��V����9W��M�'9�Vw �J�:jS��
0p�⻿8�e�C"��yخM�q�l��:F-��9�lٍ/2Glj���B-�.���C!.de�4!]������٩��0�0��x�T]2��*��~��RI�007��(؜�� �_�ᮛ��n��#���x��e2�O"L���D��מyI�YB��K*C�m�C涸�bE�����4e�T#�J��!-ɋ���p�^`K�R�	{`O� 􄍍�*��$���D�%Z_ʢ�������aG���E֨[�\m�;�IL�'���z�B>���W��.���,�ѱEv��i��iGa�n˩.1*�����Q����8��jgc{5�!�,���o�H�~>Ъ�.f1ot5��G��T����>_W�,��K�`N�Dw��F�,���C8f�V�|aw�.&����FQ�^���:`j�u�R�Ӗ�`�3�ER��˄�wA�E�F�%�X3b�%����e���VE=��8�G� jRJ�\J���#���/V�V���%�w��j-7���S��4SNVb;'68>�H��/t].����X�Yd\��2w��� l�����	�d�#'˨����%M�7�Z3��UP��i�D���I��r^�̺pO�w�,��R�{"bs�C��Rꁘ��!�CCPj��)X�0|��zvY[���j�9J��sĺ9s24�����.j�<
��k���duXpOYV�q�����a�a���p�O�&�c����[3�h'wYC�jhŤ}D�/�O7	8FƲJ
E��9��LK],��ջ�6\����:����}�=��Մ&#ɻ�Y,�J4vp����<~����{����W3�c�u�W�ܯw���a ��H�O�ͭq%�����c'�.PN^��k?�EJDk��(֠���z��w`����L���Я��h%8@�Ƭ�V� ۚ?������(�ea�Q�M&`�J�+]�3N*$x�A�`�K7`��)(x3.U���?ڼ�&0��Z�����^I�O'��H�߲+cKE�1�� \m!��D��dǥZ ��\�.��U�@��������MPʻ?��V����5� �ҳ�!��E{"�۫��E���<�-���;{#VJߺt�=��z��;,떍����z� �� ��=8r�	��r��?�8(h���<.�:��PB���;Ÿ�Z٠V�vZ�Ϡ�����·��2Ku�֝*�oq�Ą[���|�tU�?eYO�+����<#��Ns��Eit��m� ��	�����sH���Ę�y���ډ��uh"M# )8�7�H��!ua�$'�6��@nr�^"��H��
���L�0��.~.#���ۋ�$!���D9
4ۛ>�W�y1��G��G��7���9d)�p�5A?g懦�[���S0{���"�$���yI��d���W���55s�9O��RFSW�g�a#z�X�jUNt�pY3V�:���M&��Smu�ޗ���]Զ�Wm�G+��|�xE�?v�����07c S����g�q�dV���FD�E/���JPǊ0�Z�µ���f�ف�4z'�(G%Ca2xq�X��^n�Q?��ςȁW����3����֫ۛ��οއ�!�qH�'�P�rJ��V�>���pO���~��˥�'�Y%�y�i[���b"�߾��M��uX�=��!T_2Q�x�Ǐۙ�+�#�����2�Y���z��C���GjG�Se<��R�S_���aaW8cE�7��Y�����8p��	|��h���?˯�k�m�*���/��c�W�݃���g�e��	RP�Ľ�1�.y����.'>�)�t����kl ��S�1�1x����.u�K7��Bɽ��?�[�	��:�u�qc��9��z�P.q�R���׌��A���su�	6Oh�;�"7�Xl�Ir)�A��d�����=�\�i$P���ۙ�w�v�O�@EL!��"0����"�֩#��hBM�V�������6-z�f�8��*����_#H�;�����w�i�C�R*`�i��)	p�2g�Bl�t�����߇4ѬG�m�5�2HL��6$�cDxj�Y��Ӑ8���%��p��i�����pu�ȭ{t��PrRk�i�uru^�2&H�%:��6"Ec�2�6I��l�"4	�=)}5����SU�O/]}ݺ�^�:e'��o�Oy���+
�w�
���.��8�����^/�=.�A1XZ�L�&�ޏ���3�DDzpT�F[�����a�]�>آ�+�گ���m��Tn�3WV<�%A�4�
4��/�|��7���<�Ϻ��J@�c�H 
LW~�:�p4Y%
&�/~�&��q�1L������ku�1�b�h	��z�XMg"Q�W��6�u�'��)�CZ�t&	E��; ��4���I��{]e�Y3�|)3�3�KΣD+�M=����`s�jq�����e��혛y��8U�F�n��`�.Z�a��#�2Eҏ��j�H�A����T���ɬ�1c$4*����[:����oa��q�`*;�2 CO��/�q��}��:�r���W����̵�b����=ւX�}�(z$�A2w�����{Nt�Wט�h�J�B|���Խ��vm��5�~Φ`V(��7&į9�,�o <�{i���9t.�3j��9dO�Z��po��Lk��az�|�4�,}�+�Jm� �������0-s�0�VVT�HKP�F��s�{��G�T#l�&����\�bܰ�Z.�IAK��SK�����5`����fe���~�f���,�AͪQ-)�E��6�bY�� ��37�k<HX���o���W��3��b�>�m�8>}c��W@n��Xg?0n ��<v�U�K�$��ü�x(��s�Wӧ�7[��.��#���s�v������U��hY8a��@Bǿ��_O;oY�	%�9q��T�����lW�:!	CJ��q�BӚ'.(�;�ӕ	�'8i�[�=���5��|���c֭���r"2��W�:.�B¢�P�+~^Rf�X�=��A�|��=Tȶܡ�Cܦ���bp^?Vv��Ă����BkULτ0G*��r��b_3}�Q)�<����B���1��CϊٛD���x�#[X�c��Ҏ=y��O��-0
ұo��lX��LN�G	#���~��h9%��klp�"�V�������=I����U�b��3�/�P�1�šn�L�AfV���h� C˹P��f�sE�Lu
H��h���3��G)6�K
�K:���[bU��K��`�A��4����v(�줸(���co��B	���3�FٺA�Ŷ�ن)�,.*\�?XmV���z����ޢX�E�oܸ�T?�7��(����U�Vl��ŷ�f���5�J�j���6_��O��߬h2�؁W�mve?k�W�*��c�I�H�~���h���#��{Kg�W}a������x��e��Iv��t��{رs�X��j p�/uiw��7#'�!r�ӂ,���pG|�
ә��L(E֯���p�/����?����+�v��G��bJX�5@&Z"����������-�~;9۲G��d�z�vP��v+�[���8��#���p�sc�DƋT48P�j}�e%e���- ���P�k�m��S��¿�����N��h:����F�%�SӅb�pG2dXPy�ۋh�D�ԥ�����ո��`#�yj��%-}��)xR=4�~&��M�>�T��.Z�)B�����Oý�Y�\�DD|=d�yz���H:L�P3��?�ñb�����L�*��ڷ�M][ �E_C��U��OiL��aZ[������G��Y�u+�/��Q��|^��zV
��Ũ�g6����74�8Vuu�krNW�R�'����&"�\B*?ד�ri�l�xu[@����pؒ� ��;7�h�����c��� �$2����|-_K-[��1S.�����Z�^�ØgUi�.I�(ꊓ�����s��$Iō��� ��Z�<�$����װ��%��; 
1>�(��M��P�&I����0�yE��/��ژĥV��Ia�+�9��+Ѷ�6�Jމ���3�������j|(i^k�
���Y��U|m��c���N�/�Qw�Y���_|���)"�82�庘��L���l0%ՠ���Ǹz}���P8l�!��ugULD何�4ٮx���(*>{i�t���Z�F�E"��~�y�D_��d˸}�̣�=n#�@X!����m�����֠/����RfV�Q��D��ߧ��u���2O4� �_1hn6(^n�`�Y^�Mn��&��ak*U��� *�tc��.yX�]ΐJb���_��e���X�l�v�hf�6?=�(�)�Zb2f/�co�QT.S�0�E�����}6jz)M��I�~>&�2p�fo�U�>mhSIlmC��A�7|�2qp
vl!Q��7���X���U����6p�Q��`�"R�a�f���%&��D<�q��- ���[��9�~�-��a�g�n��H��.]���r����x��o!��!_������b��D�nus�k�	����O)��$W�Bǈ;���̼�u��wxla�>@*~���� �_3Ws�
�w����{����n`)��)��ALhz�49����m��-�w"�l ��`ǐ㇃��D�mL��������L�^�hx/;8<�v����P���]u�5-}���y�EI���(��kB���H�Dj�Uā�<�}4���{����% �e+<�\.��pJ<�� 3Ҷ=:eP�
J8<�ț����*N�i�ɗ-�Oj��\�B��/�n�εׁ�ĺ�̲MTNf�T�7=����.��������I-���+Q���v\��$��c�� .�֝�ë{ߗ`}?jP�;��4���(�eAO��8���@M��`���-9->u�A`{K��~9����CǦx~~�a[�����[��+�f�0�iA=Ү��kl`��^����mUT;T�:�a�YT��k+����"J��Ib��jW�*9	�$8k�5n�r|E(��� ɂTJ^��R�4&u�5�Hod����X�M�,��ڊ�
,�9�n���,Ĥ��t�� ���Ye	c7�H��c}���u~�A��/��#��S�/���6Da�d<Oi��cX[��`�5[v�$'r>.�5�τ�I��l���I����Ԃ�����j�X�@��'~��b�kd[WƫӵX�G�"��u�"T�e��Uu�:���H�-��M��S�5u#p�hJUa��iP�-�y�[�!{T��e������59 �,v����4��/W�����A��ĽGU����Iv��{�F�4���Ƃ�Be�cU1�Ϳ�a�#�t�xSY*��g�u��׳/Um����"�]�*��:����`���']Z�H۷~<���Sk?��4����NE�9���ԋ<%3�d<�z�oL����C��ݲ�VTw�;�aB@wq%�e%��ӹrCD]��+�D��a��ߝA	x�R���bd�-at��B �{��7� �C�1Y8�	@4
Ş�ܖ�}��+9�^�:=i7�� �-rǘk �Bҷ��2�� 8��u U�U���B>�%��pa��4/�V�}�e��Υ��c,OA������P�{ ɳ�`�v#���VǕ��`{�PSO7��E�U�z}�D�� �`�T���1��9�-���JH~�?N|��g��A��)����_�#Hy>	vְ���s��r�����.kyV�8و�N�7
��l֐v���;��w������"���}��X@N ��1�yj��'��h��3m	5���[�F�S��� ����|��?;׿�=	w��< !b(l�Ha�H1����3C�b��f���A�ę.O��f��t�&�^�﭂#*�^����=a�`��(Q6��!f[�^����2 Au��%k�A���Qef�m5DF��`M�K�G�5R�'=����~��|@|�'����W�&��"STޏ�N�9/�8e�ʨ����!��!^�l��vI~pY��D��]5��o�2j�d��B�w��~�p��=�\�R�y��Ҹ'�'�8h榠�Lr��+`;Os����]�7�0�xzaoKG�5���GT�*�ve��&���C��MD��!�{(m�T�EB]���QP�h[d�|�,�m��Z"I�)�:~�e�:��o�Sm9����ŗ����/����������!7��7sP�v�C��yM'	�䄯ul�Z@�[L~}�=P�!���o�d�_YYV� �� 93W$Ρi���)R�a�-��^��8.�vd�'�5�ew�PG�r`<4�0�%!�l/zM�u��Tț�	]�"$�Oi�u���[ƌ�w�����,�(c����I6-��hm?�U�P�sp�<�կS��V��<��^!�69�i�T�Y`"YH�j�5�A?�_L���`ot~&[i%w
s�����Z���� ڝΕ0�ܖRY���"s���i'����2�M���ó���u-�gb4w���l����72T��:���5���|��`q��z�"708�K�F���-:�>�>W��U�M�� ��]��\���V���s6���92��\EU�7Ӧ���۾jEQ'(��Ցj�=�Y�	t�Y��e�AA�F	2b$_�e6_4��p���������݊mJE�wV���G���]R�݋�H�Y7�!L�n����k�u�I�7����i��9�e�ao��|G�����M��\/�k���vv��"�V���8Ϝ�9�+��Nx���^x��'�Z䙩�5^E=t����7=�ڽ 7�I���:���_���@��);����/T�j�BvZA}x��1B�5J
���OQ�w�l�6���ECe�j��\lt5Z:��FMyp��,V!��!sɰ��I�ϩ����?�$���{���Zꇽ��ߦJ�F��̏J*a~��T�p�5�zɾR@&�<(
�aw�3�U��,B�(M;�U�Jut�C]ݔ��lEj�#+o���K�%pX�{�󪹾DXC��bfj����
)�QB�����"���g
ݸ^���&��Q�P�ҭ~��Q�[H�I�j&B�bAϦ%���Sa�y�v��E�HmL�����`wuY(v�e�'�8^��A�X7.R_�s0��PW��.�lO�;I��G�!��Ia}ڞ�^�'��-��~��lH�Z]��=�H]��f}_�鰡��
����v�ERu�������
2U�Uj&B,�-%����G��)�#/`H,�š�N��e��#�[v��l���mJ��\�ij�¦Y���=_|z���HCAǷ�c3pZqT�c�2��>�ic�#j��v��$���`���&�>t�̗궨�����M�ܵ���� �/��Z?P��% �f���tƤP%�0wc#��a�9��^����a�l�ʅ�+:;�%��ys��2�4[ZT#�w�����w�Z%���v�YhI�N�����[;�T�dج��Z�)�s^�:�fkUb���W�h�i"�2�Q�4�r2ea�+���S=U����%�W�������ͼ�(����M���#\ 7V�X�݃��UES��>�6Haqpz��~v���$�3q�(�^1������j*��)<�1�4���d,�5Sr'Z9O���x/�)�X��R�ܕ��|SMG=r�Xso�� ��\&�D��e�pf�����	��Z�v�VJ�F^R��\�^�/�."�{��8M$ɘ����J�1�2+r}�vSH���g�F\�X� eu�&qnY�����9�Om X����ᒾh*؊%TvU�����Kvl�PM� nK���1u	pi�s�����	�_���j�a�p� ss|5��#	(P�.<���0�}��-��T3�h�ex�K~���*ȉ]�]���f�����^�޸&�p���]���)���H�.A�;����iH��6��e�_��+o���+9Ҡ>$hQ����"~�?ċ�/r��{���!@+��>�s�$��p��w�%�u��?x��D�K�ߺ�j驢�go��)����Z�)���ȹ፻VMi�$��t<hj#���i�1MstΠpnz��s��4�ty��'؉� 9u�����o��1��������htuq�@K���O�[��0ɿ�rxO�m���򈒶���E|a��y����O��aQuc0	�f�a3���r&h���~���"&5�j��偄Y�Е�Y�SyC��vUP���4��:+N+� �lT7�#�He�)�Y�����P�����������o�Ƙnh����� �:��8�"���B�6��#����v/���S���ᔆM��s�[�ۓJ`����_����!�}+���aT�'ˈ$����a�҅�����;�������+0ߞ����SJ���,����q�[�<�o:�7`�Q��Z�X
��!��ggBt����CqY���(IT���}]�E���{@��K�ov�����3�|�˄�i���R=ף����s�� d�$Q��rNi�'j�]g�=\ݪ�I�la��l�&,���Q��OϣS��`���:��:@c��y���A���	�@DaI����4#1B����B�� )w��I&����bw�`��
�O��2k��!S�[jd6 �M�q|#
�ES$�����.2�:����(��B�~0P�+�0RZ,��ƿ��1{ꋦ��}�А��r����__��V=X0�ش`ՙJ���'Ƈ�J�"�������s9���xL�L�{�v��{�rm�<��%���� ��yR5Tv0;���P씛;|ɹZ��8���ٶ�}�p�	�xg�����.�i���l6�*�E��,g�tpv�:���ڲ�Y�_,�YY�u�s-E����"��1�q�]���m����@je��-Rĸ�M�c�h���݉9�OIL�H\�}�G!:��%j��@�6�E �C2���A����K(�����$ˡ��X�S]3�Ħ$�ꩪ�<��Ŧ~�D�M�	}d��A�.n�Պ#O�(��C�4���z�V���	�=r��z���`����x:"8C!Y�� nJ��W�q�1H��ph+��р$Z/�^�@��^4O��I����'�1ڀ��;����w���Iq�~���S}�f�iǀ:�v�U@=�H
+E�]UI�PW]Q�#�"�M6H�h�	6M��+�Z �"��9/��cD"��^{T:辔;3�)��Q�н+��Tz�&��ӊ���p1!4�e��2p]On��h[n-�ϑ�+J�O|�v\3��L�I�B��1�r՜Ut歵���V�����>c�C`��ڕ��}��0͐���J���J`\t�<�`��e#��/dX��YCr�+��-L�P���#K�T3Z�~d�CU����Ky���Y.\��u8��v�9��i]R�oJ���P�Y9���Dh�#%����
-b�)�٥��B�bZ"I�2��U���`�>����2(�u����)l�}/V.o�Ri|��Wz���M���բ8�ă��0q�Q(�=T�i��;��!= amC�y���Q�) ��z�_�Q��ȏ[V��S����� �UVa�����.8<M�BU�V���ݻDR�"Hy�w�9������my/����|�l�$����0�VF*�c�M�bӞЭ�`���J`�V��k����K��-�p��,�<�F@���l�R�*e.u-����lB���g�����$�:��vt-���JRJ�r�Ҳ��(�����·�e9NJ�ɓ���`��͝��y�@�* ���*���wi��#�M��R���y���7�m�p�v(=��7BC@��y	;�ƺ��ǝ�*�+O��!m����1H�&�Pz( c^�'~��D#P֓YZ��Y/rG�����8��.�L�D�*�z�X���lS��;`jO%��]�_+b�Z�.��"®�.k�
,(�[~d�IN<)@��cB����곐��$��;�3�:�oss�^rn�?Q���N�ܢ[����1�*�݊�%NJGOo:q�|2���e騌��dK�6²;Ǿ>�}�\�}k��=0���Y���o�d�x<<�V\��}f������h �~k I��T���bcj�q�PL��@]���ؚ���FI�!�|6�&���?Vy��4E�Ck_��*�g�=�^�]Ux��(������l���$d���']9
� �t9Y5�\�|��aF0�`����>V�+Y��s{/�������6^U�Q=�F	��t" [VG�<0��	@�9���ן~����P�o�܃|�]-�!��4��x��n�|��@hD�G@�Y�e���[��<U��wbE�v9�w�^Q��3N����<c�4����8!�C_'"���.\�_��qM�趷G+��;��C��2�)=/��K���{���n p<���8��������;v��%)Z�q�|���s�S��J����p�W�i�������{sC��\�[�lT|�W)GB�m
6c�($V팶����P����=6�=Ƒ�����ˎI,hm�,s����T�ΰA�0#���(��'�t{:�fqu�� n�̜�(�>h��ך�,C�ө���0OAQ�����	��#G��]D�UQ-8��J�L�h�o��l�!�o�A��E	Q����֨~�P���>#/�'��z/].5��D'?+l�y���Xœ��'q�����Jkd"m+���@�qa�Qg#�#����c��cBߥ˾��6��N�8A.��9|��4�����R�KkL��#Vyo|�������D.�P0�p�8�I?py��9��ǟo��� OH�s�� ��aP�R��<^O�f�	.�����S�'�>x��f9U��\��(������n�$�
�F�C�f��s���-У=�X	ҍ����1��92����#|�+��~v RY��	O:̅e{��E{�ڇg~��i7z[�X�c�vV��]�:vNz_�w�­"�U��\�p��&iwx��&�A������ny��(կ���T�m2��V�aQ%9p{E71?�J��V�7,�@~fm�$��c_��y�{^y�w 2�A˃ �XC��7�Ȇ�vY��1��'Ph �O����45 ���#Gi�ah��͓/��+XC�u�� |�=��Fk�������S��݁�_�J�u.0d��*�n�/E5k3p��3ĂJ����Т62)vB�c�e�#��ue����Ii's���:�Wv���:��݁����W/#r)=Å�?H�A�2*�'�er���u%!*��B��G�Y�r��L�B��<|t��+s8���� 6Y|��Ż�������;۰=��y��~�s�N$X�(�2�-�����l�|��c�#&6��V�5#�K�QLj��j�����`+�ǈ���Ϸ�c�N��qiʜ�&7xy; ��;�0�Jk� 9�-��^���Y����>C\��Vޗ�2�!9&�؍���F�Qí�[�!��&���:|pa�b[�Qtw�d��깛�jiSGO΃S7�D�ޚ׊5^r�g\
j�8���I��&c������#$h&�:����s����j� �{�����E�����M��K2���_Ď�=O���W��K�$MH�YW��E���#���`Ă�	.�WUuj�9�l]e��3�̋l�n"�����SO���~�xݎ���e��c��J>O53҃$?̖V��|Q��6�ｂ陚�`��|\��pP������e�\�~��>=�
Ȅp)��|~��.7s��"p�g&�l����sv$eA�����M�Ҽ�K1eL����^��ُ�({ȋM�bl�^jz�%��E.e���i� � �r1(�t�:6�V�q\,�m��`b7{��]����Hh$]���qN�0��̓�4���<� W˃&vG`��2����&���4�	��gNXg�p�2��y��i�4F� �=��Xh:���^�+} n$�(>0���:����r=�{�!u��7��M�Y��&��Ĉ�I]�uό����=�{g�
��޹u�!�bP�Mz�;�=.b_f{+D�S9}r���V��E:\���2mdXPe�%�t���ᖩ]#+9ZXq�>��Fe<س҆�Qb�����s�
�i?/4�pmE͗�!�Y��ڈՐ�,#�:oz&qhO�ZlE�yB�N�� �L
��` �[�G�:?��$�W���.�W/Q��S^7J��e�~K���T�o�<V�r��	M?r��5�wW�TT�������h�5�v�-Vr��o���B�8��ކE�j���`|������ܗ��	�SB�b}��b&����S
�B�Ō71Y�3�G\kه?�?�����j?�<,����W:$�4�%�M�e� [6�	,o���k���wF��Q���7���*&Z�}W{�$�in���K�זaH�H�`�g}~FMw�/	J(PX˷�NąƂ28�ʊH���Z�5��9|�%	��J<J�\↞��m� LU^� �"nX��}9%Y��X�oU�O����H��� �΍�����_���jΙY���~�^��DCT@ӕ�����-�Ǳ%O�a¿��P~�na�'kW�$��n��VN��*\N�)-hT��4!�3��Q.&4�=�!����3|��t6�*���>c�����-?�ߣ�)�{t�����;��7GGb7��d�ʦ�I�g�CP�p��7���IF�+sP�Ā�Z������t(��:�}W���Ӏ�PF��$x�rO��[�hm�?�f.���{d����� �|����RF�^�UZ�6���([A&f�a�ugnK��X:��E�R���ͮ���}-bi�BQ	+<OK�2�q�1C�	�6�����rՏY�>��ѩ�}��!��>�=qXHv"u^	uٺ��J^ �����)��#|I��JJ�x,3G�T}&��&)`��fTY�=	�'\��*�\�g�a'R9�)��H�QA"b��m�h�G)�v�zV���W������
5��j��!��6�$�i���1�E���8����+�3�AS�*i&���:8�Dc��7���,��uF�{O�e���bw^Vl8s�f�a��IS���=� >��/R�Pڈ͸�nr_�n�H��9�h������-�\��`�&si'c�)G����#����;4��Z``�%���Vڱ�^$}
C,�BLs
�\L���T���_K'c��х�vd�*s'?�*�<�n�|BU����Y�4����6�H�e|-�т5�rEP�8K�jضU����D���
k��*�b�V&q�d�T������<6�Ɓ�l�x���7,
@�m��_$/��Q`N�F�e3ذ0X�9+��3��)||X𚝳�/�oD��2�:Ti*�:H�s�),�#����޾����L@�k��*D���%f�<�Fe� �M�#}�ɵ6�ae9�_��E/�]]U-�Ӎ����=ۆaƤ&2��M����l���WlVNБ�,�.�^i9HK�SAsP�9J����St�*�R��o����(����!�6L���(��e3�j��B��tf1:*�T�Kt��pm+&l�C��B�����u3��cr�&ǽ�45�E�"�tI�°�zuT�����6�g�l�����$��^����ɱ��Lox�P]Tlu��������o�&�"�>Z0������}ex�Rza�]�R�؉�
PO K-��;7-%�2��!�7؊��@o5�����?���*���S �X*��U�k�M��u�ǣb������Hm@���f�ͥ�6l;�i��;����������@]�ya�Y��r'�	˺�ST�e���j,��A���ކJ��:i�D�i��Rq��T��k/=\>�CZ^C� %�_��e@��`5�u]1��>��6� ���_V-�/��p���������Dm��Is�����X3"Z�*y҄��W�� �e_W�@���������1c�Є��H*o8�<��px���h�Y��\�'"�] 9���XA����`�_x�Ų������2�'~g&���$m|�{ә�4"qi�qվ%Y�,��[޲�d����f_�h�Wg0�N��81�2C3Maj��ޜ�k���6^�]���RZ����Q�߸�˥9g��n<��Ɇ^׫�'h��ȵ
7����g������O�X/'����C;X���+E��br�V��gTt�X�)����>����Z,/x��=l��]GF�*�vNG{���	Xʾdg^�{��0kõ�m�؃��C�"�[��*�{�9����Q�.��d!������9�x�"��m< 3�[B)M���	�+�؟�0_����Io�Z�1��;�3Q%7���
��Z�<r�2�P���5s�!�b�ǁM��(m�w|�)6���1t���%���w3D��ܽ罡$��g!�jg�{=�p�W ���G�����ړm}h2Xޤ��悦q��&�"�(*[~�["L�J�y8���2�nψX�
ablK�SI��`O!�fsi����f��	z�1��a�����k��	E���	��3�]| �O�&Kc�'�m)�� ��������DV��x7�k{J��r,4��E{�7�����tzu��\��2K
^3xT����8�՚q$ ��W̲���魣fn�@˛�ِZ����.0J�f�!��~���i�q��,�+lnr|��]�1%sE;Å��r�������C�k����+�x�K���UQ9ƴ6e��u�p{���ڗ���x� ���J��D:�}<�}͕�,VI}�աv0Z�y@4��L��>��q��l�<"6Sս����l͎DyNק�>x���_(���Q�]�~���1�z��;l���v����K�Y_MW����g��.{(BR*��ddw<�>�Ӽ�v�O+d�Π�|tH6}!��nQ�q�yH�G��.ο�u��,�O���˒��]���������ؿZӞo�Zb�59C��n�u���`�Tk�@B �_�}u����U{�>�Y�=�?�n�Z'*P�9@�M&w���wv��K�p�����>;���z���q`��6�\YjL�&�l|Sm�x�zu�4ǡj�дa{�K�qVa��.���t�g�\f�����Ls�t*#����p��cw���yH�ĩ��#�!���dB�P,=�����a&�y�>W�gN��(��(L� j�=_����6x������G�GC<&���5[�d�� �l};/s89��S����\`]p��!�I*�G��.7��0y�TO�0�>��ƛ��i���0궕
�/��1Q=9��ճ�t��� �]/^�b�^����3���̋Or�î���^qNNOg.� �~Ў��7TH��6�}�U�}޹́�{�b���]���>����`Pm���-$�6p�S�13�3��e��: ��a�����|��Dgs��\A�O5�Bՙc�Fg�J�hp�,�l'����8^̦����_���E��t���Q�¤��d�^�0�eU��6�ۇf�b�
{�:�b}<����=�Z��Y��ۂg�	[u���i�2+1���S�'Q�]/��m����6"��yL!A.A���1}�R�]b{��G�=�`��c�g�e}=��(ێ��z=7�������=>^�oɠ��%kvFʿ���9�h��6!��W��$�7��jF�A-Ϩ篻[Ӧ�9d-O6��>��r���x�����}L����:��с��>�1U���[��CME�Y�2�D��h�:��,$'VS;E�u}�X�m�����l~Vfk#����ˋ��9�ݥ<�Y����!��|���P��{�A]�؉��ц���K�8.���L�^�ةAJ �ٛ�Ɨ��M(������u�ެU|�Jh��ft櫄;�[TwKm�E�����ѥ�1��쑵~�} �f�
8�-�-�D7W�lӻ� H�7��S�w�?�T:��@�r]�8%Zf� �*�Ϳv�>�����|��Q���j�m��)�Ám�
��2F�1��ŏ.#x�y��W*�T��wO��Ib�3��@IC�;��cme�τ�eΉ*{J�������:�������|S6����	���lX�#���N�ʈß�U�9j��TE@�E�rS	(�H�2���%;+�=̃�d���q�bc\�j`�ǰ������?���Q=L�fx,���kD�/�k�暜��x�=і��@P��s��z�M]��9�����م�V[߱`/��>�I���%v����(��%:�3�mp�b��1hF�}ĄN��C{�T������#���3�3��a��/�
�QoE�tr�a#�-�$�m8]F��W�[X;�'Lpf�CE'�XA��	��z�U{~tX��6�D0�8q�o(��dP�����lUT�1�%�zkr���NL���[�/��&4`*��s�ՒX�.�{���3�����q�2���q;�k5BFl���+�wL���[�����eG��R�1.�-Ysz��		R����5�7���/7�S��g���!�^�`�9k�L-P�'8	��\Gz�,����F�Z>\����DqU:N�O�1�8Q^�Ux$�p�#�F�A`�aj����5&g��!!9ֳO�V?3� �l,8<y�[���q���Y~k< ?�#P"�-��7�φ�R�͠����2m���v��D���j>P�2|AV�����X�	]p���6�ݞ��@4��I"�dg�T��X_��YC���n�<�*�uI�7;�~^xfEk�KbRK�ma�`2��֠#�;�of	ʐ赶*����@ژ�����s-�{��q����u��Q,�ŷ�Ծ�
e�Hqv�@�H�,��?g�׷G�d����ZV�i$R �Q�{��ǃҒ�	��93,����Bm�헢hځJ���&Z�#�������F��u��^#�T�vDE�<;Zƿ�Ose~9g<�ќ�x���FD/g��Z#p��A�{������_K�p�gyj7
�T���n^k�'0��1���ݦ6�f/>�u�Br[��0bɔp�2��[���|T� ���ڥ��7w���s9����OhI&m����x�4y3U����ܨ����7�yRd�R3W�pw�����fC2S?�/���kM�f<� �UWTiW�8t.�ȯv�X)�CC<�����8�jMS/ͱ�������2��U�1��8�yQ���S�]F��h�#����jo$���Q����
��쀬�\�k�-2�43�3���_ �V���9��հ��)G{�Co�<׳�A�$�$����*�p��%s�_3���A<�g3*P%S����zx���.�������ޑ�z��xj�_�Q7lC��u�27���]��a�4>σ!CH	�	�%�ra�,;��O�a�nHt�PC=СALψRb��H�V���;vvI DR� t;C�Gm�Aj�s�u��߆���	�2�f�����Ƌ�)H���p!1���K��+P�R~8�~W����¯��Cte�/�H��7)k��N�	�ʥ�����{���*\��I���IW8f`�,% �쟂r1`�� �}�¿����z�漁�*a���(۵������y�ߘR����!��z�s8�4�"�t	i��?��Gu{~����:��P�"%��͜yO��m��bd���QrY�B-J{�k7�5I�k�l1� ;G�O���)���ܚ��X��L���@�;��Y�vR�s����L�gk�e&
��h��7��Dꬎ{�߂��n=�O���:�����CX�6u�Sn]���v��!��%�y��6������p.!�=��/Ϸ�"w�i����CT%�%0����L3=�@��!N.��Hwx_=�E��d���)5��n�df0�TŹS�A���U6C8�7C;�: ��:�{� <_M.� gz����Z�S.2g�f��� ���ZE��\�U�-/9F���n��������X%r�7�6eH�7��q����p�Yi�ح��s���pI��b+��:A~؄}8���2����2�w�x���l?�5�b�0��}f��~�0+�u���t�i^��Ak�������h'��ޔhB���ly�����#�z����	iV�-�%��?@r�#� 9�*n �R�*�x��^ %-8���V��z�U�CF��ڿ7 �$Eq�PT��2O��^�K�1dR3裇c���ѯ��=��U#�B9k�A�rǡk��e �UR��hݏ�88L:�K�p�0͠c�9H��2�&ੜ�C3v��ʕf�%�F�L"$ߥDeY6�S�	��_�"!á���u��.��-�g��z����a�8N���._\�~@|lK�t͙W�z9ξ��Oj�0c�0gy�iԊEkY�l��@3=F���.Q�������]�� �~�/��/�Hj�<t�E��Bܲ�Cx�8���o��7dLLJ���JC�����мkB�#	z�y3�F?#~�IV���c��=�4���(S�iG��-CjjHk�������/[�BH=z'U����_�H�6�;���>�-SƋ���ro��Yge�7LɊO3z�yP��꓉pcK����+�n�"/�����8�R�0�s"����a�f��I4>�0A���<�VN;�ڢ}�w�\9l;os�ݞDX����Pދ�E@�1� 禶)�BU�l�|���k�hU$8D��m,�%�Л�X2�L��ao^������.<L1�AL�e���GՇ��(w5=�G9���h�@j
�\'�i�y�bʻc�9;ZL��z|��'X�%��`,RnT��c�e�7}�����4/U4K%d���Hꍉ?I4 �@HK� �A���"�6L�)s�G�J��j)�&�vAcg��
���c=89�R��~�/�l_5nL��H��(��cd�,��^��c4ђm����������'O����rim�6��?���U��6������[�\ޝ�`�<�O2,�O������1-�`?\��݊��4_.!n���� *'����j���/�T�A=����\J��qgZ��>q��sB?�%�=�㚹��h��ݺ��uf�s2\#��D:5
@`.���0��H�2߅5-���ێ���<M��Q4Z��,vRC|2�6_����>G^i�ν'�{I���W{װ^#�p�`x��V�5����(	��qm=#+D?���[�;�
��|5�_�-�߹1�b��C�0*�vܱ�[�#���1�He
���&7�[�P��wJ�,���f�N��\��.�X���p�=g|S�h}��|O�c�,� ��@f�z_�~MK2r������]���Q��Tb��q���a���z�P�īM����~�% 0}�y;_�0-���WK)�O�$o�h5���>�X�UW�z��=~�\��^�K��4������qٍ���=���j�v�/����_�2lS.�*�^לxh��l����t��3�E� жآN] kvr�Y�n:|gE���1Ҙ��8�S���uҋ���b��׼�U��߆囏��%}�${=ژ	^�E���[JC�ۭ!��'�"�b;�������Kt�޽�إ�]��������K�(*蚖�O2*8f�[�x���Bvp� ����i��8���-d,WIn���'8���4M�Qa.&�m7�����n�)�Lo&_F�Y�;ߧ�����I8����y� �Q��+m�[��qZ�Xyu��9��Jγ���]B��Ɲ�V��ii���T[�ވ���>�$R��r�H�hO6eI1�!ѻm���� z�������Ū&r��VS���a�&�.ivF!S7�rӃ��ѷe_�/,��kZv;>ziʣW�`����3;֟�H�t.=A��2��'o(����,{^�k�9d�Fz�����"�F6�br#&0�>3��8ή������Gm�ZM�S��s��C��_�ӑyrӨk/��N��זt͵��XA���}�I������`���_���T��ؙ��oר�Q�3��X�K�E�g����0�R\Y�Nt���)ѕC�$/>v���L7%Yf��l��W��F)_��qQ����&r���/_���1�%�ȁ�7�!'��s's	�|�Fp-׆�'
v�'��:/n]����� ���f�Z��G�:�(��0Wگ�K�X�Cyct�/W��+�6~�rE���Z�I��I
��Bb�k`���;����፬ݔ��j�QiiD%��^�p$�.��5v�Z5�9y��wBK=&��А"�UE���:��k���HzV�9�o���X��.
6��bpMI�����♿#��t�`S������R�L�n��HŠ�o��na�,@r�
·�!{[�%+*��/�����a��h����\@/�wt f��c�Wnhj�[ce�Q�ѡQ�#������+	!�;�<�u�+i�\c�	00�}�4<��<&����H�X�'F#lYܾc��-�p$}�] ����é�a�P��@�k@��o-��/:��t"�{X���p.v�r��r��/��4h��v9��u�!d*���f���ϵ�8~�(2�
a��*��Չ�M�1O�Z�/�rn�%���[�ܮ���
��Łm��HA��n��k���d��<�_��Q� L�����/֌��($��(+�[I���QC8e ��Q]���O��??K��8V8�>������r��k��0Ҝ�Qvq��Դr1C��k�^\�y��$�A��	���c�DI� �e�=_�	sK�t����]-w|�m�2�XJ(�r�5C�4B�$����B~��/Y.�����$~~w�
�\YM��R����S���=��r�]��#"�qc옣uK�����RMyn�ړi�d�Q�?����$�eU�n�d
���z�mnB���/��!jHbꁫn�)Rqk~��ie���Z37��LF�3
��O�*��[��/n�"��ح�p��u��p`Á3�R�4�ܠ2�AA���\^3��T������i��0b����,Sh��ssx��~R$:� ���c6u6��������r�*�٢xS�O��F��-�r�.:�}]L�G���KOe�y��
_$Y���b盳��Gi:�~N�z�:�Z�+2�Jг���{V��G��=4@
aR�\c��f~�VQ̨h�oM�q��"tާ|�	#�� ���%���E�:�Q\�1F�oǟ?_��j�+u�_��|AXܲ�H�ε��>5��������f��f�|ŵ�n~�$�W�m񏤕kM�km`�m>pFz�M~@8�����u԰ڔ۫��h�"��P�_�X'E*���5zR���h�,)�.���g���ùaQh,ذ�L�Ky�5|�����(*	%_G��R�/4�<8S�d5���I��>���g�P���~��"�"���Ǜ$�'z��(_=fs�lH�S���H�-"�O�O�����a4E�AD3��W<�]�ff ����ok�&�L$�x��o�����+0��z��_M�`T���F����9�ym�vm0�%�j$����cG�r�C,��%�g��h��s,R��u�h~�84a1�F��h���]X��k��X�U>2O�U����:ުH�I��b�9��G���u���:��MfX
B��-��l���3�ѯ7�G����Y!�laL)-A�A����f�I��i=����O��9��f�x�6L���K����V�����.��pr�}��_4�	���5�f������|]y�<�4qf��pv/P`��,�e��&J�[~}���k�xH�*�JE��_��&F߮]������|�Z2�Ǧ)J�]��Ϭ��'�֢&��dc�:-��v�_Q����x
�n:��R���wD��}��r�v�9K�P���=ٳœ���P��tH2Ϧ��L�O�D�/��
��%�d����Q����|4�L�y���8�F��'Y�����''��5bk�C+���W�~����2�#�,�E����ڈا�'2�;��`EE���Hٗ�M���@�B��3I��]S���H���񪷹{�ҩ����lQ�$��N��ps��?ⷽ�?h���|����{�H��H�e_�3�r�_hxEq����j�v[���!�%;�U�H��I�����$��(�^G��EG$�#p��(4�I�b����G��Q�
�KwE�L��~�_�H�%��Ҏ[���!���f.�LT��!H�B�	7^����B�`ûb�V�*?f��|�u:u/<J�����(xv�
�,�k\���,��s
�[4)�ʑ�d�����$���i:�$G\���v[���ǒ	a[����^Z1���4�� ��P"v�j��o��Byץo�JO���>���J�B�	{��7\,��� ��ŢȥNV��ir..`>���������b ��+?�%��?V�����>�x��լ�������~��t�̵����Z�f���|!��Y�f�?l� Jr��	}>6/Yp�Ω'J�E�%�yi�[Z5~	oMB���
?�źjV��Ca��t�s:MӦ햌�����p�ṑ��x�\�r!���%R���	XdOe��(�Evա����7oiO=E�.��zD֗f�
��O�,��E9d$@�Mo^	%*D76�	�{��zE��P�e (��9si^�M}�檎P������߂v�C����n@`�:W�� o�B�yvc�n�i.�g�fT��{�?�D��Dpx���KV?����?�ξ�Ͽ�Al@A��ɦ����W�/Ux���)��>J�X7Yy��^`Tb̉ �,i��؍�μ�� ����w����mM�nM����'���<x���f]x�v��$��8z%<�	������@u��#�x˨є<���	�Z�Fmr{v��s�u��qB�U��ⵈ�-�ݥG����c9^�k�!�ia~[��7l���k�>�H���v^�o��W����/��=��?�ΰ���[T�T����`[RTw^@��Ԓ2����7���b���!��6ޏ�I�$9����mN P�̖3���^h��~#�dü�̂���v1�No���4��naB'�p��=�0C�	��!�q9�2惿t�+ۇ�Ϸ�l]#�#��r��f���ݪA !�6p1�Yrp=�NzU�(��O�kF�X�Dc0#��f�e�Zg�ѡ�Y���gޗX�Lf����S����gM��TK��`;W��=r@�q��R!�|M}��#���J)��wf~(��������hk�v�+{n�0�_/\�!�|�U_4��ɟ�V�S��A�7A؅)��:�ͼ)qE��a9��>o��K�M�K�3r�j>��W��Q�6_|��6�_)���ʏ�^"�[ʃ4ܹvױ|�}SV�krQ�k|���tz���k� #�aVA7����1M�����~��)n���L��ӟ9� T.7�c(Y1xr*�ɣ�1[�t�} �K�b���*����?}�e]{6���,�u�]l����y�W	��Me�}�s�Ś�����V�΃�'a���q���_R��*C��@�w�Y��v��8���7������6�A��$$�g�%�mum0Z�����c�~���Y�Ƕ����F�D���θ/�A�l��<X���a��'[o�/|�z=�"M�@�ҕ�s�v����s��4kFH����k="�"�����m�c;��PV�4̽P�N��'�doՃ����^�[ v~���G58?t��7"��LC��PɌ�U�yu@�cS��+X�%�-z~l�u�:2;DxF��5��u(K^g����m����J�U��[k�^6of�����>|>-f-�*�|��ϔ0a�#���d�C�!���ٳ������"<|�ᇳ��b�a���ꭨ���:�4���*�8r;{Kw�%�aF�l�K��$Z�U?�Ӎ7j8��U7M1�&�~����~��B�e��ͨ�8�]u�/�9��TNy�o�R�4IܚXm�w��m��<vbw��.�9��#�����ҰF��w�n�$�+�\�%��|��3��nd�C��n�����h�{ٲ-�cG�gJ[�p8
,=���1-L��C��9[P�I�U�#���u�?�\ż*��,Bgr�p(4L�@�F9�,j�?o3�}*eJm�����J�]@��J:.�e\i����Wu�;�VSz��t��5H�6n�_@&r��ɻ�z�Y�CDI�1�~W_�ƌ2BD����� ��	T��o�\�[[�kN�W������!Ytȯ���(���,�������n�qԍm�+pfTK�5�u�-a��+����2_����	�KS��8�0"���	S�Q�~�M��ؔ�|�hgD��� �!m��n��{=�x��C�F̊��z7E5cD�O�m��I������NU�g{P�Ⱥ��>�0b*x��Sz��j:�9;V@��Ͼ5낌�@�����!#���U����a��֬0)���93~F�:�9J���[,1�\�+�ϧ�)M� �����+����7�EI�D5"�Z�w�t�xx��xc�7�#"����MW�h_ �w8}��H��tri�z�r1Nh�jD��1�2�UR�d�J�#��>�#D|�e�l}?�\%����BZ��ߦZA��*�&�Q���)��׸)T0�BHO,����%Lv�=aK"�X!�&:�ص3rtf�?բ]�9a{�#KSJO8x������\�F>u�+��M��Do� ���ǡqA�
(�8z�:4��c7�EN�Գ���t����X|�
I�X�������,rl����"��=��@��Q�@:O?�+%$]G�|��?OG?��JZ�9W,���y��V:���2�`.�V����r��`�2Hʀ@�{�_��k��E������!A	oCQ�F-�e;�%�Z��V|Z�=+��kEꞛ[կ?~�f�ʨR�w53�����-�_�S�;J��m�@D:�0Q�G`i��h�}�؁�ر���X���ecw(PJ��a
�FQ0����RgX2Qz����.�X�T�{�䦖�q1��j�q�&a6�~LW���(h��(G��������6as��O��C��g��(�׺��\jj�����l�l?�i�s9���y����H�A�t��0��/���Q}��k�n�
�@�c�5)�h<��BZ��Sc	�WW��=
��5s{P��0eӡ��=Ժ��G�Pk(ɧ���!#f�7K�a�ѼB���>G�gPk���2�K _�����~�;$q+ikw�dQ��;	�ɴ���	\n%v�f7�� �8�q����ym7$qy.ڌ���$=�{���xNj�`=�?ى�_�J�����lÿ���]8�9��9|�܅+k|�]%R�Va�i�k�Y�)CTG�
���8mǠ��П����sB�.�0l��1p�|�)?����B!a,��CO�K�r}d,27� {��/|7�go��t�\֡����x�z�:!b'��*����2.��v6P�+]�7��A�� ��BVc�LRA�������|� os-�[ �v��՟9�\Yu��ݔ��ѿ��נ�Gf��%��!"���;Lvg��60E3[��g�p����x�+tPm���!�t� bt�5����Y���/�L;L�J���a'0�1�/��,|���b���([G���R����9=5����ח�H�b�e��6�\[��7~��X�g��zB6GI���q�:��y���it?���ҟ�諞Ｉc����v�Nx�.2ޟZ'e��a���8C������5��G	�8Y~Ҫ���K��Sf�-�G�
;FFtHۏ�L��G�N�e��Ӂ{�
!RԸ�I ���ș�t��i�5mL�����?�<*s�a!�_�I��Մf��]&D�i��*��;k�]xo\��:^����ܼ��</��U��or�$S$�zJ-���Us���<�<v��a�`S�o��[x'{�T3-��g�fŐ�2.�(&�&��,a�>*�m&�vۊ����j]���c,��zD"�M��4_G^����T�<i�u�ޜ�S��]�G�Vb��SW�`�@|���6ApDwW�d�ř�Ƶ��ˁ� 4��,�x��B��`�n�5Kp�\� �0;����P\u�Kj,W����f$ Q?������b�vjZxi������F��/�;���N=�L�o*��