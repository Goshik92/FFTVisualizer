��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�T0������[&1hX�O�.� ��$�u��Ծ�pH�Am�2���}"iBrNC�l���R8�9mg�Z���e] ��^�+��p�D{��I�v���n���^8&ީ���&����	�&5�nV��V�Et4�>Y/�|:��<R�����_�D�L㨷�;�F�����W !)qZW�7��w�5���N{c� �N¢�kt�O+�!�	���W�͠rV���e_�+�WUiJR���7=�[U���݃o��)�'�/�d6,�?_s�=YB��k���&͈��:��6C#çsMP���H�HÄ���|���̀�G Bؠ1Ǜ;�U�V�Xʟ�=z�� Г���J�os��NY��;=�Y���+ߗΩ�\��| �!k%�]|���DՉ���1�Әs��j`�d���2��.;���jT�9��3���������P{ �-c/�u8�+\��(��)��]�̜�dJ����햯����ډ���xj��]��r��U8'�vD����/F��/�FSu;C�����Z������u&<��z���h���T~�+�٤'��$[��'�S7u52̞��oO͜@9$��*Ͳ`� ˆ;�So3�$zm�!�;�; ��M��uF���/��Xb�����f韹>�~-f�z.0�d�0Pqg�|�jE�m�IgO���ax�n�u�ǁ�SIei�I��5�n�9�:D4ۮD�ɮݤj��ǣ�l��?���+����+�t�30�6����3�[]����M/^��c.���P����Y��y콚���m�-T%Xn��p��`��=��n( ^��#8~�}ψq�P^����%�r���_�a�\�L�?��:��˼�� �KK�ۻ�]���~��+`��N�lh)��^˝�k�,X�g	is0��#g�氶n�>0E���|�K��$1k}��s+�mR������ZVF�;��AH7�6[��h&Ԙ��|��Ji��r|T4R;F�%7}��2��݃��	D��i��-��RN���')��MV��2�K|���t��f�\�5=*�OI�B���I������\��x)欍{������S$�F�t���m�����$���<5��k����<���`H��T�7�cR�O���.�c��'�]R-��^��t����[����3���|����<j����<8��Ե��L���7�(�n��^]��fہŜ�Z�Ld8r��۟�&���1Y�7��uh��g�A��l0�?e��
�PO��IF�[��b)B�Б���&�%e���&�>��2�Ey�O%�m���������Z�WE����e�
�?L��	�|~%)&�MZ���z����+������S[����[�,����*��0(Q�de��#��(g�������@�-�p���&7a.�CE�a?�%������W��>
	p���F��!~2�/�lDs��ԋw�!���G��P�d�{��n�C��}��y6P����u'O��x�0��`FR�AGO��*z��5�7@+u��ky��ʼ}�������@�Vtǜ߹�3��/��ҿ{ŗ���	���;^&����1�'tN�Â�/�󀸆P%��g��*��3	�T�މ�~iR�o��8�S�����-�g��3D�Ʉ1d6ʻ�Ž憦������M���鴎Z@jS�B��[�n�ɌJR���$ŧ*Dݠ��-��l��^G�K��\=�/XE�O.0����Q��gh3�+BV~6Ia1�u�W�@b�U�=
C�p4�Iԡ�0���"%�QT�Ԭ��ʣ�%Ҭ���x\I��%�ـd��|~4�w��3�5�]BK�$#SY�i[�)��j*e�1ՕzouO�����ȡ�]Ϲ��v��xe=��bx�<z1�'��n?WTG]� ���Yi�	$F5��h�[������
�ԌEyY@1��(�I4X	�;��k8���{�<�kI��e
�~L5�^1�R�/{H�M�zB0��fWǒ��C��y[�5���l�Էf;�).�-J��� ��M�|���߽I�d_4	R���<�A=��r�+h�h���dcR��ӒT��<Iq��{�_u��;�~�nJ\�*���ҖzI~��趛��x�
�?GM�����FO�~6�*��*����=����Y���ί��\}�eJ��d�)"1�Y��VE)�	/J���AcC�m�b���-/֥�ﮣ�짌��H��i#�Q~;����>lp����F�J���I�ƿ�)�
�؁G�-���{�M��>Y|-\�C��,�V��rm=�� �;��Xΰ_��:�	�֧~ى�	���CZo`�#j`ܺ���6�	3dO�G<��O(@ϖ�5�@5�z/�#֚D xZ�h
2�-�A�laE�oSe�]��~��U��@�I�����U3ނl�2��a�����W�{Z#.e�G"��đ�.��ꅶ��i��;3�%x@xfh+'}���ﾇj�\_�攆���v���Y�Cҗ͸8�s��g��s�;���_��b�twp��E���,!\�Ѧ��1�gt�86JK��(� �3��ʇ/}X�8��zP��Ṋ��I��C���ʅ�"D�J_2�LI�zF�P]pеd�����5���Ԟ�ֹ���:��z�^������{�I���r����=Rx&�vA^W��K�L�\E� ^���^;��#C2,I����) �m�Z�#0tn�3���%A	��2��4pY��W�<���%�H���l��t��F�^ږC�SX
�$�����[���e��C<�u�	�شm'Ch��W&�l�d�o\Փ�$PFm��<�h�,T�'�%n+2�X�Z�7�l��-�5�S�P�����e<+���y�|g���H9,U�(/�@CRr��=0���݉aC$����g���-�,��T�o�	)���`��"/f+:yN#^�5��5��0\�/�x�ѯ[�Ǧ+?9l}�U.;��� �|�g�=�'��=���1Bc�ʭ�f(��)�S ñiŝ���l� �2)�I`.�[����@��#}Uvt�,5�e��[�5�$ q �|��e�L-��;�.Q�u>*	�혴�I�ڭ�io�F���;�´�w�!������س��Q�pP'�T*-7Ħ�.>�d�d�+?��"U���_k3��Q��/������K�sc���Ӡ��~��2f�;���i�Ī�ЂT��_A;6.WB�7�B�4ɧ6`�y���a��El��̰�3��J�g/��_-�?���|�MX�2/�OCT�;�AA�ӻU��-��{��"ٽ2�~��Zrg� ߙd�����b)�t�3I^QZ�V!��� ��,E���H�oKRǞS�Y�/��;b�ic�'-����S�R�z��(m�!^ �?��b�|3�3�
�Ҏ/,\�i�T��\��9�����s�C:\̣ә��;��&�n��l-�TO��"EiW�|��C̖�a5r��L��k�9iɼ-t�����o�w���Ҙ8�
dh0iMQ6�ڣ/����Kn!^�P�ro���[v�&m��j��4�oZ��[=`xG���<�wSO�V)�xc3ڏ�����wi�Ah���U"7n�՞��L�IT����*��sC����������	{J!*�M}����*ŷP�= �[���7���R�ۧQ�-W�M�2bF��%ʳ.OyB�53<x`F���#V��}���*z�qΊ}�I�gDF� �@I?��ʕQ&g�U~r[�k��tW�Ǌ�N���5|l�T��y���R���i�i��l�h:�{�q����dq?Ml��k��>���w�7�� c�o��Jkv�K3,��$)�����b��%��[��>�={Y����0�R
U�d��7}#��0���x�^�K�d��+-���cO��ż��xnڻ��[�RT7�(��57�o0n���*޶9�! �k�5NuY���Ӽ�1�`{Ao�K�7�4m;J,�C�o�eLa9����u2��f�3��1i�P<5��|l_)�ߨ�A����	���#a4�0����q(rj�њ�u5�L[=���}�ŉWs�	��8>k,�Q�g�r��J`�D��Ah�;�����&�9���,�Vd_ٌ-�/��	����vW�0t,������H���� �o=�V�=.ŋ�K�����H�T��[����֑
���ʻR��H)S��B�&@�a�<pܣ�Æ@����A��@��ls�V�)=9{�%���`"��Yb �rC�g���(�C��tvs�r��j��q�|g9��i�"�7ę]�[��h�yR����8�s>[�*���;�U����\�)x7ټ|
�R�lh�t=����ޕp�B�濨%uHt+����QlN�����w�|�������qb�ʗp���� �VP_H!UDk��<K���<i��>C�TU-n{#�ycE�ʲ,躟Ŕ��lo`	����>����j�]f��)�Oh��r^{*�-�oz�.R +|�_n� A���]�x.�S�f�Y�g��8��5�Ա�9�~0߆�Zh���>1�Z_�*/3�,c���Fݿ�����裩r�S��rq��������l,^��h��H���4�{�`�y��'	�X]�r-���{����|k��REvv�㏪��*��p�Č�� �6F����+��ѕn��s��W���k���H�UT�\��'����J����'��z�a��c\�o_����؁�rf.�･��ҭxS�^���l��K���*ή�#�\�vb��C�.�6���a]��`M_���}� �PD�t-pJ�Ɗ<J�nZE�+��mƯ_A��p�I?ͭb�z� ���5�t�mz��X(�����{��_lZ���j<x'����B.� _a��#���!��r��Ͽ����S�p��E�W����>8߄�wf�o#ҷ�ⱡAw���l�0Z*M�hd-�<�v��Ŝ;��C����!��hQ��tw�$5W�[��͙�4��k��}��	C��H�X$�Y�"1��� ���� ��e�`��;/�)�ޘ�[G��]���f��}��ȅ�8k�-����N�Sm4�����U:b�zR`��J�יwoD�����r��bd]�'Z����5�\M�-���ݙT��q��$��,�2���E�[��Æψ[RPTO�rw~AvRT�lʋ3��5�lv���6��	�r�\�}fdd�媺L�[2�Gཙ枿�JQ�f�2?zmd���z��1p�=�['S����8��,g�l;b�)�P�G�XޭA��W�qp��&}����F�8/��e�RP"= �)�8�؁Q�p�g�KhY����Z���%�i#�����8�r���&��������32vTSw!�^�vREj+ ��9��Qu\`�.^c�p:��?N�ْ���\+v�$�M�s�`4�?%e�d�/#���W���F��w��@B����|�j�s�SG.�9�`�dP�� ���'�qTp,,�L�b(b݌��d��ڒ��M�|��V���cr��ݖ�A,�#�wo/��Zw0�]6r���,dJ�r�.Mqo��QTI;�:��l��s�+Lb,�Q��+���d��� (�K
h^FGQ�;)��� mJ��;����d=��)�*�AD¥!�\��}��a?-�Ug�T�o��������F���~u�������r=	Dy�]���*h�eMa�;z@�_���Ѽ�q��:b'(D&�84�Ⲣs�q�/�6yW���GÿD�&è3���ѣ�L�e���F&�.#U�~�+�睹� �)�!��~fX�XO���C��yz����f;�o.T�Nv�4}&��ƢQY��=��x���?�!�W����#]�\a$̳
���?sҶ{��@�ݓ[uLY��n�]�ޜ�YN9�41ȲzO���RX��a�D��Gr9w 4�^�Zp�I�5�T�U�q֧�ֻÝ�"�V��r�/ F���j�iG��f���U��?���qc�h�ql$��U�ת$��������_m'�_�H5�;�gA��0�ybws%X��p[����p#��wX�,����"2�]wxG���T08/�z��R�P-���%Uj����ۏ�YjB\����e ^����A�J@#����^����}u�]��D�nh~v��d��5
�L�ɮ���^��x�͂���͚S0o��F_e�,��b��K>d^
�h�9�þZ�@>��\'ǫ������͔o|�Z�N:=B_s�@X`0��zEf�N�/T:��f����0����̯��)m�������+KA�zz
7e�	��wn��^���;�0���R��id8�E�T�e�IJ=:8v��M�=RAm���F"Cȁ�=eB��տgJH�v�?Q�b ��uV�O��iT91�B����*T�ե�[�L��P�4��G�ۧ2�>1^�N�)�:P�`��K�gj��2 �UR$빓���P"�f>��A~'�_ =������'���v4�dW_=�ym��YN�i�������3�fˣCtx��O�R���I؂a~�p_l��z���.����>]y̼���L�I�n��P%��9rK�{)�S��罬�d7��̃�@(w:�������rO�����2�x\�Ǧ�mY+o]Ͽ�Q�w�c�8��ƸB�L��t�"�4rƙ&y��"-%5?��b��۾�U{�bh��C�$W�kߗ>e l*콕�Se\)J&��t<��s��}︳�M���j��rV!ds;�y�2W�C?�Vk/pg�u�o���{�c�GthtU��w�du{<6"����TwII����+���]G'J��)<Ӆ
1�Bˍ�L@�^�)�WC������c��׸�%�4����[����ex]���O$�(�.s��c��>E��c�� ���
�kZ��:	) ^ߪ�����:�����j{�p�%��#����@��/�f�}��=u�&_Ec��|�b�a��wU�� ��H	�Ā7��a���Q�;T��lG�J���B	&�K��$�`���J��hW{\כ+�8�ۍ�fĂ�Nۦ�~zp�6��yt�}�gk�@���3���$��ϻ��U��X���it��;C�8๮��e�9�ڿIY$ T���q��Q�\T$H�0t;�W�6��&��Q�4�bd8]2Z"��L�3��|I�G>^��PQn}�W��\�`��QFԘR�'0��9�\ibWP�Gk��u��G~�/d��,d�w��6�%@��{͛2��ݒ�8U�\���_�'�����Qs+����G�f�^o#�O�d��kIF�o�HAC%;��xF�jA����"V'�g&�f�tLe�U�>=�q����ƌ���ZcxU�u<���w�h`E	0�x�~E���<��;��`�L#Y�v�Ua1�.�Wf��禡�Օ* ܚ�>)�՜�L���3a�[�P���|���^�3E��p_�ʄ��쟾O@b5C4T���(�?�@g��c���Q1���  ��Q����[��"!YW-l���"�P���䠪����suĥ��,5^���،��m�Go�`�H�]��$l�\xK�C_���V"�%��Iz곷,(A�X����o��jl L2���2ӵ��G�	?�E�W;���~�
����{SB���F�����~=d$�z(�d��(����5�J��C����e_N�՝g�TT�D�C(!M���x����3f��4.ik���BG����1~x�C�Vp���cb�d��Hk�O�qŢ`�ƫ:l�?E�͐�(��Q;�n\	p�X3t�P�a�8�����~�u���,�4���n� �2V!��G�Un�b}���:�Rv���x;�����}�&�����/�Mw����?H�c� ^n&FF>�k-Ϫ{0����&�Nh^���C���ti��:�6ׁ�%��� �
�I���cw����N�u�8��3�e���'��fHkI%�~@��F���L�����?~�s�Q��۽G�{3K���ix��/��d��ޚG���u�a�q�^�.�� �e�ڗ���Z#��� Q����Ǚc�᠂D���;�T���J1j����FJv�ˤ��o���q�Y{j:w�����J�KӄDU�)�B����P.ۭ}�� o�@��Z��kQq%��<s����`�`��	�`�?YVF�1<��s�ʩ��`a�Y�ˣ�קw��ӄ��!�۸�.�}T�|��j���Z���'X&bj�^I'��ݼ�p(� *�%�9��\�a������<���9�'5�^Ԝ�	,J-��h�Ӕ���&��������E9gB�������4�Mo��7=�S{�@*��<U��QW�i�(�Ҋ�[3J[��n�RV�A�}
�{~/cF{|�Khh����o{�(��R8��i�s�{(́�[�o�T��f�r�=����b�&���f�`t�G/��mex(T��jW�����x�������ugCX����z�	>��z3�v��l[��Vs�(��:���ت5��f���U���r��Id�]�HQ�5����k?8�Vp���P9{�QK<Q�Ο�DeI����U[�&+�	ؒyH��R`{!|8jH0��GEw;��ŉ�">�(C�}ʛ�$����+[���?�R���r�v����>@mi���joj�A����g��ˤQ�~����& ��N�3�͍ǧ�P~�^�Pmh%�W`&��(�b��:��9gO�:5鿶��h؂1�@���*<ܢ��$�+1�h��v��[�V���V�c�cN�V]�1 B����ٓG"!|S]��\�l�m�3�'���7��@K5䨄�^p�q���Ԁ�0���"��^���>[�7h>rJФ�Ѱ�.L6�OQf(JI��d���0/7.4�I��	8�Xȸ6���SM{-Vb8���c�%"Q�t�Q¥x���(!�Ej'�bΎW�&\��Ǿ�ۚ8�����S����sߔ>>cr�?�3�Ej\�I�9��l���O6�:�&)��!�>��Q�Qf�9�pk��k���n3���;���̜7��xna�/b�	�R������=|�Ψ����t<�s�gL)-�>�!S��v�,�|Ӹ9��'���>�h��E08R/h��H2�W��kI�ʶ���/b�B��|���cA$Rv�rz�G��!��J�1��&�P�b��s�ɾ-G	�]E%m�@ 6:�N,BEQ�Ծ�0�u��F�bn�`P��.��V�|�U�q�/�{��k�ٿ��|�o�H�+�;_�h ��sA�ũ2�?�U��ӒN~���[ (��~��L+�W6 ��R�,/��m�o��c���k�:�#%!�lE���S�*h���'q�W��'/9����{g��{l�Fe�, �h�]�c���1�Vy��8��MO����y�k���_9~�qT��#M�#�H|}08�bnxݢs��<;{�3z��F5P�4E΂d��������2���sinӻֵ�5Gn\�J�F����=�t� �G"K�tg㰝���!�+�o�"R~g���,Dg�a&�s�o�ErYg�a�QA�W6�*���9�rh��)�iWs���h�(1������3O/�ʆi������(K�T֝fT�l�b����bPE?ϳab��&)8�ÕEٖ�X��|m"Sm>'�gZ�fȧ<Y�!�����
�C�9Ϭ��N+N�|�
\'k�b4ӏD�r��!�?Tr�b5Oh#2>1X�c	�݊|C���0����0xh�X��������R��?s��^9�uV�/�H�R�s�`���@
:�;%��7��7�y��W��1�R�3�@��W�'����h~��밸�7����/F�VC����5�1M3�9v�re,��?a�9�{�� �j���]RJ�HK{��|v��\������^:;������.B��F&���Q�p���O
v�T���_���4���Z˓�P��	i��R"=�E#@�u ��}z��R����%H�"�+��
\����P��O&�"x`�ujr���Z��]�f�6�=�a��W��0��99`N,���UÎ�	Br�|8u0*1T������Ξ�$��t�Eu��6�4���.�3]�s�X$�� ș��,�U^�������_�g,��ӂ��'y����aj �?bz4���Q�y����Q�he�?�������و@I8�� ɳ��t@.L�<��d��g�ҍ���$~�W��{���s�F/��6]f�C��C4� ���>A5k3�fq�}�~yJ>xO���.U;�f�s��>�~iP�֯W*���ZgɼȩZ���O�i�"�n2�gy)^]��Q�G'�"��ff�����9M�"��2u�1G�G�9vX�Ү����6Հr1R��|�M7���������s�+g���h4���)�7m������mP�Xا�x�ݮ��G=�n7�So����^q�3H�$U�yeq։P����u���-X���L��~.p��S�
�?1f6�@&U���Eu�߾���� #���+m�jX��%��qm����_#J{�5����x�[���cWN��
��� h%�X�xM��� 2�>P��9Z|t��tjA_ˡ8���q