��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ��]��Xȭ*�Cf�*`�'/�9gS$��Sh��f����n����+EhM�j�O'�yz,�_ ���)ZN�6��dQr�p�x�y�C'�m��H.@'�!ѽ��Ќ����M�P�;�{��3�OT����n/\�@���V�F�	G�V��]� z�`t���y[q����a2X~�*���O���k�<Ζ�?
J��I���iR��eϴ�J�Ij�Je�V�e��JB^ �9�E�|�h,����� �������c���k�zbr���A�5b���J�f�"UP��"� ^$wW�1�t�Ў��	�/G>�ڇ�[mȺ��j���K�_���)ϕ��4�����k-�mVs/��͆Cw�$U؇�/4dY���J�=������ ��e[M����
㌞c��|?vNqs	U�{)�ic=�$s�o�����F�/�������.����^+��t�7I�ΏY}Ҩ��)E5��'K��z�F���40�m��G �d~��e�<8��a��d���J�A�i��4�[���a���~����Pz��������*=���{��Mn�Y2���}A�Z�R�+X?��
��F��1�
 }��M�t�ڑ� �-��֧iյ�A�kϟ���f�h	 K&z;���d�IX����"d�TM��{>4� ������C"��U>3��K�;�0�~˗DO(�8	7�<T:�H��(8���v=�yX���^
��>2�U/�����T�9�\�ԍz3�g�.����\ډ�L���n�G�\��F���ډNR�Uxǉx�.�Jys)��@p; 	�{��#2{�u�B{��<ӟ�;$������;2������(����������#-�L��	�3�0.c08ʑ�Q�`F�&������Tb��YR��c(�P,d�)�%Ar+�]8�4�h��i6����R���}�}�'R��D5ɐ%�+��]k�1s�/��z%F~�h���5��)O�6��}�ށ�TlUx@�]�3Yd@\�C��5���ѧ�
%�Á�H6\�\c	�C��f�b[�P�o��=���!��.	f�ḵ��V5P�p9]��|��D����Kۨ���W�h:�3�V|�g�㳤'(�YE1*V����L�x��G�[��Ӧ&լݫaIC����<�:���)#�@����^`�^��f?5�C/8!Ia��W�����Z�����7��:+����K2l}�`�LꚀ�'�Nt߶>Z��Jz�f:��I�������zJ�\��Jk¹������
m]�Ta���t�8��v^�F����؄�jd��3�����*�w!l
�i.�	p�Fv�� %ܕ�RX:>��E|D����_�"ix���|�8X.�
D��㥴j�8�TI���O$XܞO�H��NnÅ{��Q��j����KBf��"���� \��,"��Ӵ��EB�_�'�݂�%�PZ2�%V���2f�f��??�;#&�U�� z&��i�s��ƙW���0+8\F�/["�EN�
�yw �����Θ|k���0k���2@��?�V�يC�NZ�7gM�p�E_ �����4e��v�9��� `ޡ�L6��_�Z�4�6��1�)Yue=����罣��& �S�x[�3*LE���	wy��.l3��p���=cI�xǕ!�\d�8�v Tkͧ�s<�4FK�V:I����"�D�D$*QY[�v-��=��[��9h+��j�ʇ�0�^[}kU+3Q���խ�A6���AݘJ��+gڇ��٩5�Ib���&#��;%Ż ~S,�@�$��2��*�quJ�8IT~����IgN2��8HiͿ,�K����K	��TE���N��l���i���E����g��V�8 ��o� ��!�23V*�<��qC�E첗R��[B�sQ��M�Gu����I���g�d���x��.���o+����K���_i�E��-Cuk2�j�h<o�� u��T�?#r��D��_u2	�L�o�2�n��'i1(��цMP/�z�a�_MvN!�&�'x��/��$�D�I��9�Q�Kl�T\Ss�M����F!v�y7h2~� ��3J�� �L(���Mt�;�M�I�����a��E�8'I�����C�|F9-�,{��cQ�+���4�*i�K�9���bti��,�B������މP1���"���N�_I�p.�+�DKI:y#M�v�p��QJd�С6�2���>¨���M+)b�֚~�N��]ubk.ϩ�uE����VL�7"���^:\s1f��):%��Z�����*1���]E#���,��f��*bU˿k��h��6z�`+��(��ji:QZ�!m�S����ڊ�	��/��Pԑ���u9�"5N���=
��9���\��ʾ%,��ǎ\��1�����k��������31p�D�nd�&;��~4���}�s�3�/�q����3Nck|�.��)an�����U������⌺�_�;��M�2�(�z|�ytbX��d�7h�_�]S:�xy���Gctο�hy��.6�į�����7<�D�~(`j�t�����K#�kgW�(_Ƕ�"��Wy�޶���գ%7���<}���QWA\��ʸ�f��q�c�R�˕J�[�I���K%�u5�M��-�92i��N����)شf�%j2<?�f�Si*�,*���F�g�L���g,�sOܿI��C]�j7��?L^�����
�,$�4 �]Y&���v�&�B�t#b���[����p��FF>�Sr�>�E���,rPZ������>m�_D<M����ӈ3P~�h1P?'��F��G�%8�B[lJi<��4���G�����5yx�� �fޙ�/���x@��%�{j�k�B�1qygt򂖣+�cf�d.r�¼{�V���5�)y��(�Sm�y���n�u@Z;�Ų�+�&Y�(���z�=��҇�cT����^��G`�5�4 9�?԰�PG^��F�L��N'=�M���UY�����`�0���f\Qqdx��8�q6!���󊻠A���]o��%��(��z�,%(N�r:	���Y�n7Ю� ��Qz�m3?1��В?X�;�O�.,�=����:��;�J8aI[;�í8t��.�#���yK�`��n��8��uv�`'�E�tީ�N%?������!!��^��A��ˎ~�c Va�u~SqBa�y���ȟ���
�����:a�Ct��d�}���<��w���0��|�h:�ۍ�P��1/��tϏ���C����o��&\��]d7p���EÌ�$7�{4������y�*cW��ASX#l���/}Y��2�>Q�@[;�t��Kc��d��Ct�=�AE����S=]��y}\/�?x�-�)�,�"@F�6/$���kl`L^;D�^��Ad:�ʭh�G�*Zw�5��C.��-��u���{��_U)L��l6�FԵwr2e?���9����h�G��5��{�>��S�R�o����'�n�2^�;1�*<YT����_9/��IW�	�p�'��;OĠ�z���®�b?�1�V��;UI�����Ƨ:��|��ٌ˞_�m�I�(�ꅀ+7�m�<��qe��:�z��,bU�KĸUs�穚ʲ�o�f8���O�B(�)���-��^�p}�.H�爟�
���R�GK�)+�(L$j��Ş2s;)�G�B��-^���e�N��y[PPA�8�J�YBűDU�错�J5�c���^����ɿN��viq�m%0�Ͳ��ca]M��|��a ji��P��G}���q�;I�F�����;�H�������dl��0��j���g[��-���U�]߂������#7!�o`~�pE�R��8��J�w������:�g;Q9���?m����o$�<����~o{��£���8s�*Ay���a�;����1N�-�z:\�y��(��V0��C��y�eC��8�@�O�XR�TGSy��M���@Z��)`��mXӧ>�/¤���u`��c�p�!uXV�BdJ��,��N��d�'s:n9d�5��{y��  ���@d��<1\ŖI]�9*ʴLxpl���Z����GX�����aQ�xZ���Z0�d�o�~ᛙg���8Q��v�D�(�ե�XWN���]_��I�����9�]��i�1���(�C�hEI+e���H�6���!!�t���	à?3EX�I������8�Ux$0|H1��bN
-�'�<dce�Y�C��m���A�����(,UG$䒓�6��Ď���$��e�Շ����1�m��@IZ�U�
����;��F{{�(��(�]��qw�_d(=�u%!��Y��2O��-ҝ�͑ i�FK^�#T֦> �y��̙�������AFi2m4��3�6���g���՜;�|o�{�r�Q��,�\�-�I0�x�x�Hx|�&
��.��$���5��Y2['��iS|#�,̤���	f�K�3��J#K��x��K�J]dC�K�%�6Ax��숁�l͵:%`6@{H��A��v�����lmf�C���oW +�M�\�����v��W¨�V\~&�d�1/0�&1�g�@����D��QR�3�QF }p;��ן���;�?���ϥ(�L�ib� �Օ�AF��!?�b}�mkEok��8_�����H2�"��e6�I#���dP�b�*������.64���]b��J��⥱2���&�ǐ}+�A��x_��b�FVMAM�rwe���:�Vr�y]�����4�P���� �6Ը��X�-�����-A�H>/�u	�a�F�?!��b�ɔ��+bɰ_�Iv���
D� l�;��1�7v|�	��~�$K������_� �!�a���uL߹ĿR��uyB���?+p:6��H���.�Wv�,e�8�tv�S�
�����?պ-��Z{t5f�aF�%��'6��`S��TP��L�H�����(�=��Vt�`�}1G ��i�vd�N&�$($gJ�w�=��\f�-���>MaD]m)�9���]�l�F,ۡ�$q�=c�Y^�|�}Mv��<u2�T�܏�8/���n��.�o@ˮE��}��[Zc��kM�"D���H(h�:mYH;�����8���:_���&e H�.�w��|��2f�-��Ȕ��u���?�B�����7��)R�ށ�+��4��d��I��G���!E
q�Ps;
SL�p�,�C���J{��fs�*�/���Z�7��������d�2`�����Q��>���e&���&����Uܲy�S��W]
2��i��k��[���n����X~��<��P�&�������#Yl��cG�ݽ-ԗ�"��_u!�6�*�k�Sa�]��|��CNQ����Ƅ�)��J�2|	��@�B:8������g��B{a�f�x��[A���4��@��g��#wqm���L�a"0,���Y�Na�پ���}�����*�������}��w֢��AI�\�;�8�52+Xh����Bf�� uϰ����7�G�:��k)C�r���y;o�"OsG���R�Lߕ%�oIL�s|@э����7����?��	ýt�=;��g�絚����4�A0�$�	��d?��։�be
!>��� ��MP\:�#$���o 6�AD!ݛăg�I� �`aj �P.>ѭY�������U'��!�Hʼh�*pd.h�\�+��A��\��9�'���fr��\A���q��������&d��_�D�`;�� h	����T�}�Oy�W9|��m$���V7L��'K� 3[�M׳x_ʧeoB�@TVU�mg�t��F�ʯ��q��2��l�A?��JQS���=q
U����ĭ��O�uW��$��n��0�',1;݁s�	���(�c��9��n%���	��Z�����5
AZ �*����g�00�u�����tR)�G]Cl���}2hUVJ>>�3卺-��f/�f�Li<��Vxޖ��2�ч���ı.���c{/�m+k�zS���qQ������i4W���qM�M)�<����p�ҹ���.��ó	����y��w��y�	��[�2�2 �X�B��'��(�֬�_f/X��x�G)+�F�LP]���Xu��՝������̀��<4��l��"nk�j������g�zr�ǆP�V�T&�?��O���p ��tF�qb�&�C���K��[B�)�ila�'<��Q�>:�h�M~�<^[ШT�	j����#�,��tu�#����gs�0���4tC��10�Jp�������:���aa��}5J�!�jW1^������%eeC/�ДE����9Q��2a��h����T���4|.���w4XW8��S���/[������r��ґR�c}��W>� 5k ����94uFN�S 3�m8�m:ܙ[Y��	�Mo/n]�z-���y&� ��B�+�s���ط���|���}+��p��̈����I�rl�]����|Xs����< \��|�*���m7��g���0jxp�%ɹDk����^a>���x��vqҡ�n5AMR���]ٓ�6a�rp09���*�
��7��%���s�#�V��D�b����(�֡�O�A�y����5���C���$!#���M��ԍ�Ś$:�'�F�=�=��P)!ck돾Y�n6)��/�z0K�9z=G�6����@����?;*��Y!&�-j�m�;U���ȐOӍU�4�B$���:� �9�k��%�������]CԂ���Pv�◸�VQ�4�Q�_zPI��8�ڟ�-|̠��mU������9���?�5�d�P��G�=ԇj��lQZJ�UH�����"�kD��4���U/R5� w��#����
���v��u���|^O}b褑�/f��)�5�@{������wM��M#@�d��-�ĵqŁg>��Pd�⭬g������������2��f��D�3J
�-�X�<0X|�vN9���mWv=ѾP���%�����l��i�W`oҹ�p����[�j�ޙУ<Q��
�kB7=*e)S��a�������A�@�-�-�WŖ�E5\�I���*V���u}�e�1��D�'���:lw�_��8�kcފ�e w-1͈i�S �*>��U������Y��&��z�Nj��N�򩨇5��7K�GE�"]Xf%���ͶYC�+;�ڰ#��1�xT�A���L�fO�t4�@��R_Z����<>AQ0\�̂ �[�X8�#i'���C`B��.t��.!(�A� P�����d�L���f�>
T�;K�ef3t�s�p3���Y~P��8\�!B���eM���:��xv��c,e7s"5	ì�t=z�<�?!#A��@���̵gCf��>�Z��'����fL��AJA���}�R|B���i��iQ�Y����$�
3�	\��jZp7�v�$e�_��?L�Ĝ���	o��,pid� Qߡ~��5��h��z(]��ņJg9�f�`��o����+�Cp͵�p3�t�v�C�'(j��=�e1�&"x}#Y��MK�Y/���ꙛ	%�:]�1�)�$���M�\�h�&�Zz�')�A �3مl@�D�Ԋ�.�W�8L�5���ᓔP⸐2['�Y�j�o��i(۴q��E�mG����W�YM��.!�'`?3G��6,�eb�VhHb(�$J�k�2����@̰�M��^�[�x��
���{,�D)��O/�ι�l~����R������N��9���D0�ZYIVn�"��|i�9��X�i�E50?�r��}0
�N�n<�y6��WX��+
f���+� d�91�7����xԷ,����i[����):ͬ�e���v��{J�(s��K�g��O����ء Ef�&h�
��>�=�a��g��"�:3��KW�"K���"8)�V�TLQ7
(se�����&�2��� ݲ�=�7�J��z�Bɸ��e�E�MqUزT����+4�g� ��$8ҋ@?n� S9�X�)��P�k�ZEW��:�ڹ�p��w��&�G!8����zOHOB-P��K���h����ѼM�\�9s\ɜ@�W�ЎR@�#��~�mȆ!�B����g}��y_��p���������w:uYN�'_��s3��3�z�/0�YA8+륉 ��[ْB��%��Oe��j1�\]�[/�Z�:e�����U�����n�i�e��T�f4�K�zW�)�~(�t�ú����:}�a�}u�uy����X���m�+�����|��(͉�PA6g�º�(���-`���ߗpt.R�'��f!��7wϽh��Ah!������r�ب�]�q~{dz�S�yY�b�z׉n�R��?�؜(b>����[+��w�_��T�d<E!pO�w_����+M��v��?��K\�j�;x�,p�[���O��>��ZEB'�jCt�\A�����Ƹ!�9AG�o�GP�ߋ:,�[	���O2������M+�V'#X��-Z6�_�2��\X� �M'�ҍ>�M
<�l<���bV�	�Py�x���F�?B�����1�xe��I�|ϒi�`��Z�.���iۮ�3��R��-U5z�p{�t`�iN��$����l:��@�����T/��m���܉A�d.	
m���#��m���Dz�B���Je�S�lTu��y�ᾥ���'ߡ����V�ږ.�y���ͳ �=ĈzL��J+%����ĺ`��?�l�(�eT!��a܄�����$��\�"{��Y����@�1�Iy�>-�m��P2;�X0�O��'C�^���s��i��8(^A�j�1ɹG^?��6�c�j��[N�qi^�-`����@�yL��)�Q����e��V�/���ꊆ�!��'=�䅘�w
�AJz�Кմ�� �H���$e���¯���q	�PY���
+^�?�JϠ�c���PP$@�j�m� .�׈���e	�eA��!G��ſl�R�'RV��uMGI�ѷ�E�̥.�"�{�47�xg�$3t�O*]Ob����W��z�����jጥ�	Q��c��*�l6���l}�L��<�>+�3�)-{Y(����_�jA���cih7 еθ>h�Ǐʞ�8��D���s� �����ܬ� ��"����'lM��~�v�ON�PȪ��g��V�q<.ݭMC��^�ځJ	�h�����	���B[O���A�u���!5N�8���g�uA�Ĝh
0拢� ���=����M�4��N��puVa���[M���t%�:�p���
��Z��v�E(ݘ��"�
�> ~���Y�4+/ ����@�D����`q���nw��Ju�J�6�����|��o�U���i�3�t��9�yx��y�ԱZ+���A�=����{hJs�&�PKe�ޘm��C���φ��r�[G`rKw��jK�q��hu�>6?�j�ʺ�)Idyz*l6S飭�a�����}�cЏ?����u�B9�~-[ �4f�uW� �ղ����d��̈ϋLZ���~�A�>6�	W_��5��~ɐ6P�>��LOA�9S#vN��3���ة�v� O�_CM��Y�x��}g�%�|���x䒻�6��u`���^D�b��O�FxU������
�6T�����N�󼍆���A��\����	S*hغ?v{���ʪ����IЫ��o,e@C\�8
z��\i���wX�/�>pS�>[M=Ϊ�'1P ����|��rRuW��������ف]�� ������CtKH�ITR/�~f��y6L�{fid���Ws�@�co
q�H��e���Q:�W�=��T<������3QV�@�[��G�e?Ah�~�Z,�6�����yԜ�X7l%���kBa_��(v2mQ}�[<��w��.Y� ��(�`	��iS���8��d�<.�?�fH�K����"��p�pt0��aS��8�,s�D.>�:��H����?�\���� ���Z6��X�t}/�s�p�<�U�o����tN�zD2�7QB��4�;�����6�2?�A���~FO�r;�� ��B�m"a@�NW9u֡Ot�~d�	cJ�������b���"������uP����S���y6W��T� L�z}����7��Aa)5�@,8���Gv/���7��qFG7�}�+|u�+�һebRE����םed��	�ō�&M�*|K B+�QB����LD}�faܺ*gh��1m���d�}�?���ڕ倇���Qc��-g��`���=�J�
��a���`��I��мj:��q�ZR�F��Gя�w�K�`$���'ѐ*5lxq?��8�Os�K����~S8ֺ}㒙B�m��'�j�9#�B�Y��t�/¯aE8_����2�<�4��V�:��Z��~���Q�Y�=��&P9��lKz� �b4T�ow�wEd���˔Ɠ��8�)c���1r9��J�Z���|'�Vz�9�;�SC�Q���.�U%~,���F3L`���`8��W"�2V��m��,G����%2��\���{crE�p3�w��O�pa\�gn��mUQB���:8YL�fc	7;gsD�e+�u2T��΅C��9��{���d#Y��x�tO��aj�����8}ݿ��]����S�gLG1V������[HF��:3�n03�M[
�%������nU[p�Z�XGw��F�l�����`���%j
�:��]�ɨ�'��B���G��J�����ڻ֘(U�W:m4��1�uD� b|�]�G-VЖ/O�?���'N�{�s|��� `���r%e�����^�������5����sl[�;ᖧ�'�1\%����[3�1[4�:�i��ܷk�S�����nT:{.��G�ĳ��@�:Lw�Li� �^��u�6Ƞ����YOۅR���:pl��J�����`�����ŀ����1����D��0?rͨ�ˤ���[I��3FK<1^E�`��_W��]�е����A�ruG��=T�aP�9�S@6�i�)����ѭ��O<)v��p��b��b<!�K, ��?��8Q�t�QX�$��t;σ�F�TȨ��#��_a��[y��z{��6T�Y�q�����MC)6���Q��
if�BqQ�����r]c�1��l�dG[8��R����z�N`���w�����h��	& ����p�d���"�г��
:󃕅Xw������,��v���� o==R������i���W��[�"�iw����2uP��-[�jy�D4-�yM�V�=��^v�=��2��e�D�t���<Ź��*Bϼ�,fs�N���QL�~��1�b/HѴ0&=�>Jm,���g�mFر�GXS�Vwue����#j�	���6�X�2�6�c�
��O�R�fnX#ʿ���ϣ4)�A�~�L���Q�
�]�M�Y�8 \�?2-Nȭ�j��$|�_��?�)�y@|ɷ^����aeG�I V�+;�	n��@�x�d��3$-C�\��g���mZsnv�ʪZg���K��2��&r�88�.	V��Ji{p�����M ��"�o'!:
Yrv�y��Wc|�4��_٭�R埜��q[�.(7Ր8��i���Jy.�5^xoCe�'�DMz��Z��d#T�dI��(6o&�c�zz1�l9���X3�����"f��[9�/�M�,)��1t���"���@)$r�w�"�bc�c��v1����R,��B]b�����^�6�V��{g�\��Rh��Qc.���}��L��QCgI�W��ng��l��� w��(��:Ďh� G��%К|�f����C�Z/�v�xXG�M�7��{t
}0����,GQ>d�g���J�&�<U9#����� �d�~�2�d��ǩXaF��Ѭl�RGB�o9�l��I-[y��+�e�ą��$��$L�O[�[��<�FE��|@�4�U�42��yd!f5�����G7�(�� ٬oC���m�H��ŀ��:jN��ov��و��,��XƆ��Ĥ��?�]��M�.�g���p�s�Ig�;�~�Y��n�*#&('�08�[2��!���{� �O�u�,�C$QZ�$WT�;`�)����x��XQ�Cƨ�{�B#�&�=)�<��[�}��v���6nE&c�Y(�C�d|G������2�5�����j�ow�r;`�������B������~5��$�y<���]�a�6���wa��0�޿�'b��td�!4,�E�
��e�N��υX�4�=_��)�:�5�X�:o��p���W�E�qmFp��ߢ�B�/4.�s���xO라��Q��&��8�!��j�`��e�O��KLW���	<�U�A��6�pm�t�0!I��6N�����`(a�Y�	�BRT
�@���Z��\����Uۤg\�Y"���׎�,����6��2?�t�h�cz%o-�������?b�t�H{�{
���C�9�-��5�O{��R�� ��E�������G(���BnF9�`�s��r�z��=-����hǁ�J�?6f'�N�e�m�+�SI�ui"FQ8��|�bP^�Rg{K ��u'@��3���4��r(x�)��>�B�*S�#Ӵ¡H�ɏ��c�ln�@� ��g�֗K"�,�T��G˟@��"�)�jB�4o䇅�˖���Z�҅���k!Q�W}�gqK��yW�N��s�7x���t��/���b8TM?�)vq/��(��K/��Von�1[�J�{�]�oV��XD���:^�n{,�elF�o��Y�=Bc��ޥy>	L�a�U�Q6:kjT`�/n8�ԧ�����V"&�v}�!��C��P=�j�/����칃}�)�*�Qt���Z$�����{�-h{I��T��h��T�qW5ťGUt �X�X��74��H�X�U�G[��,�I��+H0p�T �s����ʈ�7�毁D=�V���u��U��X�?�eYX���m{M����Q����(��[��f*�����c�c���G(��_X��S�=ĴD�[0����7�
�����]��+�1��gQ�G@Q2��1��W�m�"��@z/����ŕ���\��`�o��B�[#T~�끈���?���~�D֘�ո�;�\�X����!��g��q�!6����D�������������&�	�0��V�l��uJ�7�[���(og	ʨ��G��c�Ơ�]9p�x}G7�S���vkuB͚KС��QT�����/<<Vj&ߞ�����6C7Y��=L�譒�������}t��8��5?��l9�*Q���Qa��-$�P�R�$cL��s���(���.�ͤ�m�M0L��g.��*�WЍi�NH����h#�TXƺKȫ�j�� rPr
V��:I�F8=�n𥤐��!F��@KI�H��0�m���=����TAJ�(��v���iV��_a�����k�����ȋ@������-����8��4�H�6Y�ܸE�8�-r:>17B��{���������[�=�}Z���T�|���}�]�7�6߈�-��޺������)^N. �ANѭ%o�L�����N��3¹���9�xn�¡ �c�_�8��ߏ��>�G� G�w�X�!�z�u[�>2��t��?\�'�(e�b��-7����ͪ4JD\($���.}����Bf�X�����E��l /sG��s@�A���7b��a��H�g�է�={)�������.���fr{#�������/6Q6�	1<�P*��*j�������r=�ѧ�Ӯ;V��_��cq/��4Ǿ����n>Z��Q��8钿������� 	q�"�P3B�P���`��֧�FN)�$z��9�{éf��������z��Ck�9T�|n��d�����Wٟ{4��1�+�)\W&�+�R�0:q�u)��YP��*w�l���dA������֪��!M���i�տ�ٝ&ŗD'$SP�G����LJݻ�����1MO����p%�G*e�׶94Oy=��^�Vhi<se�.�`\�b�����]Χ��5��9yq�r1T����΂J+%��JY��u��%r:μ��I���!�}�4�ſ"��I�1Y��Yd�tJ��T~t�����F��SgB��'l��=�!�F�lfT�ZB�؄��A�kWY�,Ɯ<!FY9)�b%��
�l%��?����L5���J�V�g���X;��;Wy��\�5� a,��9�>�|E��w���b��먔��B]��b��A�V�����z!)kོ�m��l������n�;����p��[���%h���1h��S�;*@�{�2���� ,����m�6�eV����+y%�8̗�+�;�����I���m��^��@�2��Vt������f�ɍI�X�A��NPs�S7�urX��1�$LK���>*�;��A��KP��j��SmL^�r����ͭ	�zd��S�&&����fO��8���	�!�]T�Y�Qհ�"���TL��s��0]&ڴ��[�Oh!���ڥ�;/�XN����!?��Bשȩ�"Y+,o��|6�(�'��E��`k�n��$��l���8o� 
�-)C�'L�˙��?�}����8k'�ؐӽ�j�ϔ"��?��3Ǽؘ�t t��G���t��0ۄ��.z�\�>��T�c/�K����l�������^�1˛�麭EA�_�����ʎR�`��ӿ��&"��lK�~!yL�����9;����DA^�� �?���5��;�a��!;iWa�~�<G�|�4��+����5TŐ�ُ�t��O����]\7�B(��'5o�h�/@��_�����C9XNS@��uG��9C���vmi��] "q����9��x�8C��,����$���W��ʹA�$/��-k��M#O�D��[�U�M�v�M��*��F��E����tQ�Ψ�٪�FK]�?��W�����"�*ϑse�9)�@�o�y�����a���D5_��h��xn�g�*E���Yt�N����"��9T�¹��ť�h_{�d��Wy�_��y_���F�6D��dnѪ��k?��*OG2�w��yQ�Дǝ%�j�����|�R~�t^�
������~;q`�(�mL����ݾ�U���qm/	o�%�~)J�[K7K�R�X�h ^D��g�����	��s���Ȍ �ݑZ�F"�3��]g�N���v�\�Z|wͬ#����b�A?F��;���#|���\��h���8���������B?�^��R�^�_G�Bf#,7g�dĻ�G��{�F���c���e� �K��|$��+}m/��������@zu?�WY���v)�}p�;�_�3�m�V�H�_k>�Љ��W��?�R(����0Z�.�r�a,�.��^k;Sdל���z������'��w��� J��?|�ՄC��7���y�4�谳9�wuf(�cV�E�����M��2�*2�V�����Z]���{}=�rpd��������06?���`#|m;�*[Y3�`mnqˮs׿W`��́�H^1�����l��][�8Pｹ�x<�7x�/^t�h�8~�t+���P�)Ս�����&J�\�%����!�r��1ZB�{k������~wB<��gq�b%��N�A�G�K����VX�V}�Ώ:o��,�+(e�`�7��[���ë�}i�f�o&�=�R_[|���u���N�+�� �Ϩ?�ĖYj�,�����C�x����MTfY��z��;W�w�:;�_�A��+����;�Z6Z��>�u�S,4�8.|�?��@�L�S4�K���ӀM��X��g0X?G�ޝk!"r;�2ѣ���d,�q�wPoSυ+�pLأE��w��<<r�4۔�G��zoI\;���2����^� �+BfT�p��G�{Ɯ���?cӻQ\��s��ѱy|P#�-��Xr,��i�O/�Qt3�]�C	),�!Pi�uվ���F�%c6���o#γ����3vI��ʊ�ۛ:���0���'	v]	�C��U�����8�$���2si6�c�k�#*�ɷ>���� ���n����;�P�u�=䆷���]���L,ĩ�4C��n��LbJ�j��\72�(��1"��Mƅ�}4�C�=(�v�U},`Ϫ�5�۪Ɛ���fS�>/�Rt�x�{
�Z�ܛ{nY����-��t�4{���p�&�k���-R=%e�X�NK��&I�~?WMu:Z~֢	�ub��$��mC����X |��������	��CU�(1�	|��"���R8kE���5�U���c���AO��>�v.ɺC���������\̈�r�+*�yŤ׸����~��,��>ᕓMG ����]����5��l�d,?ԗ�3���/�.��E Hn����n�}��f�-S��Fp�M�����$�~�	�-s5R$�"D�������'��.�6���)�w����BŎ������k��I�xŚ��K�u�ׯ�������ϟ��Kx��F�$�$\M��x�k'C��3��mxp����H������_��O&�V7~� �_���H�=�ip/��*�=�n�AK�����r��7a)���?iV���t*�:��R 
��S�{�a���m��p����k����( 0	�6�00mG�Y�rY;�BRZe.ɐ���kP��/�4�ᡠ��̺�%�.=��o�»B�e�@U���&Ƥ(~��=� �|�ǧ�[;Ꜹ1@K ���ؘj`����Q<q(Y��4J�:�"�50�|&_5x�U�M^Z�r�e4�:EM2<Ogn <�y>���;��Egm�i���F���l�|�Q�w���**�jx�C1 }$�G�Ԓ�m�1�«S��|~ :jr:�
_$�}!%�mn��M��\��Ĺ[S���Ȯva��"E�P�:�Y���
|hn���#�U_�X�wM��u6�|�l�A�ƒ͆ �\��f�=Ϊ%�4���xz���M
{d�6�`Kq�=��SѠ���tDuKՋ5������'n��{�����0��>��%�Cc`a̓[�����MF���YMK�)��D���.�#�a����
n�B1���kT�X��  *�k��e��\'�H���uq�����P�����T�^v%�
j�:�U�)��h��l�Ir�� �.5n�Aٸ���O���� � q'�{�Qo��=�Z��G3��ķ���_�7W� @�,��Z7���p����p61u�j�B��r��V�ٰ�K~�0yM�A���������L���ù����q��X�H/�z�	ur�ڱO2��?�C����N�;�� �2�4k(@�i���P��8�S�ĔJݑ��f�
$h����*�LR�nuS�1��P�x^�j�������Y>5+�-�<b���A���ЃPd�W0:s`Q5V�<��ʬ�=?S�<y�`
�S��~����)w��ni��5��(�٬I�ܒ��Ul+�Y�T&�1�!]k�JQ��m<o�!r�y�st�g��Z��P�F˩�(���F�=�ȳ�΢�E�w5��97��M�\e,�ڞ��JQ��2��Ѥ��͚���߻p�8���]x�ߪ�6�q
e���"|��$O<0�'�9��t�,mG���9����`]�e�X�$l�ȵ<�X<U@5Ds%���>�PvQd$������B��_�B�Lj7���Ka5�4�%���V���\R�����ƈ�{�B���7������e�~��RVR��	%�F�?�����4�['�+H�MT>�c�i�U�1�����V��-iX�;��c���/XR��m��.`v��Qp��:Ӂ7{�I��C�6l��;������鍽p�Tmv��[�޸�S�)�����-q�11�)��Э_�v���k��傐8Fm,��52�:=ޛ^K_�8*'�1f�me3+�{@���."C�m�Y4�M3"�/�B�r<Z�Fh��r`�g�.�uǳ_��#|C�L�K+��%�4KV����o�]�3l,��aۯ�� ��=���U�=�ő&۳�����\�}�1b djN�X2 ������Uk�Y'�bny�NGM�<�x� �؍,��;t17�u�N�a��F�+���
�w1��v�E͆8���!=� c���V_���$@C�2g���Ȯ��}ǵƛ��<�Ψ�o}�����Qv���N��⤛Su5^3�D[�d��Ԫ�K�����U��@v~��#8� �!�~�j�v
��s:9��'�v?�o����c��r���2w6�䣶���`��6��������K}�?6o\��̢W.j�S�w�b8����y���Ŀ0����O��ў�oh�]��)Gӳ���5���� A�g�s�����8K8�}"s�`��O���<�LW%�=Ch��������G��|��������j�Q
��x�����u��4�SN3�܅"Zm�tg1� ���H�/�i����j-���8�jM���{i7b�d c2�b���~�[;�G�ƻS�eΝ��))[ޕ��1�w)�m�:&	�S�?q8 L�bf������ăˀ�9��%�`�E�"�Y0�j\�}��V�Hn*�H�'Q��Tg� ��~��l��6���ͦj��![����Lr5��
��Olj"�b�u�$.�w�鳮����(.EXi�)���&.ܠ��7+�,���٠ӀBA�7Pָpy||Cx���L�G��7���v>=���Kh�_�D�iF�C�I�{ϧ�U���={I��#�KKy���s�Ʀ�0C4�0�>~���ه5���ue����:��F�?G���ԫЖjef����.s0viI��:�^��U�r{!������:m�Ӛ�ձu��u�{ɿ��y��oI�eG��8�D��L>$s��i��I<�G��.�Ӓ�n�T����2M�bM'+��q�����3�P��_I<3�K�1�'i��'�XD4���d<A{�^�-���y��u� 0���r���ԾW]�vQ�m� 73+�,�F\�ro�;10��_�r~�����(�7�}4�MfwEd�����!D-�2"���}�w�U��e~s�f�zTﰷ[[��W�V�g��Α/����J=�԰D��?c/�ͲϠ�����QB4�x���d@l��ʙۋrZ3'芍�W6��8st��S<"n: ߴ�����ܫ�,�ҁV�m�����5�;��u���p�л��M|UڍI��)Y#������U������9&��>��q���%�"P DÎ�B��O	���>3,z�/}��rQ�EL�����k��ۈ�) Z7M�V�ԍrŦh)��/�@��=��hft4����JGo�a��Ga؆Ā������}>��&?�#�J������2U���M��R^�P$'��}�uM������Y3��k"��ܪ0���8�sOO��}Q��	�2���kQ�U� 0!3C0��K��X��S���W噰���-�����-D��w�w����M2�_�S�oX�FP��:�ڑT�8��'�C{�	�'���[&l���P��,��#�Mösy�%~�c�����mKߣ�_��������{G��<�Va8�:��Ў]�I�N�Fd5Q_��g-�3��Bl4�7�J�I�[�ϮM�J] "����KR�5�V����g�� &�Sx0e'��*��M��Wc��5�s�7.']��"Q#
����t�AeJ&J=Ցz�4�Kk������?�9�>�Q�.���q=�p^���d��.�����]���Ӌ���&���"�9��5��=��Ca����.������&���C��MX�P���w�?rarĚ��=_\�O��Q��G"Ǐ��w����{�ھ~;���|�qYH�ԣ��?=g)��5�V�4������#������odA7���*=Ζ|��/�;D_k+<��.-�HiBZ��J�ܾ�Z��!�6� 1� �B'[�m�B��;vRVM(+K�+� ���ڻf�ߦ2G�E1����$�Nq�b��z�,�|K;��@��(X��F��M>ql�M_�^(�*�X�C�e�<����S�}�)��J%��
ư Ms͠����3���Q惶I,c���_l�����se�`x�540[�&L@�P�<�s��k|#I��os�r��|FN�+�|wY��]�/ƙ|���e�H�X�gE�[R`���eƋ���Ҟũ[�+)��e�!�E�,�|�nzD� �`l�LH�������O�}=\�tc��i�����x���m��n][4v1�/@
L��X��Ԫ�S����T��^�(EI#�s0b�n�s3�/_��}�}$�L���tJ���ſ}$�C�z�������r66!K$�����;�dxp-�b6�F�����X���l�vݝG����b��:\�G��$�����5�NH���q�y�PvЪ��w�,h�M��&���с̅8���?�϶�*��<�~�����ߚ��D�����l�!���Zo*���Щ&2�K����{m�x �"+0������_����6�2�{�9x�������c���V!��t��(Ьod�:+�����+|y�D^C��p�w�a$i��{�Y#!��2!���	$d�&6EF��]o��>�1��j��f���[KC�o( 4}-K[h��	��ƛ:�洸;��݉���ӊ�&>�-Q�W{����������;�p__w���[p��*�v�	���V�] $v7݈ץ?�L��-6MI�S2�'h�W.ӱX������gZ���c!�� Y?�L���(��Pf��~��{�+��_&�_y��xZ��}�Z�@�o�E*v���[���ΎO�/!%S��'����^��6��ص�<��/�C�����]��
g`�?�4rz�+=26����9���ǈ[�[\�Dܴ��o�Av����e+u:u�i�T^���f���;; V�Ui��m~���ݩ�n�P���P��چ���.���p4~�vG��� L���Gnֿ���w�����m�
C�*��a*�_��!�K���G6���^㒝d��HX�r/w���"���6���D-��k4C�ي	�V�]���KF�����?$�C�n��s���A׍�<Y�?�P��:�nz<�'��'l��+����8��+��^K�-fY��+�M�R~Mؕ=ִ���Co5��G}���K��E���C���o�D��d����i*K�~���=�:����esX=Y6.��r�D낾X��J� �((=$�Dsڟ}���a���z��2\Feɓ�K�/�l�O�[��Rc���.>Q�1�2���+^b,a�d�q-@�Fe�̰��.'����T�Ʀ��5&�cz�L:C��rz,��+S�:y��=��mD;qi# ��-�z�٧�Bfd�rDu��Cl��Cq�o{�⑲���2����Cr&�G���<B���ʻ�%���O�6�ٓ��y��?09�u�Vk��O	���S���p����>#:a��(�ç`h�P) ��CZ:���[��C��<!����ڌ�&?��t�
����8!<x���U����Fuꅱ�E�7}x='!Vb���)�QGو#t2-�q�l��� ���R�blF~�Rt/P�
E�hC�M�	FD�u� E �tF�'t-)�K�|��l}�g<s��(�u�d_�i��Ģ�A��x�K�1/%\@�h�V#��mb��l%���z9��V�"]���υCy��2���gEL <	=j1��]�<ג���W����e�u%����Vy����pE϶ـ?�V����ksM���.u����Cu��oq�����-}@H��Gxh�{��v+y���<�3�_\���ؐ��M��TTӛp���dl�����������c�ӹw`EtzG�Wх.��:�X�g�J�Œ� <ͯRJ琗.�[�yV%�W^�;EI<	OuK�*��'4�Y���\���V��Ӽr�f�˸.��qEjO�w��|/0KCt�ʠ��ͫ�aB��}�GǊy^>���A�g���KT`6��Ғ{�̪� �H�d����F�t��)�������&��._�9�ր��#�;|bư|�z�Rmt�|)�WC�]9��"c��#,�م�H/�/j��b�77�2�V�8��lV%u�C^θ,�*�.���D��}"N	#3�N�f�+��Isc��&Z,�xKݟ�?�l^��.8<T�=���2�$Z_n�i���	ڧ��l�8�8�J��1@���+�P�%�C�Zڼ�-�u%��@�L�?���(]�~�,<������1
Q�{�!x�Q�`?� �$T_$;���
�_�����y<�I��G_5�O���ő��x�ۇ�x9��r���V�n��z t�S@v#�=܈��v�E��ֳ-	 â=\F�a}��i�CS*ۣ�Û^)�=Twף�>��"z���3�3�U�k�s�~�u�P�Q�_7#�͵�(��r��p�gd�qa�MC�[�M���(
�"+���A�2����c,�\o� Lm��{��iy-�����l�����kE]�	���Γ�>�uD��9(���x�zx��d�?g���^�	�=�A��Ϧ+���ʑ�R�{g $v�4\K`m[��]�h�6�잍�V�����ǳ�h������$E�A���TOL"%�I�0����h��R����0�aBݙ/�)t~�=	:�T�&Ƙ�7%,��%��*�O#��� �s�=@�8 �`�4[z�1��� dX�[M�_�����,o�ŏ�\�{������]��H��ݤ��iq�>F��6�d	�i�J{۝��F�7�N�G�f)����㢄�J�i= U�%�B�|�1���\�"�s����#E��J�լ���	̨��AzB�Kk�r��?lf���A�|XW��Ͳm!q�%�8����N�x|�b۶Nt�e�m\ݣ�&A�C��.ye�	N�� �>t!����=��E���a��Q3��t�g��M�1,��{�S0UQ���C��+@��=vH������<��4��v��b��o�g%5fBDm�&���{�� _2�j5K���PD����t|Ӳ�,���ו��S ��gD�?&�D;��'�l!��b��,泐�-�����irU��,yKC~��`FABF�+Q�J�|:�Χ>>"�hxϿ�" �`>�~V�����^��`�F�J�hW��s���x��]W�)�s���iw����VN�����G��f)�A+ͨ͐��gs�Ts{��1��YPR	�Q���F!˜J�y!.竞�z�	�W���Js2(ն,�t��qrߴ��k�*�7�O/m����Lk�3����	xrfw��.��i���A�
L�P���[��)�wy�DR]/���.4?���؛�<i�WeГ��̄k*���r�T4��^��g�\���1�ސ�#�"-U���>y�yv��>d�5U4�!즫1xa �<x.$�d\��;-V-����z���s|�UĜ�u$��fH��-�,6�y�f��r����B��,�������8Y�ߺ�e�X�SU:���nK�\�mL�T��2I�&T��y��'�����^o��+;�A�/A g?r3�q�tJ[����#5�;Ν|v�ﺰ�j�Y�����ڎy�; G�ڊQs2�wĚ�$�����H�n�m�a����	�B�a��x+k�o_�}ԥ��9��
�o����4���&<��p���G*y���i2�}9_ĵ�J�
սD��׃�>��.��I4�\��f��M���TN��ݢ<��0M��tނ�X��}|���B��Sϓ�����(��p�O&�"9�Nҟ�O�ET�t(�D�k=�>�!�J���P&nW���g���9�����叕F J�]�Ua�C��J��$�ӔnN����?���6\��e��"�.����{�A���᪙�ٵ�U;���16��,���!����t�1��a"/�x�Χ�^>�S$����8{��>bRTa���(�~���q �Q�xv:E�\�`�Ò�������f|��Z�����=E�&������Ŵ�"�]���E#�pϙhdXH����*w���JH\�L�u5�o陣�2ԑ��ȅ�O0��v��N�Ȇ�U��Ȥ d��S�F;77z���W~�o0�W�a�*Hc�D~�Ӏ�;'����_y)Q���k8L�O�Ι��L���B�G'~/4�IU<e7�[�x'HVبI���[�Օ>���?�bX�O��[٬�_׀R\��,������Vyy�De�(�RJo_�����ʥ����%�.)=J@�T91�P� ��S�����JF����m���h��t�
QA�r�	���_	��<�KW���E���*�"h����:�9Ց+���q#	��&+E$��L�\�0���E��=6���0)O�9Z��� rWHDm=XDo��g�lh��������o*���DSV�y�`�zW�l�D5[�}��LJ�"����5?<��Q��H#��{%ms�����ݲ�5�oS��3a�F�Ao��jj櫦����\���������c���4�Ұ����$qjF0��j�q!}%�#-K�P�@�9��D�1(�ݗ}�O5�*��-�3q����	������F�f� �Iøc��+��gi����Bc+�3O��X1z��7�sw�����	6�!߲D���rZ<)������(o>����;��P����pD������ũ<��՛�h'#T�.GBc(����V����������7@h�Ys-� `QU@�(��1c�]M��j��7"���u���QC	��W��3�rz��#ݺe ��mx�� >�[u�����*�3
��N�9�X����o��v��Z�ߠ���<_��":"m�fqQ@s&[��9&���)���S����@�V���/�KP���s��N��{���FDݩ�ʊ���"[H+�ę�I��Aʹd�{Zљ��X��-�uy�`����$+�>�=�.<�p���3��Cr]��5�!�f˷���t�@g�1H=}Fr'!���YěW8G���kM���?�%�����x<���/�����3̋���20�wotI�t^\��K��8m�x5菿y�AQr5�HA���I����4��B�-T!G���/�9AA�����'4O�������y��1�{z��%%�H�C��Kњ�D7p��]�{�`#8��6բn��.�6�����@�a%F���3N��в'�G�KӬ��Qj�D�*�\bJ�
J#�ẙ��Ǆ{���1�l�o����ߝ��3���a	]1�r��?8�qz�^,��g������<e�Δ���:�B8�z��+����������o�K�I_ɫ�8ަ����k)�i�y�F��Q?�r���I�]���H<�<*�6��Jv�@��9%tYn�d&�˓�M��t��#�`��k�7_��2i��*0��Kk�y�T��c0Ha��xįN���/I_HЄ�xl�ym)��щ���Mo�V���.��F�����C�N��?����l�(!3>|���N��Y�������s�p_�>._��fѰ�'B��ڠ���r	 ^�H�|z���Lv�p[IBl �f��qܹ�����;5쐭\;A��W����-��r䙂��0:Vh�1#Z[`\�	���,O	�G�e�o>J�ϸ��d����Z���nG����]��YT�0�ojcS���w2�ed��K���c���e�D��HB5��h�W����p���h�7����g���25q�`vl�e����;�  �����n��q��Wr�׵ū`&�IZ+��?��J�]�"�b��.�V���EH��1q��S��"XT�[�ۙyn~̩���6��Z�����?���0:Z��v��j���2�'��u���ɣ(�>xp�;<������+�ޙ��uicQ����΋*?4�(�e�;|>�H�)���G���D�_��n/�w��U���~��_O�c���\����p�������`�����hp����K��wop�FW�$��H�&*پ��atC�#��\_��w��y�~����E��cȼ>˹&hw� �rY�n:��wr�n�S��Cf��?�r�Zg-G�s��PU͘�)������r[�Vo�H��ɬa�=38�u�؞��ݿ4;gh�N� ���ڤ� ��U�q2�>2=_���a����u�ƨ����@m]S���6��:�R�b���-��yR�����ǆ�0�L���֧���q��U�5vD��G��>k�ܥ*��C�{d���5���ǛE�x��y��.'�j�vyf5Iw��%�ю�[ԥ�lP�e��Lj��`#�~r�xDH�vEI�H��R<�M03�K�B!.O1��Ach�6 � A����T�FV&�6��s��Z$�,�����>��X�L]M�_�QZ&L��b+Ӷ�?��r�1Ɂѩ���ͧ���%"$JR1����g��ZW�'��
�����54U8d��"��&��0�TR�pI`)��~�k9��Ь�RW쑛'����,�3�u5H�Y�[_Q�=�����л��}�3�Ʉ�ţ���qAv�'�X8)�^�� �.�gB�4XC�u���VU [�nH��*�!���!���x�oKk��Xv7�h�<��ئ@0��\<��0�X�C�t[#��p��d���Jx�w�9�%>'�a�8�1�=��'��n���7᚟�J�cxfi�NU�mm~e�����o�4s��� ��Y��_4g�%���&P>7�5�t��3��T�*K4�Rȶ�>̚��c4��Zs��̐�E"���1��-c�H����3�.
%�9�iE@ V�"�=Բ���n���W@%s-
��d���Ɉ[{hw�!"�l��U9Cq�ɐ����f�QM�L�qc]m�C����GҖ�.��q̅�"ഒ�rI�7���rt�����;M��D�CRA>X���ʓh���u�f�+��ݦD����ՖR�� �(B"��-	��@�.s��(>�W�m���3�[�'��j�]P~�Z�������3��4���Za�ѕN�f�q���1J��>{�	�,���F_��v�܎@��8<,���雳Ok+�R�ɣ�Bl�WN�gcy��8�I�|�����X"����t�&���Q���ò���(xN_�h'�"��I���;���ջ��ʞ�҇ꆓ����ֱoQ���CA���ARߪ�F�F��XD��I^���u��w:�߹鯬d%A�����~A��M?�M�")Nt(u����-�^UZ��52ŵd�<�w���[K�Nx&�p�O ݷ��;�^$"�Ϲ���� /��e���ex|�X��JO�'f�Z�٧BC
����F��z2^exiҦ��9e�L:ʃr�s�@H�y���Evdɼ)���x����[�nYАW�a9GaK��c�]���r(�3�iy�@/�맨kud���N(ԠNdΩo��Q�8PY�@a,Gy_ԽoY��G��a��``8�1Q��GD>�.q�����k��Zt��Gk�C�fUV*F��w�m
����y��]�������F<R>�D8}�׻�fD�w-c5�]"QXAe�$�2���oڟ�ѱ�'kB����K����NG��1v��<�J����������o\��c��X
w0��7��gSE��v�Sڰ�hu��`$R��o���N�~ۦ��"Z>�����Q��º0Ė�g�I?�$b�>�kW֪_�����l�ݭ[.��򼐡�|����S��?r�I���g��W�V�ӽr��fI��.1FoE����2�;#f��1� ��,#��>�2���*�(�X��}���9�4)b�\Ǚų�0��ԛA��Cщǉ�]����OY��aę����W�F�Q(_T�8l �V�2O�ߕ�$�x��X}`Y��h����ӫ�Q�'x�O8J.���������E������SXPl�T�[f;>�#��9�zB�ls:o:�?rSUY�c�߬c@3d�����G����5�W�t��җ>F�~�������*H}T�S�<a��^c�<ב��o��5a�	D�#�f�y$o������O�&��eM�<�H�w4p-/��﾿,����Ԑ�������W��9v�,�1w1i�*�G���Y7��VF�쭮5�~�K���k��C�c���Q���Db�}*W�ɊL�0�uw����d�s�`d�(�U ��p�E�mV�W+rVܗ.g�5t��	R���0�>쫑�ΗZ��q����5|����~������[�Y�^�=ܰ�j��h��.^���|O[���(�Ie��]��,��-���`��Y���Z�Y@9��%N�1� ���E�F�<�?����E���n�9@{��g�a!�0�?N�}�J!���(7���L+-�6�"Ή5'���3E�V�U�ү�Y���x熎��M���4S	���ظ��/c��X�=� ���0|[�����&�cX8J��1�)�]�F�á���[�&�����`��G����c9��P�F�w���giǮ�g�fDv�V��B!�c�%��v^���o4���b��#��Md�hԽWLͅ$b�A��;mr�_|�Ks���V�k5]n��(ʤ��zS�A��-~�}"f�x�ma�����#S�<5;��I���*R� �7EA�&�ybp�9���t.m�&nbN� �g�����$�v�^
�5��#`�g�)k�a�I�������w?�a�Ʋ�r7�u������.h���լ�hNB�'�׆jJ���n�h��X�k+Lf�Ǥ��说`C�����Pf�+�T��W�[ɃC����s@	�/�!vg�aq��p��$W��Ȅ�DI*I��H4��.�JW{ [΋@@]�������o9�	��lSÁ5���B� ��p�6;�㱳����;t/F�5�p�}N�v����VX��q�p�w/����H�~�tg�ʶ��J#�5r�:I@j��w����n�NN�e��l��\�Ƴ���0� �.�6�Y�3�?p��R��E��2f�P���S�_ndl�fٚK����I�5�-�����v�`j�]PJ�|����A!`/�I��r��L=��v�P�!����ہ��r{jz}kj~�:��8��F����WB�D
��5noI�!$ �,�b���Hy	�u�t>��|����*5S��9x����J��x��i<d����j�i\٨:�uB0~�7��V�r�[�B��c���Zg�
�Rye%_];w4%�k�Q�AfZ�0����� ����\��5]���J멷��62�����Ej���w܏�kG0
i�(�X��	3�Z���~&��%a�������^�łxkCm���3t�*&O�+r\�lr�l��Y)��Fh��uq��N����՗�o�/Κ@(ٙ6�[���\�������+��r�*�Ɓ��		#��~˴W3X��A0+W��7�gN��t�e��0�&���n���T�7�m�":���g������-2b�11�r�LX�}��7^F�&��f~,g(J[����3�8?L�}�.�F�
&�d�xn��5���x4�0F>�}dv�Y����:ݺ�*A���u�#�n�5sr1)a����$-SL%[��M9Ͳ�n��"�A��9�����W�9��O}���
7��V�ݜ���i�n�i�ߣFLd���z���d��B��|! 2�	8�$�p�M�w[��I	}e**&|_XͶ���E��V���T9����*%����צ ��E)^<MC�����dgq��%íT��k���l\�@�&m��J����D[qN
?�O6�� wؙb��l-){䅘T���
Gp�*�K����xߙ��˦�3y)�2y,z�qf�!�@��D�L?&�u��ˏ'��*L
�!/�/��W]����fQxm�X=^�eC	��$*�xU�_�J<���i�Q�r��0�������r[_O�ܚ���V�&����Ͱy�)����H���W0��\6��P��&>���\�٫��Ӥ�j��dn��5s�+u��>�BަO���H��iO��Y��tz�膬���v>�%n.�uNq|�=I]y����Z��0P:�>$���/O�������6�f(�)[b�r]�����|3��O?�ޗ��(��ge����<ԁ�$ 6j������ΰB��J;�d=f�e��B���S��"6�'�='�3�}����*~���F�3
p�&���/�R'G�`�`r�Z�_����Kr���|0Lu(1��ġ�Q��[�M�䁄*O��K�Űg�Ӽ�u 	�X����NE��H!����7�V�e��I�;� >맇ܩc�Z&�k�E�
X��P�Yk�Mp:R��<���8
���R7���W�y�ȦE.�W*��F�v�6D�l�
MC���I��f�-?V$�ѿ��<;����`���OÓ�T�h*~���C�w'
 ��9A� r���'�]xY#�j�C_�!�&:u�E�F�kD���ky����O���Ae5��<UހV��(M'g{ZE�s���#���v���y�^ú�	'0V˟���|���";�<?L�B��KT�� d�X�}>���ֺ0KgL���n�t	;��/�VdG�o D����
���So�ƃ��?n�,d�����-��|�&E�y�*����Q��e?j����Ю����^��l>�c���Rp��*�����!)j�V����!������]�,9F�њđ�����W��@�%�+|u�y��wQ@_�H<�s��[�B���T����I���9��V�<7Tw��t5���G���3>$�ӏ|�ǤmP�7Ot�]��>�߇�b=�������\0��G���H�$#L���艭Gɽ��.�SI�&��`��6��P�?3(���K㗉&)��Pyf�����52���<�ɮk�y��V�ʟ�ύ�o�<v&�Gۍ3j+Iq؆����������O~wX�!�|�����뼭$��3m`�mR��	U���p�S�N�v��0�	��ƈ���#,
��2�>���̀������.x�J�FDTϺ`��(1�0ʐ�w?L	�-ڈ͔��Mǖ��B<~�lH����<��f3�F�u� \JK��,���J�e���}��6�>_�K�ya��` ���7$H=���s8�1O������JN� �HP���H;DJ������JO�q���$Ǩu�%�>�6��|���Z��n�z �ث\ŽJ���`�z�<o>B}"�_�%�N�X����#��\����W��̣z�P�.��":0��������o-���W$�
������HV@ϘU��|I�Sx��Al�qb�9�(������D�N��d��w�<q��~��o���1�mee!zD(�C}0��a`�ܘ��dA�&�&_�F��+X~K��ۻmX��v��_+>=��~��מFN=m%����������a|��NU��U�:�S�R�k3�.F�ku���Y�j��j���Ka�l{�*��B�R�.�h[��x݄js�=��D6�#�ރD�Hjȃ�ɉ~�m�&s�{�Q�;���L"�Ӿ�QԉL������<�ϓ@��m�;>I���nT�l��m�nZ�ԭ*D��ɤ����;�e1~�M ��R(�D��U#�`������Vh]^�\�*����6�9R��?�E>k��(����1���'�+]�>3:?/����y��py�f����O��(�2=����z$��ȑ�Jv�)ōΞ��n�Շ输Se!������}�3�Aݎg�sr��� �o�߰��a�úȊ��s�Q�ѶC�M0?��Wߜƍ9�i�9�yR�P���T���>�P�WF»��<����P�Քن&PsME)O�Y���a���Q�c5a��xN넄��2	��wt�e�qO�S�Ȣ�_�5�#z���7g���)��L��H�P���ةh!\��nŜEِJ��=^@v��:�66������g����W�J��7i��`]a��5q���TeV^W�����r�9�s��Gu��ٗ�:�$Ql�Hεr�DB�7X����1�}qr�{<�}y���>Y~H6������M�?Y���I2Effbeu`b�H#M���V<bD�NY�_A�4x�����#���%�o�0��S�����iƻv��*�9R�H3o`4���ˆq��Xw��?8S�C�
�����E�-�ZKg�I�Zm>j^�}��H�`�wl�N`'��)R�O�)�;��JI:6N/�:|��S�.N���x�d.5sǔ[5�8p��ߞ�}�����{D���kG$��X��q$	��j�?Dt��N�� �P1�V>���.��EY4�Ƶ�y ��-���0>UG�}MK��v+r��~`6���,��V��y�?V��1�� �7P�O�91%��V�` ��wg��"�N�F�d��f9qe�'W7�3<���A��_��W�`�o�Q�R/8����iOV`��+3^i.������A��#��F�{8��u�h�� ϸR��͑����@k�]a5v���8�}�ekx�q0��}��=�s�%搆)ZP�v_�[Pb�!i�{'k����5�2�2�KW0�ae��k�[,;o��M���Y; �(��`=��7W���nػ�7Jl���n�Τ����_�!f��,����BW�>XS�1\����Xl��������A��?�I��k�Q��4JZ��>���_�*�]����mP�"d�!.�ۓ}0�j<'��%ȃ���)*��=]K����6�����>;M� nH���ń-�{8[ӄ��교s)�!9q��M�t��>���L��
D��f$��l����m�s�Y�s�9�˩�
�X����@I ����S#���De��hh܍
*d�a����P�L��T�NAs-p���dm�Ҧ!���(愔9���Z��ӏ����x� _G���Y��YRk��f�TsߋS���fڶ��˥
<� g�b�ީt�l�"d��Dǳ,*Rw�aF�<܅E%΍+!������S���� #�'?f����c�/9�k���(��I��BlFh)�K����.�����_�A��M Z#�Fn�W��]
!o'ڝ)n8ؒ�d�%��n�m��,��k,��c]����Ofɗ�Rt��@O_�����p��S�v��b����	Kef^��\`�&ս��1Bx� ��=9��������l�\�po7}냓���X�J���?�-O����<9�6r�󩎰���:�2�	$��Xܵ��(U&� ��ދ�B�?���$�^C�c��x���4?z'G	0�݊n<͇��� X}w�6��@f1L�߈m��,��{`%�����|eE3��|_<i����E����C�d����YB@���N���=2�l$�L}j�v��fF�A���"��A
��v[qAS>��?u�58*�&�i�AN����BE�{Lڝ�Y�e̩�Ɇ:�D<kK�8���\��[��O�N��ʀ^ ��Dn�@��e9k��o��QB�?�/tK�B�l{�c��|����*���0$��:�`;�-!��ϸ��l8I�>+"�����)��ߨ<�Q�s�d�Ζߌ)|
��}���ȗC5w��t���>%�q,�|�ᚧ��ָ�,��XA!.��,0�;Mi�.����^F�a+�K1����A����BEd���s�7���F��k���� Ǥ���z��S�UL�9� ꎖt�#�y;?UE<�;(ϡ�(���ȏҐ#Z��ᩌ������l�X#<Q���1wx�|h��ը2�"8��aAq����-pk�zb�3���"��*��?>�H�gk��@�y7�X�D��L�X��.�B��W��#½G���Ρ����H�3�!FyE�jƦ~ga��6�r�/
���;ۃ��Q���3x_��#�f�0��N��*�`W����h_�E$D\��#[���2�������-o�^F�\M�䉍�̯"iZ����ʦI;��SqEDj�X
E��Y{��L�w�>������������c�0:p��$
��):��|��.��f�+x�ԧ&�ӾfL���p� �a����j� ����x�w/�vw���\���@�K5t�jF�~��MٮБ��mӕ
�
fs����!i�H���k`�yZ�ab��ц�CϜ�)C��e�V׮L�HhU'����
��[N�.6�X󲠱���l�	��O�]�bh<x��J9���ž��{���d�EO�.GR��j+�Fp����ږXd`�9Qh�P�G�r-3[8�2
�e��m�q�e
�Ī���[��o�5�\/�M��$ݾ�s���,w����V>l�S�d~g�X�"�ܼ��Xf�7���d�α�����G�ˋ2�K�HDh`����(�@������7pj}��:L��3�{���F�Z��hG�\`�+�*j�\i�Pg�Żg���F"���,Ӕ�Q�d��9Ah�i(�sO	���4�	FW�nq e�j��<"]��O���?'wd�������5Ӻ:y�`h�L�nh��/e�5-v�ȃd���L���Ø�wvY~�]����ת�] pT�̀�"��.��#a�E����  V����]���2��W�>�t^?�9������-̻`t�9�ǭ#)�N���2Y'ȱ+~R!�X�,�TW����(/]�(�𖂞�}Z�)Y�n2��-���c�ޣ@������tWv?�ط"J�|+�K�m��ڽ�vȒ#�����e[4�s�L���'I&적W�ćB`�!�ƴKF�y�4��;�W�c)����'5�G�����q�z�!->��T�����-q��i=�[w�ſ4�/>h��Yy3Z%0����e�2X7kJ�7|_F��l ��%��oO����4�ڤg��/�A�EN����c�7�)X�NO��dF����<uA��[��D�>�C����51����z/p71 ��c��F�v���rp�])�����n�q�OA�Yk�c2l�1�i7uw��|��� ���t S̳�!2� �ޥ����<o�\��g�N����5�Pj��Y��Ԫ�F@ �Q�c���C�Ǿ3�.�������ņ9M�)7@�и	���.V��6�A��Y��H����Bdb����G;h��86K�]�H�h�t�8��7�+�`N]6<�03�;�|�䲹��<Ƙ��#�E�E1.Ff�bU|V^H|�[l�Z�f{����b-�;��w��Յ(�/x���6�W-��5+qn���,ح��Ё�m�	��{�|�>�@����&�$Ir�������@l�E����@Ms3���� Aɒ,�3�:U��&S�(m�m��jK6���|xLw��Qd?�j�gWAuBW�\�l�H�FN�)���$8���I#�R����L.�@,�Ё���!��ZrF�3l�VڮND��5y����m��O���2�f�J�癢����#*B8^�[	�=�R:�Ӣ��b���1��.�1w�
�c���4bx.#%����Ƶ��_[}���\�� ����
��&9u�nv_GJ�bR���;�l�� ��)ߏͬU����L�Y�#�~��.�.`o��-���z���P�/s���؉�v^��{��7�j������K�89��i��q:��z�f$�	���(ŝƭϥ��3�<��p���>2uh����н�T�Q�ܩ!b��}��֒�tmC�5���HW��o��P,�a�@+o��x ��}��]��?�gl x�O:.��o���3c��Ī�޵���$U~�."X K_Y�b+X^�3��u�+�~ P��V���3]J��q�V�3�(u"@����\�h��m���
��~ο���o�a*y�A�-r{ھ�'�\Y�5_���[6�
���u@��nUYK �3�^��^
�V���tF���Y3C{I�U��^X�i/��~^P��sv�ܾ��>�#v��k}���k�{{٫No�����G���m?��c�=<���*$���f��=>������~�K�n=�@�!�{[e#��Qc�ø�9nS���+4�L���������W �#�i%���>��5�>�[����j*C�y�%��pҶ�SD�O�$gm�ދ1��_T�ݬx���PyWt=�'�u�:�ӝ;�8]��G^JT�/o��
�����44 ��:_���I�~���T�yӃ*��?}ɘ�}�t2�������CWm����g
�k�ǵ����i���Қ��̫*�6�7$DH�BC� �i�5Y/P2d�	�AZ.n���\�lِg�3\����t>��\�>z�~�#\�,T}�$����(x��T{�,Z�Cz70v4��āq��,9걸v�Uk��V��c{���*�1��uɐ��.���'�Z<���K���W��V�]��_��-w�g�y�G��Aׁ�+7�{�4/x/-G��@�Q�<����b��4!r&�� �dď���˨g�4/ԭ�mOh��+"_w)��9�)�,1\��i�ߟ͑�w�����>�:�.Q�p�Cݺ����u��Z�i�����c�k�*{R�t���W���Ed�#���4	�Dݤ*��榝De� x}V�G{{�v��Ԃ7&p�f2P�Oڂ���t���⣝$���C��	�2MA��~R����uz(�J87�S�,�N��3����Z����rW�_�Q~�YkjA=b��$n{��e��N_�:l�3K�jt�>�X�U�����3,a�	��F��lO��mujr�<l�.���f��ʪ���h(�i���M忚���Y�1b�x]����m�צ������OgR�ρ������w=��Bb�ȢU��p�s�Bg��a�?���d�n�L�#�,�"�ԗ�zU��D]O�="<�f 
��0�Ӹ`�Tjh�'a��N��X�TjQo�ce�Ż�Yb�ͬ�����|�����Ӓ��$E�����e2v�i�7#����o$e�FO%{HZ0��E�;�+��px䉏M�f�3� �~���k���y<Q$]��J����GI����̜�7�\�d��PlcRP��$<@��ؒ�O������$��Fo�jy�[�lqu#C3r���hp�[c�Zo�
�`�y9?�CW�q���-��@`�Xy��@�t뀌����LU�	�E�5�/�o1x���Y��3Q�u�e���(D�����a��+��{�1S?�D�cC\��<�� �K�T�1~bj��֥v�ڌ�濠�?�B@W�WI+WIg��{��iʍA�c3Z8�`+�!����ů�.i�����:{���'�A�EŮ��>������=���=B��Q=��R,+��x���##��-�c��A�{��u���Ll�-�-_�_a��I�*
!���w�O^�ɫ��k��,K�h����#.��9�V4K�ыZ�k�ƾ�PNi`�Kdw��%��3f(�M�3���|��T� ��Sz��euO9<�fIY�Kې�D�5z��ihu�yhf�NF(�V�������M�߳��ة��;�`��=_�o��a�b�E�X}�B����Ճ��b�1ɬCo���V���|I^�ۤ��B��:ju�o��8��Oܰ�H�_�1��"!/�OD�nϘm�5��0���^+
������;����/�">���葮u���6����~N�.�^i��Z�0P���Y�"(��{�����l��r�1%O�{������VB��^���7�E��6�^�酔��<L�ؗ���e�z������d_b���H�}�-)�_~�6F��;K�G$O|W��ߒ��z/���G	IC�a��N���>����t����2�oD�܆T�"H��:���ЅΑ�x�ׂ���p0E��.ue���:�N]<d�&M��q.R�B�(cWm���'!%Y]Б�`��BNn��M�۸�ל���=�ay��M��q{�%�wY9k��>&!�Q�j+�e����w?�zKςA�B��9!��h�#�_��+�͞��֜y �IС*��S+��76�+̕c�@�`�-M\���(�χ��̹��P5@�Bv�kL�"��P+a&�3��� �:�-8��s�~pu��Q����렌~)���Տ��,���б�x�d�� ������P��Y�C)q�T�@K���*:W�+�E��k�9Y�
J�D+��=QT�'����▔��*C~���8���P������?� ���`c$7��96�r_w�
��슮�s��������C�K-�k�P@dS�� ��"3�z�y�A�[�b������)�?��ן�K�>>�Q��Ez�cw��Tw	�L�� d]����x�z6"@���!���5�G���;2���~_�[����kC���/JP�Z����5QK��mU��T<'�fE��qx�����<7���5�5̕㻷�Mt��+�n�g�>K�L��}�r���Ҳӂa%O���d~0QC���:���J�hć,.�EZ�]��O5�������M%����! &��I�����ׇϫΔ�����.��[ 3�`��׬����ɥ̶	�<ӐI�C,�:'�B��3�"͏��s��\J\eL�j$l�qh:I[��,���R
B��ic9�e����dU���3������΍���5� EƷ2v�;a=+����#K]�?+��	y8Ŗ��Mb"
��ȴ�8�aҿ]�Z����9/"<�ݼ�.?���K�pu� ��pV��Ƞ�2�+�}����6Lt����{"�+	6�@�)���(���'���ĜT��v�L;�ՙ8 h�����G���)��9�]rK�V7�P嚲	���M&]��[Y�վ����m/Ɂ3"}Z��!���1�q�8y��1��G��؏F�6��x|�N\��'C'�tY��*"�%�yt�L��%�eT����G�F&��&X�zr���˳zu7���P"�`p�����V�ZI<���I}2�dW}E�Nkf�E&3�B���6jN{�%�O���~�a�PU5�:�k�"�^�b=n\+a�la�0�q�a"Yk����cU85�7d��Э��d8��ϬD1<1X�@}J��d�D��/^��D�2�ūT�wM\�5Ԩ�<�X��j>�ҽ��+Щ0��㱈�ԹF2�j!wg	_���nX0�F^�RB��T�ɍ(_"�L�[6��x��P������k>�s��z�Z������F�I^�ϲ��&�}���p�k~\��Y�!�-Q&��{Vx�ǘ��t.��e����)Ws�7���=nG�_/�P����4�jvF[9�ɐ������&9O� T�{#ѻt(&'�gIj6�2q�Z����,�`���'�eD;�Q�/��!���ۜ�[�nD+�J�!�9Ω��J�����gů���i��)����	��n7}�UL;�<lb�	�~�m?u�鯧��5Uc~�eyj	=��&e�YW1��ñZ�����p+GM�rnk�ώ�"�$�e$��%3^d!@��_�(���-�I�2�i��N��d���:�DLh�ܩ�M���#��[�F�t�|(�ZY��PG�)ZMH��%��;�HE|D�����P&@����^�j�j6��q�z.B��-�����"j���)s勎���T��A_;-�C�~`r��m!���@JЭ��z$כ�j(骏��ޖ�n�u��g��o����Er-�e3H@��&�C�±����$��lk�G(�<�6H��B��Z�
�i(�(�k��O`O_Z���Lg�?W����T�H�� x98b���$���0 ;�FM������10��I4x����O,,�x�|#+��g�	���	f[�M6mÐ�k�K��5[���Brh�i��jεKEHKj�g��֫�۠m��q�җ�+�4� w�W��Ě-�U�%X�q��h��h���{�i���yu��\$�������]'�t��Ԡ�O�&��n%�wQ"	0e��/f ��%���Cν�s��D��g)$X1�:�G
$D�QF��RXJ ��b���w�>^���#=��*T�[)�"���~�;� lB-�"�jx���Zp��d Qy�`���:������C���k+�C��U�@��?BY�w�E�Y�q%j�[{�wr���U-������k�]��`�N/����Y���'C�>�Nz���=�B\z�Z��@�9)�G��u�-��a�t�s���������8��7ӏn ���W���b7��V� �9��f���O��#NT
C��v����3�[�g6b��fD�t�z�k��2?�����+�v$)�Y.����D Q�7�H_�P}�������*Y�J�MM����A�͒��� ]�
�M��(p`k(/:�������%���9���k�}�C+��wɡR��w�cZ����c웚���dw<��zw��Y1��ɣ�ӭ�M̉4xT{�rv4��=ˮV�}R����qbTϛ7V���1I��[숩Qgu^u��1�^��tot˽�\e���};��H��A�QH�!Z�\�T����	a�p�^S�R�n��f�U^��ʰ��q�H��9�����ǌ��S�I����>k�kF��@�fL��B�/����٪ ~�=E����: ��7��e�/�R��6>^�ŋa(z�V��)x�b����CE�+�>�D@�Ց�T��u�f�G���T(�g���E?����Q]l�P|�ߊ'1()�h�w!'4�G���ۨ��^|k�Y[bz�N2P�G�YT��;r	�n�r���b�2�k��޷?SW0���41o�D��F�F���tf���M�%�(]O���~	�^�c���s�yQ�~C�{��됢p�}�1U��0 ��V�7�'jˉX�5�t::0�x��TN�"ߧV-,i=EL��:Sޱ@�>�H���� e���LK9��t<N�#+�ﲠ<[��mW|�������r�S�ڐ�ɕʿ��a���SO��N�+�����/�>ٴ)�EZ1�*G�#�M5*n����<��ㄻN��9OK>_�м���þ�մ�%t�b�z|�}����iT�~0�iˍ�^�k�\O�%�$+9��tpp�+6e�>�<�U:
����̲]J��ެ�����t���á�De��/���|@p��3\�˩Hak�<'`J6'��\�furga�풞/.���o��S��u�ϣu�����D�tS�������S���_A%��w�5�zEŭ��6�����;�)l��S\�n�0��b����T��F������;`��%:��������0ۿ��JqVNv�j�7�e�\��R�83�����0�
��� h��i�x�k�Y��9a�Wkh���<���Z��8��6�},د�kc4x#rŰ
�t�MSe�P�~b�V..�W���@�̚�h��|=|�yGH=��F�!����������e"O7�,�J�i�ckG wMUU�����u�Z��<�)�/���I /X����a���?� >fذ:Z�!�~d��YeG����;��PP��O��ؓD���_B����w�lN-��!V�hkw�� `w|K������J`� ���{R�����%Ɨ����y�XB�J2�H �E����zٜınD��#Ec�5qX��t�\~w��e���)u�Wk0�L��m�6;�Z2ǣM�d��Ome�׽$�Ec�ZGZ�%?p9$E1�W�M�����c\>	��.o�����<���Q����f��h��t�`�qϿ�y��9��9���~�GD�ː}y����]�E(xGݣ�~�9{���^��N���?�F�=�}�V7��#�"����xB�ǜ{T����	�d*V�Z����YtX��_G�ٱ�6�)3��"�W$��Me��S�W�)QE�-hCh09m��gb�љ�9!±(�t��kn���n��6�s�K�.��p>��:���/�3�K��0
x�BD��Z�4$Zim�4#�zW�p��>�����,�}�T��OI��6.��I�+Nw�[}����B8��ݗ�1R���(ď��/A;���4<��Q� ?�.z��ϦÂ
I�8)�`OO;?d;�2���,����2��eE�ٌ�'��c�l�V��g>��k9�������޶:�w�h���������H���� ڞ뮋�$A}n�B�R�br����щ�Crý��j�h8M��h�Z��G����)#�/5��
��Z�e�~�*5����GN�ꍄZg��TS��>EY�D���������q��=r��sxyd�Ti���g�\G�'/a�GЫ�-�Vta��ڀ,:���)����H.#�����dk�������ٳAn�/y9�ɪ$�����~��)V%��yBpaC1^��b0��#F�X���fu歮���� ���\�����]f�'js}1�5�mxo��|�X��n"�,o� ��6&�>�Z~j�m#?7xF�^��"�'�'k�pjȯ�]+Cc(E�}���Ze�5a�����ه�I�O�����k��P���x��{wu	 �h+4��~�ˢ�Pm�%�[��rU��b�}�]��C�PI��	܍�P֙�v�4���A� ��&Rh���3��i$d H83�輩����!оӴjG�X��ϙE��!m�Fj#��$ا�Z��U��gQ��p;�ҋ�苩��V���/r�3h3J�|�DZ��浴�W�P�0Lw����6S�V�(�8��:��F�dR]�n����UV*������Ok��3Y�%���>�u����� y_��[����6	��;�Ndђ���Ɣm�о��DrG���=��O�Ԕ���0L�2"��x���;D�o�T�P���2�?s-�VV)|��ҿ�wIm�A(S�uS�ɼ�&��?�@*�g�ѝ(5�&@�;���,��-�xl���߿��H�Xn�����X@��=�Mcpx�ʈ�O̿����Qy&O��D!>2�7�a���a�:�_�*=њ�7�$(�Z|bӧE�=K�7h�`�OP���Wi��-�`��\vJ3�Z�l
?����K�XBAov��oyC%
zNʔ�O�6̮�ڸ����p:'t�қ�/�J����.���fz6��}�V��!�^Gɾ���u$$��]���qL�@D+��AE�����Y>Z3�r5t�^
�=Z�{�%�;��s/mm�Y��d���qQ
��5����i���^�t�o���(�G�f&|�I��Wλ���r��\��F	����������Լ�}��@��w0#"���b���s"��~���E-`�ϖ���ZQ	h�b���`(ρB�<,������E�WÒ���_�
ۅZ�_đ^X�<]�b�O��nM���=����i�&XN-_�ĸ��KֽŸ���J>m�dwf��Mtm sWU��}nud��|�������3b�a�#⑭��U�K2�y�T�o��������C7�M�K������ �G��h���c��Q�+�$�s�hLqUZU�ӄ�r:0CRj�|��y~�&4'����`gK�;(P�F�*��H�&L����b�3�_mŠ0�`o8���Z�I1�r��p�{U]������%���F��/�i���'T`�����+r�v����#a�c�$D?Գ<������>���U�.A���\�����Q���]U5���7��l�Q�ι�$)r���(Դ����4@��qH��p�m�&��\�{ئ�u'm�54�}�Ѝa5�Dm@q'���=\����=e��}��ğ���l�X�|�/=]X�c�:"���<s�k����b%���7b��t�G;K"���bH@>;Q��yZM2��P?��c�P��N�	$( ���£ײM�a8����2	_�f@����mB`��x�p�ሼ�W�>�L�#s@KP�����[x����v�o�-�:Fq�����f�낳\�� ��`���<7}Zp���ߖK�M�F
KK�`�W�#�Lu<���|w��ȐA.6��Ƒb��x��=��Ҩ�r�Q9�R��?y��E���L�^߫��������4��W�3W�_����Y���͍���{v1��`����nIx��+�e�/��rM�6Wg?}zt��(��`FE8W��w�L�)>�x�+��Fь������P�{��