��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>�;�Í�|>�qT��>�[3�W�ry�cˀ�
��$� A!�J��^4�<��(o ��ڞ�yW�����ķn���_.���)+� *: �N-\�z*R��h@�e!Q9
�}oWio���r����m�顖<.��J܃���b|>�c���x5Q�>�����bN�6�{>
�h
�F�u2ӊ�h�Μ�2,��ւ3��Xp�Y��z���u�{Ƌv���NVu���(�J�GыM�R~�՞�1Jf]^�V1[�\a�yJ�:Q�$�[��E�����-E��H˽W$�.�>��u�l�0�&��~J�	�������r��l=�ۧ��l:���{F��)��j�Ĉ�c5��1Na�� ��j��h���dm^�#�e��
+iX��C�/s��8]A6��l�r��V%	z޻ �*�n��`�QT]�/Ʃ>{>7m��M҈$n\�j����,_D6�~��w1:)9�a��Y,T�i��H�q'<`#I]�^O����<#���afK
M��Zm����2�L0���'�� m��E�Xw�GN�1Uw�Q:Ġ&p�	����<��<s����m�f�����3:&�eϏn&䄵i(X��[��ڴA*7@_.��!fʔ`�02U�wfͭ8kirqe-A {+�����s-��)��=D�Pk�}⤕hv=D� &`�{�����k��6�J���9$�&�>�6��a#�ڡ�u��t�jAZ����!
g-B�(�`�|������3(:�*ߏ�z��EѼ��q�8�܅�_Ak�P�	8�D���OsjZ3�5�t��4��)f�/0���&����`�Y������Z��AO�bD�T����"S(�2��8vOmnbW�K'�<�S��Τ+61���)/v@ z>�J}}]�����7��4'OK�^�.9.0�v� �-�ȗ�� �H����$h��E�u�n�f
��+�7���)��<�3u<��)�-�7�f�F��Q&ש��jٗ�L1i�Lf8�A��'��G�KI}�a��O����KA���@qz��-��������E��%Z�}���b����~q�#:O�?�]�zil�_�����YGڄ���Eɂ���Q���u݂)�)L�/;�oQ�*ǳA)�{D���q�\�|g|V��I��`koQ�8��b25rv#z�T�۷��.\�24ֹ!w��գ�h��K�\��|��֋�F��7W�����Չ�C�� J �C�I� ��}F�?��Yi��O-��v�: 8�p�v����~F/�������!��٧�܇(�)��d����Гޒ�o�}=�^�?Lyΐ�`��-�]�$���pJ�&��Ɇ��ԥ	{i��T�x��B@���zNN��f�7��h.�i%�=-W�i������5�K�� �o$C�e�4X������
H���"�EtC�����zP�a�K��~��욹�B\}ϙ!���]�H���k��^��d����g����`��p�&�%��#�{%��G���!T<���J�N���EV-�ҩ+�"5�a*�p��7f�޾Z�x�t�ܓe�0�X�w��R9D�=�Y�g?ހ`VH�|Ś��^fL��ö�Q�.��ӻ<�fȺ9�Z#���'��8��Б��㪍�����UV�`z��M�Wd��mgl|����2c��8�gztƹJ=��b��`��U�p�<�^}���[���"{<^+�ޤ�B�"g�}[� ��:,���n�G���i2�����{��ğ�.J�D�U}�q�'B��&l�̉�ѼQ/�@<a�#��t���#r�)4]%IpX��4Y�N�=�~���AG��^�Xzf�0X�O�`��UV���� DP=ZAcsBI1��jiF�Nz;�=��2Q����ryS*̫2;�*�@�ҀW�lK���`�� �RxG������$���-�yDW��	\��v=�o�W���Ù`��eR. �q�DH�J��4[!�R7i������Э.-�LDb�g�7mN,^^׹S8�<���8/�P�@�*����>Jǿ���Ձ�؜V \�4/|x�cm��_�����t���E7����Ѷ�+�>$�L?�s��#�<�DJ��Y6L��(6�Y˾*�f���+J�s�힑K�����䗴�4ϏO�{pʡ�&�*�v	Fa`��?�8p�j��4�R���/��q �"TB8(*&g��i�Btbu�~��=�^БOX�r]9�� ,��dfk�W�`f�ј-*@g5K��a���$�C*��z|{�#ZZ�"�$�LA- y�	(,6k�|���=)?C��e4D'�(�<DAn��G���+���Uo�.��w��	��ݙ�q� Z�%�b0����ҐI�e�
A�Q��^�J�j:@Z���u���_�*���.N�JЁ���$./�Ix���Ĩ�(�!��~������A1 �ө�9~Bf䀴�"��p��	�A�r���!j�Y�{7n��dY�T��`i����������\s5e��b���01T챈�-�e�K��P�(�#Yq-Z���&��\��%��`3�n8��Y!��V6��}Y�����y�]+���-y5lQ�9�>H��V
��_H���\�L�@��jY]�N6����d���A;�l/ka���y�G�3���y��ofy
�.�D�� m;��)zp���y�5�pL�.�/Τ�)�p�|M�Z!�/{%�C>��n�Q|˾G�~�uأ��?�nX�鎈�R����isP�-�i����B��
�5��a#D�ސ���،�Vu�P�ʖ�p�9�s���!TJܗ O�
r�������� �+�E!�JA�+����m�l��2�i�T1�� 0t��1u9nމ��%r
a� ����B
�F<y�]��
�%�a��'ԃ��������G:�@�Ѝ�+�bj�`��-^�{D8ָb_�C�@�1-:��W�{7<��z�D��͠`֑��jä!  �f��?k�R��?�\|��z�"ǹ�H�Ԡ&�����m\'�@	dL��s��A<����n![��M����#k�y����r#�G�;ٰ�F��RZl���`�����ۡ�.����*圢]�$GAܳO��Ai��[.�U�us�|9^��3��d�5�����a~��߳J>����<ldI���RDZ ��eY�[����Q�<�g[n�I(�7ܫu�)���.R��G����\1����H����o)����Hk���������~��W�����p�4�{��r���x��U��c���3S��d@���6N�K�3����s7�����ջ�a��9���a#�M�pGY#�Q�%���C,�`��|$�d�Y�V��_�ja^Xթ�>��h�$ǞIv��Բ� ��6����`�E���t5VǸ����1������ϘWv�9�U��Ҥ��f��~�pB�#��ܖi��� �,�oh��+4wݩqQ����x-�ѡ��	��i�q�Ӽ��#[~�FR�j͟B� �w����MIkha,POM�f� �ϓ�`�<b?���8�x*���\��b�u����o�_�3h��7��u{T~Ɂ��%0o���c�z�j*uf��7�^L��MZ�,���j����o���3�y%!�Y�S�z��Bx܅��\��Хʱ���� E���Q��Q@B+-nY�'���y�3��H�A@m�M��!,O���p{����ę&�iLe��f/Q��l��E�� Z�����t�,�b�΋�2B{̾�h�wK^ޞ�Bqvq���E���P3\t�7)��8�Og��~h|g g�����Կ�`�Ƙ�휱�����?wz���