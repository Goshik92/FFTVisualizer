��/  �ŉ�䗗�[dw�'T^��s1T��MrNb�x�>�l�&i�e�����ֽ	�<���%��-���]��s�c%����2�G�:$�uT�k��8��g+78�'���û�t���6�45k4�c�{�U��.�ƈl�T�o&�C|$��UGXn�W�^K�.#�訆2U�X=�ߍܶ� ܚJ��\�H�Ř��# �?���q{@B>8t�T��}��ӡ��[��ߞ� I��^�W᫐����k�SŪ�L}�\e��!WV�!{����"�W���W���O�v"��d��|Ѻ+�$t��>W��©<+���jT����sq$�tc�t�
x��f���p/�2���5{p;�$uCb&�N��q+h_U8#C�,)N�S[�r(>��`HX����5a8Sjf\�|Vv �|�
���ۧwѸB�;Q�)�q�ǥ̥N�y�7x�S���1+��Aҏk�A�hg�S����	�㳰SC�����Ylj�;��Ɉ/yl�Xь�}G�X؊����;�'��VG^:0�y��F�	���D�:j�k̷��u��F'U��X��ù-�h��b`f����#0.�w�N�st&C��Z�V���!: ���X���h��.�u7x/���,��� e�����엙,�Ѳ0������)��������in��&�y���F&�:������q�q���y
9���`�}��f��9�'S}�@ 5�U{�]3O:���[��x�+U���~�v�_}v)�>��
��%����:yxjD��B6���P^-��T�/{i�M�;�X#���"_lAMP���8'����e���d�X_����"�D[䄩�^�3�J���SY!��qq~�����T다�|�d�*�d��m��c:�n��^�+����=^6�zٳ`�H&`���5�[��t�f�o��o���LO-�Cم�_ρA�plX�vV]d� �710�6�')ߤ{޷7]��W��v��b����]ᨔ�3e�67�᱊t��V�V2��t�,��-�L��LM���4�+���f� �~�6�%	���9�NM�8�$/�^ږ��8ܛ��#K�tZ���	a�C�67�T�^JO���rB�M�$�^K��O�==�Dg��9g䴽�ԧ�3A��k�T�<�v��;*O��)\Y�p��]�c(��1a�����dPǛ�I�B���ώO�(艤�3�ão~k����\���~4���J�����)��55�&X�=���2��.��܇Keȭ~��[y=<��N���9R?>oȖ"��2(�f�!�8�L����w	�k�$��&�Q��j�&!`��&��fN��벌;���V{Į�x<���:��z9LK+���1��h,z8-GxIS�	�響�-AX�M]}�u)#�4T{�����â����_|�$͓~(�>����㴧���N�`d�II�m�,��G��Y�8E���'���.��n8�?��\4	˙�䧄Ͼ8�m�Z'2�C�.}UQ��]������$���_M�P�;��,&��[O��t*@R���ѿ;���I֤��ާ$�Œ��u?�B���w�I���&`�Wh�L;I���mc�>Z�W)��:��@��!�,�1�hVU{�d*�#�%��CV?�»�WD\DJA8(�ٛ�`�y�k�+Μ��!��GrI;]:Q�cԱr��=CH��C�����.��KVʎ%�^i��ls��2����yN�P��-ӧ7:�g%6�$��
���c�FG�K�k�/�|���F�g:�i���j^�f�~�k:L�Z��p8�J ��n����ewҙu���ݠ�'��=]�n@F�k�)*O&���!E
��W����b�ze!����SK��n8}�#�=�d�>�䳸�A���'=�NF�����3g���b�����q�@���;N�7��N�:����@OfH�LLb0h�;�!R���[�U��
��x��R����� �l�<d�!�,� s���MT��S�6���edd,��}��?B|�6�~�Z5�I|����ϵ���ϡ�:�Q��
�q�j�W"��7�^M��0���S2Pc�嘕~��|l�T��E$��j L;�l��2:�B@�ȠT���6�В�2[Ψ�:�O����6m0{�,sp�-1�ͻo��u��@��]��2gR7�Ds�s�n�[SL)��#��|L%�py$1Q�#��A,��X+�|��m��I�ˀ�K?*x�m�/2�x�<+�/i7T�)@�Zv��j���`��Z��7��q��� `ｱ���$C��ܩܐ�������T��a���������Ң1�h�l��%�O��$� �$C��S5c!�]@Ue��Պ,��y,:'���`��=���lo�2f�+����Jc�F	ښ[R�-�Bx<�$D��XY
�6�4�I����2�u>av<	P2���7o?
z
��7��w�@�/�����(D�A�s�[=D�;۫y2!��Yo�v��$��8�ȅ\�FP\��M:!^�in���z&}�����R'��^UP����~���ekPɗ|T
w�D�Y5��M��@e���7-�rN#g��
Y�\+���r�7?c란�t��j+�eew�<�@*{\�0N��Wa�iX�r�&]{f2�y����3���c��s0,���_�����V�39O1���`�c>l�����!}Gݺ��7�n�Y�Jur�{Šɡ}�������"�.�|�?�I}A�8���*�K�+����I�Ҝ:Y;$�R8��]��k2}��rp_?[�. '�-:L���tc��;^�6]R�̉B7­�2?y��2^�w��c�׋��U�O6��k)BoQ3�\���ǎ��p&�s'�+;ZK�,�,uɃ;��� Kk��y�Ѹ3�D�p���a��/m/�^J���Ӡ����G�3촬��G-����.�M�k���-�ZK����YCC�aY�׈>d�~�����<6n����)�f��+��Y!��X��k�\+��ﲻm����O͂�a�+��c󑯒��$�n��������Mt����[��^��ø�����f.ٙ�N7
s#�k4��ا5H�N�)��J΍j��v�� �{�`A�z��� тNXh�GU��k�h�Ԝ��G�	�ܟd��e��<���|���� �ʸ�$�n��),@�ҝF��l�ć�Q�og��K��
��VE�Kr������T�%�V���Dr8��S�=*!/m����c�XAȐ��ɞ�#_5�g˃��2֮�����Ӆ�i����s��+٠��S�3�%n��F�M����v_��m
��<�1пS]<�r;��q�8���{�nU�*�/Oҝσ��Z��=�`S��m��DuY���P�qz�x ߬^�<ѥ��Q'��O����Y�Yy5����q�<B���[�t���<'*�����T��2��_|�)ty�9�-i����\X��?�N��2�kY�}��(��uQ}�j�e��fٵ��x�<�����F�Շ���u�g�#��oǇ/�����j�n�q�4�\0`���e��wzݼ>{�W�ʖĲ����9�� %S$���2F��B$������k�*c� ��TȻ��o�� ���Q��=RG%����/�}��LG�*&�?����b���{.
���v]BewЂ�@L��m���\�ڧU?ʽai=A^���^w�(��\>�h&o�(��qנ)Wb�����	��q������T�'k�	�ч�" �B�I=��r~�R�a��ܠ�v���A�ƋЁӋLƱ�	=�)����~��"�ֱ� �Q啉�jig�����`$<��U�lhe�j6�ܔq���$�kPj��~�>��M<U�A�I��ZR�}Je-Nr��W��6.�)�uc���*�w�qm������T(�����aj3Ȅ�q��w�S*d�!,�=�ޛ����7'a�Dǌ\>�њ�lF�Sh���C̛!%��� �� v|��xKw�p:��(,�"�:�hS�Y�}�5*�+3��T����L�躎�o��k��n͇���u��'͑6??�2@�A�4�ț����ߙ����<��:��.-��ד��{�!��bk~r������Ź�F��/����c������d���DG�b8�f��D�-.�'��X"���.z}���jKe �))��5���fZ���*���%K���9�8z��RS���7N\���o����8��A�z��tn�w����u�󴄮W]L7�1�8�׳ί������/��"VEv�!X�}礊lɔ߿n�d�0����ƈV�?Ȳ7��#�fF�t-/�EkDk}z�eۿi-1~�x��4����n�~9�:�]-���1r���A���F�#�^����V�o� ��gi���h�$��s�&����\ʗ��+c�+��f)%t]6Ql�w��kt����Y��XiCq��8�a����	�1j�>�a۳*x�B# dR���"��*\P��@�i`#ɞe���r���4D�o��A_���m�|��˂���P.N�}��x��BHr,�P�9�4J�96lLV��#92G��T[��t���%P�,��߷�ś��^�֑� ���`�(�sz��-�;'�^[��a��z�O�{��CD82\��]�f� t�5Vک�-�;\�8��J�ֵ��_�={�٧��s�P�G���X(6�P�o%���_+a��Z�,���iP(2� x$�"����E��6/3,�.?�?yÞ��G��.�o��=x���4,���:aH�C���UHi��y�N�uc���lPЛ����PZaE���2Q}�?u,%�c�޿� ���: ������l����+��1�֢0��1��,��g�ƅ��f0�GI?�,&����֫F��g�������.���V�a��j�/�2k/e��7�p�3Aƹ�p�c}�Y,D�'m7x��Ȯ�������(y��a@P���c���N欜X��nw������]��ɴ���m6�cP��x���$>B��>���zY��ڳ%���nH��R�jL�?n�q����WQ��2�[���YW�J�N�!��o�0�����T��<��S���#�6SC��E�����*�b�qX��N��Ihq�GP��y���q��&�0�9����ťy���X^��ڜ��m�s�����,ԥ�F������ �=�����n�T�9J{�j��ku>mr�;2�BH�1�`8��ۺ��0/�����_w��J�Q����}�;�$��#*��M�� �?U����&�GD&+�&ޛԼ�N�m��`�W�f<�j�U��1?yٓ�{��mϻ �~i��U���GX��H$C��y��.�駑nE$k�z'iA���M����W��\T�P]}�{�L��m��V� ��H	�/�c86+�7�m�]�<E�,؀�>
��6:m��NP��e�=�|�P�'V�8>����l�w8�a��F���9��իNyҍ)5h�M_�L�W����u�.��汀����+�x���t�����6�$X����R����������xo���;ԑb�A[��/�.�?��4���ڂ0��O�m��1�v<V�!��7���4ݬ�,G1���k���x�J�Uu.�iX�p���KS�2��n�5��&w$�SW2(���(4y?������n�E��z>uV��!��
 _�e4������w�:�+�HH��yT	��#@fm��[�=Q�
e8�NF�x��<�Ʈ�憩���ᜧ8�t#�Z^9=CP�~y����1�4|4�||)��4�T�>[�jN�G���{���7���.� �ȫ�Pƴ�%�I�u�ww]g��I�Q
�d��F�?�Y`�ݡ"�ℴ��ߎg�wH���V5��Z:��v7mOE�5;L�]�)���-�H��1�b��eϜ�^�RSm����Oc</.�­V��梭��C3D��8����<5�?�j��P�P�s���H0n��-�А%Q� �'5���l^^���AQN�c�|2�pAq��?I�sBk���d��X�4H��"��%��a\�ۆ��Qo7?��&�j�����f>I/��Q��'B\���'qy�j���/��I��@�:�v
��]�%��������'���D����$���B~�d�x_���S�����>:�����l/n�xT�C3�r�@�a����O��նr�e{))[j%�Ļ�D,��ћ�E��xUZ=�g����k�Xh}��|f�<ڃ����Y�+0����!�x́�>�~��hO�qz�6�&ݭej%�F�-(�?�8�q�������l̦C�;2%�Aa���_��n��������y�pXؕޚ�[����ݼm*�0�������mwa�}��&h4�: �>K\G�$SKe�}�dof�����;� �x,�A�:��f��w~�J�2�`��)�$$��o�qb4Lo�mζ �Ǎ��~�O�����z]��!�=�3"d��9庪�W��y�N�g� E6#�kT~��>�.�깔�](Y�Q��%``�(Fu�N|v��{�,�݀i�7�ױ.&�x/i2���V����0e�F����������<oY����D���1�b"'�w1-����w��`;�W>mHm�#9OV��_*��%���8(� �c=���NE:Z	�-~Һ�v������@�qb2¡w�Ću��No��g����qĩ�d�9㵝,,��p�Ev��D��.���ԫ��'GنG�=Lu++jp�?1G�p(�TL+EǱ�1�������z�ڛ�s��M�,$�,F-L��g����I~���꥚�hQT�C��"����^K��R~R��=��">,z;�ڜ��o�w���=v���oD͖˰n����=3�X�����J������R*�'��u�,��O�(JE;>Z�'���P�����-%��ʴ.����5۸��n�"����>v�"������٢�뫷8�f�n�\����QMZdmS�����
P�|�qzZ���7�K���������:Z4\��<.��z�F��<T�q�9Wk���_x��T2��-?x).�N���KIo�!}�$(7��K��c����$쇪�F].i(H[NK�����[UN��~+&M�T�BEX)K�ēb�f�6�E��;���u8�ey���~� �0ő�h'��!����'�_��t��>��|F�8p����Ӑɳ�9w,�+~��0��h_C�px�H�����-nI���j��u�����@I{�&�"~�9�ZFG��%u @����	w{v��v�Һ�?a��5(e]<�{��P^rd ��,��n#yr�v���¿�^	o������X�*�����=�ՀV���<��Ɇƣ۷�w�Z-�x3*P���:S������+gSŻ�"g7���������+ą��!H�P�,�1U֏��̋��u�̭3�N�Q�/9ЦZА[�s/d�+�F[�*Lzj@9X�1��
�U���Z9���I2�w�^���s�U�72A'Nɘ�w�z�-����@KG��T�W�Ii�S���
�����[�Gا�� �����+�-;�O��"�/� ���)_�:��bqI�h�z%x��q��"� { �D��[�3�c���+D�r�ew�?�Or�l6�0O�}"bb�FCȩR5���f�,� �Z�4�t�g�˫¼���~D{��:>�x������F��f����zdG
�ͺ�.d9��Yd�����-s��������>��cUj;�����И=>�U���v#7����(����>���D�OnG��ϕC2�lf�Ag�:�-��Ze�J�

v���J*҈��j�s�) �p��Z���\�Mk�	_�h+�EN_>�?B6>�s��y	�ds|�_1~��Y-��J�E۫V�~��Y�2;���8ˍ	���
q�}� k}��0\�g�l��溩�	F�0�����p/���K��.���ݕ�^���6�"A��9�����8�*�W�.�[�q�t���-=�e.::��J�b��c�%�t��Y�g��e�io'K'�6T���Z%7 r��HHB� �����	�(�ao��qƙ�wlT�?��->� E�b��������W���mNS�l6}��U�|� V�_�+��*n���-�����j�P�,w0�M��pO߭����dPc��L	9�i�:��wE����¿�L'+������X6���au�Y$���6�i���op�n���ۂ�(�fk}1!v��}N�e�	�F���1a���ˣ!�驔q���$_�����Qu)%�U�J�P�M 
 ���Z��ȰƷ�O�|���H2`N�ց�%cM@�>��:�|��a����l��
����a�xY����uO�38�$���Yї�gM�3  B!:���w`���G�����q�emz�-�M�uzk?�8�d6��̋<�Md���,��q�7�O_ � K�%�x>��(�9���TF(t"���}����.bl_�Qӗ�e|:����#3������S�m1�L"�g�����X�nv��7*��%-�1���4����z �˦7��Ww�\����,^�#v>���M��>��`ǡ��?`��:RrZ�9�F������A�8e[���np���e	$�+��S�/�6'H���U�i)���EsZ��J`%��.!/����"n�f���8��;�N�#��!3��Kf�h�;�����%���9�U�ȭ��'�-��uj���܁��f[Lls>{�؄G1�l^���M�	�P"Adh}�6�R�6uԶ����%O4b@y��RU^���N��?v�!�ẓ/�.L � ��M2B���g��,���N ��kQ�q��Af��&�w���+7���G�q�X����F���R�2Ƶ�stJ�ki��m�m˥JS��ʱ@oE�3`��A$�p�f��m<�?y���WI�P$�\K�q�+�҇��:��T<�IV�sO�����.3����@ޱ3��W��`/~)�)h3�#��v��OK�s1>�<L��>-y�0<+��{�S�e"w��i>^�_Wv�����K&́��j1�|Tx�.PBqw{D{��L�h$�*��ug/����r�;P$ޡ�l�H�~ �a$R>18�[H��p��;.�$*�ǤR=�M<�N��
Һ�d�)P���8�b��ȍX���붩�q�n�-��n(�ES�XJ���=�\%19��Kl}���i<Q�i9�)wl%	��Uz����6�O��!Ќ�iYo2�8R�i蜁4Yũ>�y	��I�:RR�%����.�m?�N�>y{Fޘ��U-��R����ArHA!��\en��F��2%�n:x�h@��"���Qj��GA�/$���d~���`��E����r)�5rzA��4ZImGĿה~mԒad�dꟀntz^�=���MQh@�2��J�-j��ǹ�ǎ�S�#��%ŧ�&�040��P�Gg>w�K�C�~b���)�ۢ�5�d7
.���x8'Ҍ�Z-�,x�t�YZ�9lx�O����-I�Uwy��n(j���AWr�:��t\﫠�B���E?��,�/�g9��H�.&*��D>yZ�Z"y���SŹ�a�p�&��ǗhM������[f�}D��|�o�0?x->q�Rþ��@vay0_-�Y�.߄�}"M�i] w Tym)�+A+>k�栋�[�S�$��Qgy�3�ɠ�� 9��b�'���X{�zޫ����X��VH�,)BK��$=���f4~XV��6���[�4�i���NP)�R�0�/�\F ����J�b�$�ӱ/�����|;�d�1�2�4v"kV��
��F��))(~4s{Oa��`	7��a�9�'f]�+�CHw��)a=��0�+�7���`�x�]��:38���d!{�Σ�����[}`���8�u�MHwkYr�S�dV`&fw�ľ���[:%�ʸFx�l'���(�[�Bl:#�y��O��k4������P��Q��Ͱ,���3cR�Y@��
Y� �cxN�/�O�I��m��²��\������� ^\�sRTۍIf:`\�e`S��sn��Lx_@O��v�s+�����z�"'�4	.����ʞ�;M���u������Bm	�y�����ֱ����h�&e憅�,@�U�vZQ;P#[ؖwxM������ۧ�$�ʕ�����*�e/Ҭx��p/�p-JϫP�<Ĺa~�§�x�%O@G�6T�}��}�oH�L:2��8� ��P���L�R���:��#AQ�Mx#��Ӕ~�l:�uf��#��CvAf�]��mT��h����U���G��>�M�7B���y�x��LiAնZ���6����0-�R�a��ʘa��9�{Cɺ��C��gc ���EЎ��N$�.���X��r]T��i��aU Uig�í�K�ƾx�`@K�G	HHs*Kּ	c}M(T���^�`�k�b0^�0����G�˵)	��9������^�!�����ࣖ�-���ѭI�m����cr���?ow�x�
]�G����J%k�j*�iW5����<��1ԛ�0m+�����c�ϊ��*(��u�k����]r�<�+ >\�S� �H�k>k
�Lr<$x1�:ʥ �ڄ��t�Hk�����#�&^ɀX���_��b'�|%�}��[nA�9��k�APM�$֯��"ap��ɡ����!��<�*���0z�Ei�B6)Օ�LDClg���-W�B=ʤ&�4��q��b29��CKK�X�7�%��}�P�ngK�^2���C���w���  H�gov����J�+��@�|ڊ���Ȫv3'K�a{�Uǂ��i!(g�Ch���7Ȱ|�+�,z���u`ؓ�H�رG��z���� ��b��ӈW��>�@��2� H�M�W�yȫ�s�h�e@��-����_.��h@�J�F����z4�#�0���=Ͽ��L���/�?Q@e�-/�����tS�qz���{b|��(=t0���U��L1��� �X) "�� ~�9�M��Ѩ��������{n�e�0�P�|�����:���r
'��(����E0]�n�Չ9����
➭��	������|�������q,�\�HD��֕��ɱ��v�j��	�j�Iо���89��h�����?��y``�EML��������._ˣbB�
<K u|��)�=|�����
L�0��M�z~���hVb��$a%��4��c b�O|@'�"��O����c�2���E"vg���Ae]y��MC��d��$+��v<����.���Z�!l1E<a؜� ��6��I�PI`��O�ba�;1��\]b���$0Q�+��hΏ]�v�ao��h�7[-���K]�/�䮡���ӹz�,��scg�c.��C�*a?J�	�ح�'�m?�ֲ���!Ԥm���JeNK�Pዏf@_�:�	>�L2�5�����)�2���F�z�rP�='� ��'m�#d���=]�ƒ����f25��F���3�T�������R��dM7�{� 
�xt���ٯ�Y{T�2�Pu�ڠ�8��FFrU0y�~N�&>c� @?>^;��dY$-|H�}%O+o�H]�P�+���C�v���G�ת�uߟJ����_����:�$�ٌ>`��@��U�1%�Y�K���b_K�ؖ�������P s�4�T��N�����$�X
Zg&����I�,ֶ���2��fG��+G��4������v3HGH��1̼���� d�����W�9�� ��1�&����*+��;���xQ"��l�9���L������p�����$s|�3>ó��В�*�ґ���X|[�m�2O)=9$mM�%�4�,� ��ܜ?b�+�M�e��N��X�~���5�m�B���_F��Õ9H��okgٔ�I��=�m'+z׻��k�4�]S�rcJ)�E�@xM�,�I%���@�e�Y6M�$D�3���-�˘�1�W�r|��������g���g3�W �ϟ���l�sBܠ��)n g���t�P{�f{��Ѝ�����}��帛�;KV#0�6 �Y �O�l��z�(c�\��m�Vw�c܊��-?�� �I/��]��� 6�X�%a�K�Ӗ�y��I���n`�h���'O��a2V�@��f��]V-�K`�1��S���a#�e���<��0u�F���s)\�~ ��h�^e�.k��-Mj�EN�~0&�M���O�>�S4}q�͡�W�`�M�XxL5B�������o# &����}D�6i.-A9��ɔ��x��.D�T�_����ma�a�|��9��@�����G�����a��
Y;3A���#�\˷uqU�Y'���p�&�t)����
��I���#
�iUِǋ}x>e `D�O�XAh��⧹`�j��EP!��P�1�6'�+�����t��	є���1��0*K���pk�[��Eڹ�!;���)�q��.�ZVA�^ʑl�|*Y��p�Ӥq?�z�0̋M�
�}D����t��,���o���r4�W�F��.7�5�?^d�Z�k9&{Fe��2�-��B۵@���맧�¸��	�=0���=��=J�����`�ܜS�9ئd�D�� ��/)6ʵ���?�?,����\���{��{ĸCP��Ѷ�L	�>�Q0�Į�H+�k�}�W�*Z
^���D� �(�/_�[�q��#{@��j_��)�*� М@����f���_��d6S}w`���G��ւ���0�g]~�`�6�4Ԏҡ�E�S��I"E�R�$ek=� ���?0��+�iقlB�2��%���ֆw�%��]*8C$�Nݒ��|D�K�ж�Pߐg�s��xVd��.�{d�񀸅[	��p���A�┊�7����1�p�;GHc^�.�bga��[��
���7�`�:��綩X�,~�7]E�/H9;���|������h���O�hd���o�BF{*��?h�2���qdqN���m���ui�Ρ�1���r�$Vs^�Q*����޽$X��E�����`8�G��jBb��G��U7;3�ugX"s�F'�����e-=B!:9�z�.E��{�[3-!��8R<F#�J�>�	2| �#��/E�(��%�*
T�=o�<e*Q}��_T���J>�w���X9�4}km���m�6A.P't��?�Fd��<f��kP�a��sx�7�[C_���!Ѹ�ml�E?&��L`>���#���^��*Cb^>j��7$Ke���+��=�0χ����k�]tC���֎����;�q)o����~�)��I�D����'�$���*��(f�N����FD��m¥s{d� �^g��u��hf��LS���S�|(�W-}RTb�ޞْC�ّ�	?������&����<���d�l�$B���(iI�E?`���ޯh��GZ�<�IlS�89�UoeϪ����u��Ѭ�AE��C�ZAR�Hr҉��a����@�*�Kfo��o�*��K��L�<:�>Z�������w̸��<8���~����r��e�+*GC����Ľ�?��	�7re��ސǎr?�md�1�D�Eʡ�O��b���)�Jp�ipF+�%��|aѦ�qe�>n�c�Dg���V�-���m*t�m��-i�����)�4Qb��	y�+M�x���M�|}����vW����L~'��U!�
�.�\���-"��������]��l�TG$B����p��q�ߝ�Q�3��-� �O�J#�* ��t\�SS���A�����}�]}�>� p��پ�0��'�i�#���:���-���}�Cѻr��*`��ǟX�2׈�)��74�'d�痄�[Pm�����_�<�c���gY���p��Y����ۮ���8�P/��|p�ف�^h�}y����zLz�_��͘�]�V���&G�Ɔ5Ԋ1�䩲���=���ǜ�[���>|-m���ג{�b��r�FO�7�ݏ
%%oZ�U������jl��!A�42,�*)$���ٸ�X��:���G&��}O��s�_P�U��z����7�;E>�w�.��?�fu��=n]�e@e�%��wI>$�f �	"��+=WN��(h)A��Ys��ɹU�����^fGY���twঙ�|��2X$���
������@��V��c�-f���B�3S�=�'�2V�q�P?��` r&���o��I��L+�n��g^d�l�r�U`��;��7I��-�[]��m$�Ѓ�������� ��_*�>��m���O}���0`��-6�p���C)�m�٣`�cu"�����) �*��-��%��j�3�n�#sﮂ7	/꣥B�(9���Z&���n�c�;�z5-pInq?�=9�^1���?���
4ɔ��k")��n�w�EAmL3�Z�qD2�E��������ou���Ef���D�r:eXFv:����Ќ���Z�]h=Q�:�G��_x0Q�-�dOG���@O�8(B�t7��xz8�_\��7����W7>���h��&�D��,��qaVDX
��.͂�YZ��κp�o�-�7�W���H=Y�^�n�W9�
��W$tb�G?i���R,��܋u!TlaR����>}BB h���kyf#ƛ���.}�	����
ޠ5]�#&f�˒�R������4?� ݐ
/(艼�l-o�d������E��E��H�4��*�B����Pz<�F��� �.,I���1͙�Mmj��.�Z�����f� ��?w������X�`���@sV!��T�r�.��oo=BK�c3=h��˄��MI�F.`�c����<�=_����?���~\�4��ySB�b�~��=��7������G���8��-����|uQ3�}�����7��?��wgA�2�U9�T�_��Ӱ�$���pZ�|��E!��Z�(8��@�v&���BdtSJF%I�j��E���o��(�f��cK�sj9	��T�� �*�:��ȳ����q{{���a��c��7���f��6�a�Aptw��+��1�*=f��4��[��ͯ�ȴ�H{��Ӕ OW��]*~���I�� �l����n�T�sI����Q�4�,�M����n�{��/�u�i
�(�$���8���Ci�2[���Sc .}L 5[뭸ֱ}B����n�hb����S���3�(x"X�)�ek�Ѵ�x�b*��[gT�e��?]]��0<�����H��ƪ��0�IG��߭?7��q"� ����r�j�W�K~0�2��cҝ��t)�ө�`Q��"��'�k~�tBE���7Ὑ����?q�B7E%�*����$�u1q���?Q%���}���dQ��]�� oH��I���c�7\ǰ�{/���Wǔnm�cp9�P�_�P��
�-1{��grJ$T��7hr��F�/k7Ý��aa�&�k�D�e���#MR�g&�;]͔9�Pɼ�l�}�ԝ�lC0��%��qX�r�s{�%;��(������X�)��~CS�e��X֗��O�\;���H�A��{L�%�V8��|:�H���˚_�I���YUI�]b���W�_��l��^쁜��~2��9h�_�ԟ��B_�o���<6���<�&�v/�n�����|R���H����LH��6TQ��#�Ԣv1��<�^�C���.����-%1�5��yNr���<�J��,��V��R�����>A�|����,��fSj�=~�]	Һ�c�A��8L�%�6��[�,BY�)O))킳��,0D�N�.7���,�揬辕^fh�'
�$���]�ӿI���B����V��"�;ݒ�q��!�A�5Ӳ�z�%�_7Z�a%:�Q���+��}��V�7�{��W�F��?��4�5��vp�ٳسC�O�&V��9����le0�(/t�����+曀�]�pQ���.+�u�\�x`�9s
�kBc�Q�I8
�[�G��)�˝�o�1NwUՠp��f�,�����VX��6���bn!�e�C�O�?ɏ*�x!sE��i���]nD��B�!�=)�EPF[k�ԏ=o{0y�'�E��.�~�U�Fp��[է�-K��d�D��=���5tK��΋ѩw_Մ*{��d?��=����	�N�t*N�sN�JŰ^_����V��4��~V�n�Z\Bh���g��4<I1�-C�\-k&��,��P	�*ƍ��k
�ޒ,��)�->:��z��A�>��	�<�e]
�w��v7�G�Wi����3�w�/���C�lϬ�w�G���I��ND���#�����Lwµ���tF�0N�u� J���z���[3~��;r�!ji�Tr��Y?2��ba]Q�Q�IB�]�x��=#�a�w44=D�g֋v�S�4�����#O&m+�\����Y*���H]�*N�|*���Dy����1��^k�G��f�`,������)���W\�f���6i�,�v�>�(���T*��V����ߟ{�L��e�Y5#��6ng���T�� x�zd?���VB?�qEv=_ws��X<��.&��4�NX�����6'�����]r�$��,��I���R�k��?M�х�h�@��&XX4����5I#��c�if�r�ց������d����&�s�`Mq�,k����PN��_��imd&ά�6��f��1�)
H�rD��\��Z�ƞ���hu<�R��.�(
�B5g�1<a�9Ү���S "��#��R�Y}�Z�R2X��I����+��F�Yj���]�F�DзGtX2[��vC�;�t�Y����c4bt��nWs*.����oD���3%�m}�֔�X�e�:a,3/�2%�P�Y��uG�4}�{2��/Y�����5KLFs4���}�nH�a恍6��=��F9�.���3��`��Aʹ��:��U�)���ǯ7�\�I�Ǌ�O��	�u���5���i놂�Yn�Z�i߇�w���������څ�N�]���gݺ�"�r"�6q������0�ab47�P�$��1V�F�zL*~�bz�a+F5�w�����J�2$@B^Y�����rv&��m�Y�4��HG�4a����ĭ��[!�ԂZ�b�Z!�)���\��p(�B�&�0)��������-.�aO`�f�O1��G��"L�H�<�Ԝ�c�W+��X}���1{؎�e�\�=��z�Sδ{������l
�Ia�1�]mM<%�U�r�F�,���=K��c'�ڠ�����H�^��_S�&�S��_w��Q�n/���e�5�8p����ه<��D}�8wm������أ���ͯ���	�D����U���T�)܇ۊ�}�@�MF[Wza��B6�v�K<b�F)	'̞�	����_�ؗ��YL�a�K�r	C�Hj�l?7U�XÐ��ZOZ��k���'�Q���� h8=��?���Gl>�2*h0�G�n������T��ᯌS��� �I�.))�M�nW�x�D]��v��]�:�O\��t����霻�=K���.R�bBl�C�2M�����Er<� ?����.x���m��~F(��ךd�x��jQ����+Hį
�3ed?*�������4èW��tҵ0�F�v�v)�%͇�o��`Q�V8
:k+Pw]"WV��E�������l����{n�-�0�0|і2�w�WO���͏���_8tH�X� �_2��Ģ]l"}�׌d'���?�oT��:h
[O�]���3�|���9���o�ĸSPu����a�4�U��T6�j���>"�	��JA�\8� �v��? $mP4j7�F��o��\u�	�7]�g�kyΟ\,~�$e��\#��{���w�W�j�dEq��s�C[&����e�oR$i#���=0�R:���푦V��͎�%���m7�I!AfirvU�*Y��6Y!�7ݤ�A�q|�p��%Xθ��z��[���>�Ea�v���`�5��-a*��Y��ڟ�}]����9��2�Q��9V��G�č9�MV�o	&(�F|<�:����s⬲���!���7��`k�n�rX�y��隊����n�A��ux��AQ;�:��J(���	%o��+qp�pz5��B�`��A�f~��6�Xq�i�3������j�RJ��ּ��zȚ1Cy�sLtnuі�2t �jn�),�Ah%���e{��?��B�_��^V���|e�*��+�0�di���&���=�[(�����3�׬�k��J$:��/m]�qnyso�q/W-�eJ��.�p��B2�b;.�
M%z�R��;��f���H�W���1���c�=͜�Tr�,qL̺By�cmv����ɂx�L��`����>Ĕ�Q��%�ӾS�DpK� \Ⱥ���m���u���2�9bQ�@��Vm�� �:V�[l6����ot�^�X#�1PGTWo��e)l�ߩ<#t���ޏS&rF������g&�0�E������VW`�G7���^Wn�\O�8��ƅmɩ��S�T�jwQZ�\�h�Z&2dn��y����Eva�E�.Z0�������%rm	plA-��!m��6\9��W�A��*�����5&���,4Ӣ�s^�Y��FL`�:�,^��c��:g��w0KiB���m����&�Ҩ=h4"K��lɂ�oz��B"�,T���7�����B"��m�S\�ij|�����#o�I���d	�.��\�{��th�x�Y�*s�X���\8#b{{NZB�Wl����Q�-:�Qƣ
�81P��dg�`ݪ4q�4�q-r��(�?�!T�BI=D��*k��������&�Ȋ1a'.��dC0���?v�ib�q,��2xOi�y[p,E`wM�ΑUpuć�)�'�[�Έ�!�4Nӯ�i,7���i��p]�-���l0^l�m\X+��U0ƽ�J)�E�W��d9�?�Z���!���wd�j�d��\P0�7'�K�[�%b���&q~��^iL�[�!�S|���˯p
C����D`(8�j"/�}��h�^����������?6־U���֪�����y��P���3+�Z4���{��c>�1̒ȳ��n���޼Up�v�&zC�^�� ��=�Ҳ�#�/}�7z�����$�7��X��n4N_�M�+�"���Fw�BؼϪ����m�V7E��%��c��f"~��X�ϋ.E���8�w�r�%�;�7��s@98u�?ud���N��U8��b �ޛ��Pti��	2�H���f{c�+Hp�H�:��=�V\�Wr$91�QW���rU2P��܏�A�70%�<�'���+Af��yOm����$�rO�$��W`����/�hj\�9h�/�~=nIv�����?�D#�_ێ�Yasu�P6 n��,M��{x`q�M����v]w�����?����W�9缎�/��Q��egK{�zJ���jp��>D���#h�-���� d���59����&�V\6]C�;��$��OO�% ��0��gH�*d�GW3�-
����)���t�X��9�7͹�����,ٷD%���0�=����նKF��jv��eːz����޶ s~Qi�SأQ%U��7̀/�G	aU���:�Fɚޟ�RpEU�B�G�2���[��c�)kJ��cW9�Ǝ]Q���u�o�4k.G��/�l.A��O�՗��t0�T&�6�qpo�]�uF��?��[N9�*B*�|M�x��HV�@�荕-P��*1B����F�fq@t�Ci�^�ل_w{����)T�rmjK�Qo}�x+�_�DÉڮ�T�(�<y@�o**tW����ʫ� 	őN�`ܔE'"2�F�4#�Lҥ�&9�Jh�M��l�u\��7.P�+��6�ܬO�	�����$��e�����Ax����쉰y������ �~��&\��hK�����
�L��+�s2��c�&����(0^t���N#^v��7Z
5��{��t:���8𪶮п�t8%̼g����	��wRo5����*���8zζ��d��:/Q��D)�/mS<�4�'7�xP��ɦL�> H�c��� 衚&W�\P&�h`�q2�\��4����38����b �Pɬ�@^2�E_�]M�Gx�f���3�Շwa�����aQ_���QqL�;Ϭ'6Z�O�&�
 W�h����i��1p*/�g�ҷņ8��Oz��!��sU^۶`�Q�^�(Õ�D~���]M4jF
��<���8�ý�(f�]L��M��b�V����x�fe�WȠǭ�f�k�lD��[fԓ/~�ڬp���O��C)�`���2��Ba